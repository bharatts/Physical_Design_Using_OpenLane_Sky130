module picorv32a (clk,
    resetn,
    trap,
    mem_valid,
    mem_instr,
    mem_ready,
    mem_addr,
    mem_wdata,
    mem_wstrb,
    mem_rdata,
    mem_la_read,
    mem_la_write,
    mem_la_addr,
    mem_la_wdata,
    mem_la_wstrb,
    pcpi_valid,
    pcpi_insn,
    pcpi_rs1,
    pcpi_rs2,
    pcpi_wr,
    pcpi_rd,
    pcpi_wait,
    pcpi_ready,
    irq,
    eoi,
    trace_valid,
    trace_data);
 input clk;
 input resetn;
 output trap;
 output mem_valid;
 output mem_instr;
 input mem_ready;
 output [31:0] mem_addr;
 output [31:0] mem_wdata;
 output [3:0] mem_wstrb;
 input [31:0] mem_rdata;
 output mem_la_read;
 output mem_la_write;
 output [31:0] mem_la_addr;
 output [31:0] mem_la_wdata;
 output [3:0] mem_la_wstrb;
 output pcpi_valid;
 output [31:0] pcpi_insn;
 output [31:0] pcpi_rs1;
 output [31:0] pcpi_rs2;
 input pcpi_wr;
 input [31:0] pcpi_rd;
 input pcpi_wait;
 input pcpi_ready;
 input [31:0] irq;
 output [31:0] eoi;
 output trace_valid;
 output [35:0] trace_data;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire _06911_;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire _06965_;
 wire _06966_;
 wire _06967_;
 wire _06968_;
 wire _06969_;
 wire _06970_;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire _06982_;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire _06987_;
 wire _06988_;
 wire _06989_;
 wire _06990_;
 wire _06991_;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire _07000_;
 wire _07001_;
 wire _07002_;
 wire _07003_;
 wire _07004_;
 wire _07005_;
 wire _07006_;
 wire _07007_;
 wire _07008_;
 wire _07009_;
 wire _07010_;
 wire _07011_;
 wire _07012_;
 wire _07013_;
 wire _07014_;
 wire _07015_;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire _07019_;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire _07023_;
 wire _07024_;
 wire _07025_;
 wire _07026_;
 wire _07027_;
 wire _07028_;
 wire _07029_;
 wire _07030_;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire _07034_;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire _07038_;
 wire _07039_;
 wire _07040_;
 wire _07041_;
 wire _07042_;
 wire _07043_;
 wire _07044_;
 wire _07045_;
 wire _07046_;
 wire _07047_;
 wire _07048_;
 wire _07049_;
 wire _07050_;
 wire _07051_;
 wire _07052_;
 wire _07053_;
 wire _07054_;
 wire _07055_;
 wire _07056_;
 wire _07057_;
 wire _07058_;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire _07063_;
 wire _07064_;
 wire _07065_;
 wire _07066_;
 wire _07067_;
 wire _07068_;
 wire _07069_;
 wire _07070_;
 wire _07071_;
 wire _07072_;
 wire _07073_;
 wire _07074_;
 wire _07075_;
 wire _07076_;
 wire _07077_;
 wire _07078_;
 wire _07079_;
 wire _07080_;
 wire _07081_;
 wire _07082_;
 wire _07083_;
 wire _07084_;
 wire _07085_;
 wire _07086_;
 wire _07087_;
 wire _07088_;
 wire _07089_;
 wire _07090_;
 wire _07091_;
 wire _07092_;
 wire _07093_;
 wire _07094_;
 wire _07095_;
 wire _07096_;
 wire _07097_;
 wire _07098_;
 wire _07099_;
 wire _07100_;
 wire _07101_;
 wire _07102_;
 wire _07103_;
 wire _07104_;
 wire _07105_;
 wire _07106_;
 wire _07107_;
 wire _07108_;
 wire _07109_;
 wire _07110_;
 wire _07111_;
 wire _07112_;
 wire _07113_;
 wire _07114_;
 wire _07115_;
 wire _07116_;
 wire _07117_;
 wire _07118_;
 wire _07119_;
 wire _07120_;
 wire _07121_;
 wire _07122_;
 wire _07123_;
 wire _07124_;
 wire _07125_;
 wire _07126_;
 wire _07127_;
 wire _07128_;
 wire _07129_;
 wire _07130_;
 wire _07131_;
 wire _07132_;
 wire _07133_;
 wire _07134_;
 wire _07135_;
 wire _07136_;
 wire _07137_;
 wire _07138_;
 wire _07139_;
 wire _07140_;
 wire _07141_;
 wire _07142_;
 wire _07143_;
 wire _07144_;
 wire _07145_;
 wire _07146_;
 wire _07147_;
 wire _07148_;
 wire _07149_;
 wire _07150_;
 wire _07151_;
 wire _07152_;
 wire _07153_;
 wire _07154_;
 wire _07155_;
 wire _07156_;
 wire _07157_;
 wire _07158_;
 wire _07159_;
 wire _07160_;
 wire _07161_;
 wire _07162_;
 wire _07163_;
 wire _07164_;
 wire _07165_;
 wire _07166_;
 wire _07167_;
 wire _07168_;
 wire _07169_;
 wire _07170_;
 wire _07171_;
 wire _07172_;
 wire _07173_;
 wire _07174_;
 wire _07175_;
 wire _07176_;
 wire _07177_;
 wire _07178_;
 wire _07179_;
 wire _07180_;
 wire _07181_;
 wire _07182_;
 wire _07183_;
 wire _07184_;
 wire _07185_;
 wire _07186_;
 wire _07187_;
 wire _07188_;
 wire _07189_;
 wire _07190_;
 wire _07191_;
 wire _07192_;
 wire _07193_;
 wire _07194_;
 wire _07195_;
 wire _07196_;
 wire _07197_;
 wire _07198_;
 wire _07199_;
 wire _07200_;
 wire _07201_;
 wire _07202_;
 wire _07203_;
 wire _07204_;
 wire _07205_;
 wire _07206_;
 wire _07207_;
 wire _07208_;
 wire _07209_;
 wire _07210_;
 wire _07211_;
 wire _07212_;
 wire _07213_;
 wire _07214_;
 wire _07215_;
 wire _07216_;
 wire _07217_;
 wire _07218_;
 wire _07219_;
 wire _07220_;
 wire _07221_;
 wire _07222_;
 wire _07223_;
 wire _07224_;
 wire _07225_;
 wire _07226_;
 wire _07227_;
 wire _07228_;
 wire _07229_;
 wire _07230_;
 wire _07231_;
 wire _07232_;
 wire _07233_;
 wire _07234_;
 wire _07235_;
 wire _07236_;
 wire _07237_;
 wire _07238_;
 wire _07239_;
 wire _07240_;
 wire _07241_;
 wire _07242_;
 wire _07243_;
 wire _07244_;
 wire _07245_;
 wire _07246_;
 wire _07247_;
 wire _07248_;
 wire _07249_;
 wire _07250_;
 wire _07251_;
 wire _07252_;
 wire _07253_;
 wire _07254_;
 wire _07255_;
 wire _07256_;
 wire _07257_;
 wire _07258_;
 wire _07259_;
 wire _07260_;
 wire _07261_;
 wire _07262_;
 wire _07263_;
 wire _07264_;
 wire _07265_;
 wire _07266_;
 wire _07267_;
 wire _07268_;
 wire _07269_;
 wire _07270_;
 wire _07271_;
 wire _07272_;
 wire _07273_;
 wire _07274_;
 wire _07275_;
 wire _07276_;
 wire _07277_;
 wire _07278_;
 wire _07279_;
 wire _07280_;
 wire _07281_;
 wire _07282_;
 wire _07283_;
 wire _07284_;
 wire _07285_;
 wire _07286_;
 wire _07287_;
 wire _07288_;
 wire _07289_;
 wire _07290_;
 wire _07291_;
 wire _07292_;
 wire _07293_;
 wire _07294_;
 wire _07295_;
 wire _07296_;
 wire _07297_;
 wire _07298_;
 wire _07299_;
 wire _07300_;
 wire _07301_;
 wire _07302_;
 wire _07303_;
 wire _07304_;
 wire _07305_;
 wire _07306_;
 wire _07307_;
 wire _07308_;
 wire _07309_;
 wire _07310_;
 wire _07311_;
 wire _07312_;
 wire _07313_;
 wire _07314_;
 wire _07315_;
 wire _07316_;
 wire _07317_;
 wire _07318_;
 wire _07319_;
 wire _07320_;
 wire _07321_;
 wire _07322_;
 wire _07323_;
 wire _07324_;
 wire _07325_;
 wire _07326_;
 wire _07327_;
 wire _07328_;
 wire _07329_;
 wire _07330_;
 wire _07331_;
 wire _07332_;
 wire _07333_;
 wire _07334_;
 wire _07335_;
 wire _07336_;
 wire _07337_;
 wire _07338_;
 wire _07339_;
 wire _07340_;
 wire _07341_;
 wire _07342_;
 wire _07343_;
 wire _07344_;
 wire _07345_;
 wire _07346_;
 wire _07347_;
 wire _07348_;
 wire _07349_;
 wire _07350_;
 wire _07351_;
 wire _07352_;
 wire _07353_;
 wire _07354_;
 wire _07355_;
 wire _07356_;
 wire _07357_;
 wire _07358_;
 wire _07359_;
 wire _07360_;
 wire _07361_;
 wire _07362_;
 wire _07363_;
 wire _07364_;
 wire _07365_;
 wire _07366_;
 wire _07367_;
 wire _07368_;
 wire _07369_;
 wire _07370_;
 wire _07371_;
 wire _07372_;
 wire _07373_;
 wire _07374_;
 wire _07375_;
 wire _07376_;
 wire _07377_;
 wire _07378_;
 wire _07379_;
 wire _07380_;
 wire _07381_;
 wire _07382_;
 wire _07383_;
 wire _07384_;
 wire _07385_;
 wire _07386_;
 wire _07387_;
 wire _07388_;
 wire _07389_;
 wire _07390_;
 wire _07391_;
 wire _07392_;
 wire _07393_;
 wire _07394_;
 wire _07395_;
 wire _07396_;
 wire _07397_;
 wire _07398_;
 wire _07399_;
 wire _07400_;
 wire _07401_;
 wire _07402_;
 wire _07403_;
 wire _07404_;
 wire _07405_;
 wire _07406_;
 wire _07407_;
 wire _07408_;
 wire _07409_;
 wire _07410_;
 wire _07411_;
 wire _07412_;
 wire _07413_;
 wire _07414_;
 wire _07415_;
 wire _07416_;
 wire _07417_;
 wire _07418_;
 wire _07419_;
 wire _07420_;
 wire _07421_;
 wire _07422_;
 wire _07423_;
 wire _07424_;
 wire _07425_;
 wire _07426_;
 wire _07427_;
 wire _07428_;
 wire _07429_;
 wire _07430_;
 wire _07431_;
 wire _07432_;
 wire _07433_;
 wire _07434_;
 wire _07435_;
 wire _07436_;
 wire _07437_;
 wire _07438_;
 wire _07439_;
 wire _07440_;
 wire _07441_;
 wire _07442_;
 wire _07443_;
 wire _07444_;
 wire _07445_;
 wire _07446_;
 wire _07447_;
 wire _07448_;
 wire _07449_;
 wire _07450_;
 wire _07451_;
 wire _07452_;
 wire _07453_;
 wire _07454_;
 wire _07455_;
 wire _07456_;
 wire _07457_;
 wire _07458_;
 wire _07459_;
 wire _07460_;
 wire _07461_;
 wire _07462_;
 wire _07463_;
 wire _07464_;
 wire _07465_;
 wire _07466_;
 wire _07467_;
 wire _07468_;
 wire _07469_;
 wire _07470_;
 wire _07471_;
 wire _07472_;
 wire _07473_;
 wire _07474_;
 wire _07475_;
 wire _07476_;
 wire _07477_;
 wire _07478_;
 wire _07479_;
 wire _07480_;
 wire _07481_;
 wire _07482_;
 wire _07483_;
 wire _07484_;
 wire _07485_;
 wire _07486_;
 wire _07487_;
 wire _07488_;
 wire _07489_;
 wire _07490_;
 wire _07491_;
 wire _07492_;
 wire _07493_;
 wire _07494_;
 wire _07495_;
 wire _07496_;
 wire _07497_;
 wire _07498_;
 wire _07499_;
 wire _07500_;
 wire _07501_;
 wire _07502_;
 wire _07503_;
 wire _07504_;
 wire _07505_;
 wire _07506_;
 wire _07507_;
 wire _07508_;
 wire _07509_;
 wire _07510_;
 wire _07511_;
 wire _07512_;
 wire _07513_;
 wire _07514_;
 wire _07515_;
 wire _07516_;
 wire _07517_;
 wire _07518_;
 wire _07519_;
 wire _07520_;
 wire _07521_;
 wire _07522_;
 wire _07523_;
 wire _07524_;
 wire _07525_;
 wire _07526_;
 wire _07527_;
 wire _07528_;
 wire _07529_;
 wire _07530_;
 wire _07531_;
 wire _07532_;
 wire _07533_;
 wire _07534_;
 wire _07535_;
 wire _07536_;
 wire _07537_;
 wire _07538_;
 wire _07539_;
 wire _07540_;
 wire _07541_;
 wire _07542_;
 wire _07543_;
 wire _07544_;
 wire _07545_;
 wire _07546_;
 wire _07547_;
 wire _07548_;
 wire _07549_;
 wire _07550_;
 wire _07551_;
 wire _07552_;
 wire _07553_;
 wire _07554_;
 wire _07555_;
 wire _07556_;
 wire _07557_;
 wire _07558_;
 wire _07559_;
 wire _07560_;
 wire _07561_;
 wire _07562_;
 wire _07563_;
 wire _07564_;
 wire _07565_;
 wire _07566_;
 wire _07567_;
 wire _07568_;
 wire _07569_;
 wire _07570_;
 wire _07571_;
 wire _07572_;
 wire _07573_;
 wire _07574_;
 wire _07575_;
 wire _07576_;
 wire _07577_;
 wire _07578_;
 wire _07579_;
 wire _07580_;
 wire _07581_;
 wire _07582_;
 wire _07583_;
 wire _07584_;
 wire _07585_;
 wire _07586_;
 wire _07587_;
 wire _07588_;
 wire _07589_;
 wire _07590_;
 wire _07591_;
 wire _07592_;
 wire _07593_;
 wire _07594_;
 wire _07595_;
 wire _07596_;
 wire _07597_;
 wire _07598_;
 wire _07599_;
 wire _07600_;
 wire _07601_;
 wire _07602_;
 wire _07603_;
 wire _07604_;
 wire _07605_;
 wire _07606_;
 wire _07607_;
 wire _07608_;
 wire _07609_;
 wire _07610_;
 wire _07611_;
 wire _07612_;
 wire _07613_;
 wire _07614_;
 wire _07615_;
 wire _07616_;
 wire _07617_;
 wire _07618_;
 wire _07619_;
 wire _07620_;
 wire _07621_;
 wire _07622_;
 wire _07623_;
 wire _07624_;
 wire _07625_;
 wire _07626_;
 wire _07627_;
 wire _07628_;
 wire _07629_;
 wire _07630_;
 wire _07631_;
 wire _07632_;
 wire _07633_;
 wire _07634_;
 wire _07635_;
 wire _07636_;
 wire _07637_;
 wire _07638_;
 wire _07639_;
 wire _07640_;
 wire _07641_;
 wire _07642_;
 wire _07643_;
 wire _07644_;
 wire _07645_;
 wire _07646_;
 wire _07647_;
 wire _07648_;
 wire _07649_;
 wire _07650_;
 wire _07651_;
 wire _07652_;
 wire _07653_;
 wire _07654_;
 wire _07655_;
 wire _07656_;
 wire _07657_;
 wire _07658_;
 wire _07659_;
 wire _07660_;
 wire _07661_;
 wire _07662_;
 wire _07663_;
 wire _07664_;
 wire _07665_;
 wire _07666_;
 wire _07667_;
 wire _07668_;
 wire _07669_;
 wire _07670_;
 wire _07671_;
 wire _07672_;
 wire _07673_;
 wire _07674_;
 wire _07675_;
 wire _07676_;
 wire _07677_;
 wire _07678_;
 wire _07679_;
 wire _07680_;
 wire _07681_;
 wire _07682_;
 wire _07683_;
 wire _07684_;
 wire _07685_;
 wire _07686_;
 wire _07687_;
 wire _07688_;
 wire _07689_;
 wire _07690_;
 wire _07691_;
 wire _07692_;
 wire _07693_;
 wire _07694_;
 wire _07695_;
 wire _07696_;
 wire _07697_;
 wire _07698_;
 wire _07699_;
 wire _07700_;
 wire _07701_;
 wire _07702_;
 wire _07703_;
 wire _07704_;
 wire _07705_;
 wire _07706_;
 wire _07707_;
 wire _07708_;
 wire _07709_;
 wire _07710_;
 wire _07711_;
 wire _07712_;
 wire _07713_;
 wire _07714_;
 wire _07715_;
 wire _07716_;
 wire _07717_;
 wire _07718_;
 wire _07719_;
 wire _07720_;
 wire _07721_;
 wire _07722_;
 wire _07723_;
 wire _07724_;
 wire _07725_;
 wire _07726_;
 wire _07727_;
 wire _07728_;
 wire _07729_;
 wire _07730_;
 wire _07731_;
 wire _07732_;
 wire _07733_;
 wire _07734_;
 wire _07735_;
 wire _07736_;
 wire _07737_;
 wire _07738_;
 wire _07739_;
 wire _07740_;
 wire _07741_;
 wire _07742_;
 wire _07743_;
 wire _07744_;
 wire _07745_;
 wire _07746_;
 wire _07747_;
 wire _07748_;
 wire _07749_;
 wire _07750_;
 wire _07751_;
 wire _07752_;
 wire _07753_;
 wire _07754_;
 wire _07755_;
 wire _07756_;
 wire _07757_;
 wire _07758_;
 wire _07759_;
 wire _07760_;
 wire _07761_;
 wire _07762_;
 wire _07763_;
 wire _07764_;
 wire _07765_;
 wire _07766_;
 wire _07767_;
 wire _07768_;
 wire _07769_;
 wire _07770_;
 wire _07771_;
 wire _07772_;
 wire _07773_;
 wire _07774_;
 wire _07775_;
 wire _07776_;
 wire _07777_;
 wire _07778_;
 wire _07779_;
 wire _07780_;
 wire _07781_;
 wire _07782_;
 wire _07783_;
 wire _07784_;
 wire _07785_;
 wire _07786_;
 wire _07787_;
 wire _07788_;
 wire _07789_;
 wire _07790_;
 wire _07791_;
 wire _07792_;
 wire _07793_;
 wire _07794_;
 wire _07795_;
 wire _07796_;
 wire _07797_;
 wire _07798_;
 wire _07799_;
 wire _07800_;
 wire _07801_;
 wire _07802_;
 wire _07803_;
 wire _07804_;
 wire _07805_;
 wire _07806_;
 wire _07807_;
 wire _07808_;
 wire _07809_;
 wire _07810_;
 wire _07811_;
 wire _07812_;
 wire _07813_;
 wire _07814_;
 wire _07815_;
 wire _07816_;
 wire _07817_;
 wire _07818_;
 wire _07819_;
 wire _07820_;
 wire _07821_;
 wire _07822_;
 wire _07823_;
 wire _07824_;
 wire _07825_;
 wire _07826_;
 wire _07827_;
 wire _07828_;
 wire _07829_;
 wire _07830_;
 wire _07831_;
 wire _07832_;
 wire _07833_;
 wire _07834_;
 wire _07835_;
 wire _07836_;
 wire _07837_;
 wire _07838_;
 wire _07839_;
 wire _07840_;
 wire _07841_;
 wire _07842_;
 wire _07843_;
 wire _07844_;
 wire _07845_;
 wire _07846_;
 wire _07847_;
 wire _07848_;
 wire _07849_;
 wire _07850_;
 wire _07851_;
 wire _07852_;
 wire _07853_;
 wire _07854_;
 wire _07855_;
 wire _07856_;
 wire _07857_;
 wire _07858_;
 wire _07859_;
 wire _07860_;
 wire _07861_;
 wire _07862_;
 wire _07863_;
 wire _07864_;
 wire _07865_;
 wire _07866_;
 wire _07867_;
 wire _07868_;
 wire _07869_;
 wire _07870_;
 wire _07871_;
 wire _07872_;
 wire _07873_;
 wire _07874_;
 wire _07875_;
 wire _07876_;
 wire _07877_;
 wire _07878_;
 wire _07879_;
 wire _07880_;
 wire _07881_;
 wire _07882_;
 wire _07883_;
 wire _07884_;
 wire _07885_;
 wire _07886_;
 wire _07887_;
 wire _07888_;
 wire _07889_;
 wire _07890_;
 wire _07891_;
 wire _07892_;
 wire _07893_;
 wire _07894_;
 wire _07895_;
 wire _07896_;
 wire _07897_;
 wire _07898_;
 wire _07899_;
 wire _07900_;
 wire _07901_;
 wire _07902_;
 wire _07903_;
 wire _07904_;
 wire _07905_;
 wire _07906_;
 wire _07907_;
 wire _07908_;
 wire _07909_;
 wire _07910_;
 wire _07911_;
 wire _07912_;
 wire _07913_;
 wire _07914_;
 wire _07915_;
 wire _07916_;
 wire _07917_;
 wire _07918_;
 wire _07919_;
 wire _07920_;
 wire _07921_;
 wire _07922_;
 wire _07923_;
 wire _07924_;
 wire _07925_;
 wire _07926_;
 wire _07927_;
 wire _07928_;
 wire _07929_;
 wire _07930_;
 wire _07931_;
 wire _07932_;
 wire _07933_;
 wire _07934_;
 wire _07935_;
 wire _07936_;
 wire _07937_;
 wire _07938_;
 wire _07939_;
 wire _07940_;
 wire _07941_;
 wire _07942_;
 wire _07943_;
 wire _07944_;
 wire _07945_;
 wire _07946_;
 wire _07947_;
 wire _07948_;
 wire _07949_;
 wire _07950_;
 wire _07951_;
 wire _07952_;
 wire _07953_;
 wire _07954_;
 wire _07955_;
 wire _07956_;
 wire _07957_;
 wire _07958_;
 wire _07959_;
 wire _07960_;
 wire _07961_;
 wire _07962_;
 wire _07963_;
 wire _07964_;
 wire _07965_;
 wire _07966_;
 wire _07967_;
 wire _07968_;
 wire _07969_;
 wire _07970_;
 wire _07971_;
 wire _07972_;
 wire _07973_;
 wire _07974_;
 wire _07975_;
 wire _07976_;
 wire _07977_;
 wire _07978_;
 wire _07979_;
 wire _07980_;
 wire _07981_;
 wire _07982_;
 wire _07983_;
 wire _07984_;
 wire _07985_;
 wire _07986_;
 wire _07987_;
 wire _07988_;
 wire _07989_;
 wire _07990_;
 wire _07991_;
 wire _07992_;
 wire _07993_;
 wire _07994_;
 wire _07995_;
 wire _07996_;
 wire _07997_;
 wire _07998_;
 wire _07999_;
 wire _08000_;
 wire _08001_;
 wire _08002_;
 wire _08003_;
 wire _08004_;
 wire _08005_;
 wire _08006_;
 wire _08007_;
 wire _08008_;
 wire _08009_;
 wire _08010_;
 wire _08011_;
 wire _08012_;
 wire _08013_;
 wire _08014_;
 wire _08015_;
 wire _08016_;
 wire _08017_;
 wire _08018_;
 wire _08019_;
 wire _08020_;
 wire _08021_;
 wire _08022_;
 wire _08023_;
 wire _08024_;
 wire _08025_;
 wire _08026_;
 wire _08027_;
 wire _08028_;
 wire _08029_;
 wire _08030_;
 wire _08031_;
 wire _08032_;
 wire _08033_;
 wire _08034_;
 wire _08035_;
 wire _08036_;
 wire _08037_;
 wire _08038_;
 wire _08039_;
 wire _08040_;
 wire _08041_;
 wire _08042_;
 wire _08043_;
 wire _08044_;
 wire _08045_;
 wire _08046_;
 wire _08047_;
 wire _08048_;
 wire _08049_;
 wire _08050_;
 wire _08051_;
 wire _08052_;
 wire _08053_;
 wire _08054_;
 wire _08055_;
 wire _08056_;
 wire _08057_;
 wire _08058_;
 wire _08059_;
 wire _08060_;
 wire _08061_;
 wire _08062_;
 wire _08063_;
 wire _08064_;
 wire _08065_;
 wire _08066_;
 wire _08067_;
 wire _08068_;
 wire _08069_;
 wire _08070_;
 wire _08071_;
 wire _08072_;
 wire _08073_;
 wire _08074_;
 wire _08075_;
 wire _08076_;
 wire _08077_;
 wire _08078_;
 wire _08079_;
 wire _08080_;
 wire _08081_;
 wire _08082_;
 wire _08083_;
 wire _08084_;
 wire _08085_;
 wire _08086_;
 wire _08087_;
 wire _08088_;
 wire _08089_;
 wire _08090_;
 wire _08091_;
 wire _08092_;
 wire _08093_;
 wire _08094_;
 wire _08095_;
 wire _08096_;
 wire _08097_;
 wire _08098_;
 wire _08099_;
 wire _08100_;
 wire _08101_;
 wire _08102_;
 wire _08103_;
 wire _08104_;
 wire _08105_;
 wire _08106_;
 wire _08107_;
 wire _08108_;
 wire _08109_;
 wire _08110_;
 wire _08111_;
 wire _08112_;
 wire _08113_;
 wire _08114_;
 wire _08115_;
 wire _08116_;
 wire _08117_;
 wire _08118_;
 wire _08119_;
 wire _08120_;
 wire _08121_;
 wire _08122_;
 wire _08123_;
 wire _08124_;
 wire _08125_;
 wire _08126_;
 wire _08127_;
 wire _08128_;
 wire _08129_;
 wire _08130_;
 wire _08131_;
 wire _08132_;
 wire _08133_;
 wire _08134_;
 wire _08135_;
 wire _08136_;
 wire _08137_;
 wire _08138_;
 wire _08139_;
 wire _08140_;
 wire _08141_;
 wire _08142_;
 wire _08143_;
 wire _08144_;
 wire _08145_;
 wire _08146_;
 wire _08147_;
 wire _08148_;
 wire _08149_;
 wire _08150_;
 wire _08151_;
 wire _08152_;
 wire _08153_;
 wire _08154_;
 wire _08155_;
 wire _08156_;
 wire _08157_;
 wire _08158_;
 wire _08159_;
 wire _08160_;
 wire _08161_;
 wire _08162_;
 wire _08163_;
 wire _08164_;
 wire _08165_;
 wire _08166_;
 wire _08167_;
 wire _08168_;
 wire _08169_;
 wire _08170_;
 wire _08171_;
 wire _08172_;
 wire _08173_;
 wire _08174_;
 wire _08175_;
 wire _08176_;
 wire _08177_;
 wire _08178_;
 wire _08179_;
 wire _08180_;
 wire _08181_;
 wire _08182_;
 wire _08183_;
 wire _08184_;
 wire _08185_;
 wire _08186_;
 wire _08187_;
 wire _08188_;
 wire _08189_;
 wire _08190_;
 wire _08191_;
 wire _08192_;
 wire _08193_;
 wire _08194_;
 wire _08195_;
 wire _08196_;
 wire _08197_;
 wire _08198_;
 wire _08199_;
 wire _08200_;
 wire _08201_;
 wire _08202_;
 wire _08203_;
 wire _08204_;
 wire _08205_;
 wire _08206_;
 wire _08207_;
 wire _08208_;
 wire _08209_;
 wire _08210_;
 wire _08211_;
 wire _08212_;
 wire _08213_;
 wire _08214_;
 wire _08215_;
 wire _08216_;
 wire _08217_;
 wire _08218_;
 wire _08219_;
 wire _08220_;
 wire _08221_;
 wire _08222_;
 wire _08223_;
 wire _08224_;
 wire _08225_;
 wire _08226_;
 wire _08227_;
 wire _08228_;
 wire _08229_;
 wire _08230_;
 wire _08231_;
 wire _08232_;
 wire _08233_;
 wire _08234_;
 wire _08235_;
 wire _08236_;
 wire _08237_;
 wire _08238_;
 wire _08239_;
 wire _08240_;
 wire _08241_;
 wire _08242_;
 wire _08243_;
 wire _08244_;
 wire _08245_;
 wire _08246_;
 wire _08247_;
 wire _08248_;
 wire _08249_;
 wire _08250_;
 wire _08251_;
 wire _08252_;
 wire _08253_;
 wire _08254_;
 wire _08255_;
 wire _08256_;
 wire _08257_;
 wire _08258_;
 wire _08259_;
 wire _08260_;
 wire _08261_;
 wire _08262_;
 wire _08263_;
 wire _08264_;
 wire _08265_;
 wire _08266_;
 wire _08267_;
 wire _08268_;
 wire _08269_;
 wire _08270_;
 wire _08271_;
 wire _08272_;
 wire _08273_;
 wire _08274_;
 wire _08275_;
 wire _08276_;
 wire _08277_;
 wire _08278_;
 wire _08279_;
 wire _08280_;
 wire _08281_;
 wire _08282_;
 wire _08283_;
 wire _08284_;
 wire _08285_;
 wire _08286_;
 wire _08287_;
 wire _08288_;
 wire _08289_;
 wire _08290_;
 wire _08291_;
 wire _08292_;
 wire _08293_;
 wire _08294_;
 wire _08295_;
 wire _08296_;
 wire _08297_;
 wire _08298_;
 wire _08299_;
 wire _08300_;
 wire _08301_;
 wire _08302_;
 wire _08303_;
 wire _08304_;
 wire _08305_;
 wire _08306_;
 wire _08307_;
 wire _08308_;
 wire _08309_;
 wire _08310_;
 wire _08311_;
 wire _08312_;
 wire _08313_;
 wire _08314_;
 wire _08315_;
 wire _08316_;
 wire _08317_;
 wire _08318_;
 wire _08319_;
 wire _08320_;
 wire _08321_;
 wire _08322_;
 wire _08323_;
 wire _08324_;
 wire _08325_;
 wire _08326_;
 wire _08327_;
 wire _08328_;
 wire _08329_;
 wire _08330_;
 wire _08331_;
 wire _08332_;
 wire _08333_;
 wire _08334_;
 wire _08335_;
 wire _08336_;
 wire _08337_;
 wire _08338_;
 wire _08339_;
 wire _08340_;
 wire _08341_;
 wire _08342_;
 wire _08343_;
 wire _08344_;
 wire _08345_;
 wire _08346_;
 wire _08347_;
 wire _08348_;
 wire _08349_;
 wire _08350_;
 wire _08351_;
 wire _08352_;
 wire _08353_;
 wire _08354_;
 wire _08355_;
 wire _08356_;
 wire _08357_;
 wire _08358_;
 wire _08359_;
 wire _08360_;
 wire _08361_;
 wire _08362_;
 wire _08363_;
 wire _08364_;
 wire _08365_;
 wire _08366_;
 wire _08367_;
 wire _08368_;
 wire _08369_;
 wire _08370_;
 wire _08371_;
 wire _08372_;
 wire _08373_;
 wire _08374_;
 wire _08375_;
 wire _08376_;
 wire _08377_;
 wire _08378_;
 wire _08379_;
 wire _08380_;
 wire _08381_;
 wire _08382_;
 wire _08383_;
 wire _08384_;
 wire _08385_;
 wire _08386_;
 wire _08387_;
 wire _08388_;
 wire _08389_;
 wire _08390_;
 wire _08391_;
 wire _08392_;
 wire _08393_;
 wire _08394_;
 wire _08395_;
 wire _08396_;
 wire _08397_;
 wire _08398_;
 wire _08399_;
 wire _08400_;
 wire _08401_;
 wire _08402_;
 wire _08403_;
 wire _08404_;
 wire _08405_;
 wire _08406_;
 wire _08407_;
 wire _08408_;
 wire _08409_;
 wire _08410_;
 wire _08411_;
 wire _08412_;
 wire _08413_;
 wire _08414_;
 wire _08415_;
 wire _08416_;
 wire _08417_;
 wire _08418_;
 wire _08419_;
 wire _08420_;
 wire _08421_;
 wire _08422_;
 wire _08423_;
 wire _08424_;
 wire _08425_;
 wire _08426_;
 wire _08427_;
 wire _08428_;
 wire _08429_;
 wire _08430_;
 wire _08431_;
 wire _08432_;
 wire _08433_;
 wire _08434_;
 wire _08435_;
 wire _08436_;
 wire _08437_;
 wire _08438_;
 wire _08439_;
 wire _08440_;
 wire _08441_;
 wire _08442_;
 wire _08443_;
 wire _08444_;
 wire _08445_;
 wire _08446_;
 wire _08447_;
 wire _08448_;
 wire _08449_;
 wire _08450_;
 wire _08451_;
 wire _08452_;
 wire _08453_;
 wire _08454_;
 wire _08455_;
 wire _08456_;
 wire _08457_;
 wire _08458_;
 wire _08459_;
 wire _08460_;
 wire _08461_;
 wire _08462_;
 wire _08463_;
 wire _08464_;
 wire _08465_;
 wire _08466_;
 wire _08467_;
 wire _08468_;
 wire _08469_;
 wire _08470_;
 wire _08471_;
 wire _08472_;
 wire _08473_;
 wire _08474_;
 wire _08475_;
 wire _08476_;
 wire _08477_;
 wire _08478_;
 wire _08479_;
 wire _08480_;
 wire _08481_;
 wire _08482_;
 wire _08483_;
 wire _08484_;
 wire _08485_;
 wire _08486_;
 wire _08487_;
 wire _08488_;
 wire _08489_;
 wire _08490_;
 wire _08491_;
 wire _08492_;
 wire _08493_;
 wire _08494_;
 wire _08495_;
 wire _08496_;
 wire _08497_;
 wire _08498_;
 wire _08499_;
 wire _08500_;
 wire _08501_;
 wire _08502_;
 wire _08503_;
 wire _08504_;
 wire _08505_;
 wire _08506_;
 wire _08507_;
 wire _08508_;
 wire _08509_;
 wire _08510_;
 wire _08511_;
 wire _08512_;
 wire _08513_;
 wire _08514_;
 wire _08515_;
 wire _08516_;
 wire _08517_;
 wire _08518_;
 wire _08519_;
 wire _08520_;
 wire _08521_;
 wire _08522_;
 wire _08523_;
 wire _08524_;
 wire _08525_;
 wire _08526_;
 wire _08527_;
 wire _08528_;
 wire _08529_;
 wire _08530_;
 wire _08531_;
 wire _08532_;
 wire _08533_;
 wire _08534_;
 wire _08535_;
 wire _08536_;
 wire _08537_;
 wire _08538_;
 wire _08539_;
 wire _08540_;
 wire _08541_;
 wire _08542_;
 wire _08543_;
 wire _08544_;
 wire _08545_;
 wire _08546_;
 wire _08547_;
 wire _08548_;
 wire _08549_;
 wire _08550_;
 wire _08551_;
 wire _08552_;
 wire _08553_;
 wire _08554_;
 wire _08555_;
 wire _08556_;
 wire _08557_;
 wire _08558_;
 wire _08559_;
 wire _08560_;
 wire _08561_;
 wire _08562_;
 wire _08563_;
 wire _08564_;
 wire _08565_;
 wire _08566_;
 wire _08567_;
 wire _08568_;
 wire _08569_;
 wire _08570_;
 wire _08571_;
 wire _08572_;
 wire _08573_;
 wire _08574_;
 wire _08575_;
 wire _08576_;
 wire _08577_;
 wire _08578_;
 wire _08579_;
 wire _08580_;
 wire _08581_;
 wire _08582_;
 wire _08583_;
 wire _08584_;
 wire _08585_;
 wire _08586_;
 wire _08587_;
 wire _08588_;
 wire _08589_;
 wire _08590_;
 wire _08591_;
 wire _08592_;
 wire _08593_;
 wire _08594_;
 wire _08595_;
 wire _08596_;
 wire _08597_;
 wire _08598_;
 wire _08599_;
 wire _08600_;
 wire _08601_;
 wire _08602_;
 wire _08603_;
 wire _08604_;
 wire _08605_;
 wire _08606_;
 wire _08607_;
 wire _08608_;
 wire _08609_;
 wire _08610_;
 wire _08611_;
 wire _08612_;
 wire _08613_;
 wire _08614_;
 wire _08615_;
 wire _08616_;
 wire _08617_;
 wire _08618_;
 wire _08619_;
 wire _08620_;
 wire _08621_;
 wire _08622_;
 wire _08623_;
 wire _08624_;
 wire _08625_;
 wire _08626_;
 wire _08627_;
 wire _08628_;
 wire _08629_;
 wire _08630_;
 wire _08631_;
 wire _08632_;
 wire _08633_;
 wire _08634_;
 wire _08635_;
 wire _08636_;
 wire _08637_;
 wire _08638_;
 wire _08639_;
 wire _08640_;
 wire _08641_;
 wire _08642_;
 wire _08643_;
 wire _08644_;
 wire _08645_;
 wire _08646_;
 wire _08647_;
 wire _08648_;
 wire _08649_;
 wire _08650_;
 wire _08651_;
 wire _08652_;
 wire _08653_;
 wire _08654_;
 wire _08655_;
 wire _08656_;
 wire _08657_;
 wire _08658_;
 wire _08659_;
 wire _08660_;
 wire _08661_;
 wire _08662_;
 wire _08663_;
 wire _08664_;
 wire _08665_;
 wire _08666_;
 wire _08667_;
 wire _08668_;
 wire _08669_;
 wire _08670_;
 wire _08671_;
 wire _08672_;
 wire _08673_;
 wire _08674_;
 wire _08675_;
 wire _08676_;
 wire _08677_;
 wire _08678_;
 wire _08679_;
 wire _08680_;
 wire _08681_;
 wire _08682_;
 wire _08683_;
 wire _08684_;
 wire _08685_;
 wire _08686_;
 wire _08687_;
 wire _08688_;
 wire _08689_;
 wire _08690_;
 wire _08691_;
 wire _08692_;
 wire _08693_;
 wire _08694_;
 wire _08695_;
 wire _08696_;
 wire _08697_;
 wire _08698_;
 wire _08699_;
 wire _08700_;
 wire _08701_;
 wire _08702_;
 wire _08703_;
 wire _08704_;
 wire _08705_;
 wire _08706_;
 wire _08707_;
 wire _08708_;
 wire _08709_;
 wire _08710_;
 wire _08711_;
 wire _08712_;
 wire _08713_;
 wire _08714_;
 wire _08715_;
 wire _08716_;
 wire _08717_;
 wire _08718_;
 wire _08719_;
 wire _08720_;
 wire _08721_;
 wire _08722_;
 wire _08723_;
 wire _08724_;
 wire _08725_;
 wire _08726_;
 wire _08727_;
 wire _08728_;
 wire _08729_;
 wire _08730_;
 wire _08731_;
 wire _08732_;
 wire _08733_;
 wire _08734_;
 wire _08735_;
 wire _08736_;
 wire _08737_;
 wire _08738_;
 wire _08739_;
 wire _08740_;
 wire _08741_;
 wire _08742_;
 wire _08743_;
 wire _08744_;
 wire _08745_;
 wire _08746_;
 wire _08747_;
 wire _08748_;
 wire _08749_;
 wire _08750_;
 wire _08751_;
 wire _08752_;
 wire _08753_;
 wire _08754_;
 wire _08755_;
 wire _08756_;
 wire _08757_;
 wire _08758_;
 wire _08759_;
 wire _08760_;
 wire _08761_;
 wire _08762_;
 wire _08763_;
 wire _08764_;
 wire _08765_;
 wire _08766_;
 wire _08767_;
 wire _08768_;
 wire _08769_;
 wire _08770_;
 wire _08771_;
 wire _08772_;
 wire _08773_;
 wire _08774_;
 wire _08775_;
 wire _08776_;
 wire _08777_;
 wire _08778_;
 wire _08779_;
 wire _08780_;
 wire _08781_;
 wire _08782_;
 wire _08783_;
 wire _08784_;
 wire _08785_;
 wire _08786_;
 wire _08787_;
 wire _08788_;
 wire _08789_;
 wire _08790_;
 wire _08791_;
 wire _08792_;
 wire _08793_;
 wire _08794_;
 wire _08795_;
 wire _08796_;
 wire _08797_;
 wire _08798_;
 wire _08799_;
 wire _08800_;
 wire _08801_;
 wire _08802_;
 wire _08803_;
 wire _08804_;
 wire _08805_;
 wire _08806_;
 wire _08807_;
 wire _08808_;
 wire _08809_;
 wire _08810_;
 wire _08811_;
 wire _08812_;
 wire _08813_;
 wire _08814_;
 wire _08815_;
 wire _08816_;
 wire _08817_;
 wire _08818_;
 wire _08819_;
 wire _08820_;
 wire _08821_;
 wire _08822_;
 wire _08823_;
 wire _08824_;
 wire _08825_;
 wire _08826_;
 wire _08827_;
 wire _08828_;
 wire _08829_;
 wire _08830_;
 wire _08831_;
 wire _08832_;
 wire _08833_;
 wire _08834_;
 wire _08835_;
 wire _08836_;
 wire _08837_;
 wire _08838_;
 wire _08839_;
 wire _08840_;
 wire _08841_;
 wire _08842_;
 wire _08843_;
 wire _08844_;
 wire _08845_;
 wire _08846_;
 wire _08847_;
 wire _08848_;
 wire _08849_;
 wire _08850_;
 wire _08851_;
 wire _08852_;
 wire _08853_;
 wire _08854_;
 wire _08855_;
 wire _08856_;
 wire _08857_;
 wire _08858_;
 wire _08859_;
 wire _08860_;
 wire _08861_;
 wire _08862_;
 wire _08863_;
 wire _08864_;
 wire _08865_;
 wire _08866_;
 wire _08867_;
 wire _08868_;
 wire _08869_;
 wire _08870_;
 wire _08871_;
 wire _08872_;
 wire _08873_;
 wire _08874_;
 wire _08875_;
 wire _08876_;
 wire _08877_;
 wire _08878_;
 wire _08879_;
 wire _08880_;
 wire _08881_;
 wire _08882_;
 wire _08883_;
 wire _08884_;
 wire _08885_;
 wire _08886_;
 wire _08887_;
 wire _08888_;
 wire _08889_;
 wire _08890_;
 wire _08891_;
 wire _08892_;
 wire _08893_;
 wire _08894_;
 wire _08895_;
 wire _08896_;
 wire _08897_;
 wire _08898_;
 wire _08899_;
 wire _08900_;
 wire _08901_;
 wire _08902_;
 wire _08903_;
 wire _08904_;
 wire _08905_;
 wire _08906_;
 wire _08907_;
 wire _08908_;
 wire _08909_;
 wire _08910_;
 wire _08911_;
 wire _08912_;
 wire _08913_;
 wire _08914_;
 wire _08915_;
 wire _08916_;
 wire _08917_;
 wire _08918_;
 wire _08919_;
 wire _08920_;
 wire _08921_;
 wire _08922_;
 wire _08923_;
 wire _08924_;
 wire _08925_;
 wire _08926_;
 wire _08927_;
 wire _08928_;
 wire _08929_;
 wire _08930_;
 wire _08931_;
 wire _08932_;
 wire _08933_;
 wire _08934_;
 wire _08935_;
 wire _08936_;
 wire _08937_;
 wire _08938_;
 wire _08939_;
 wire _08940_;
 wire _08941_;
 wire _08942_;
 wire _08943_;
 wire _08944_;
 wire _08945_;
 wire _08946_;
 wire _08947_;
 wire _08948_;
 wire _08949_;
 wire _08950_;
 wire _08951_;
 wire _08952_;
 wire _08953_;
 wire _08954_;
 wire _08955_;
 wire _08956_;
 wire _08957_;
 wire _08958_;
 wire _08959_;
 wire _08960_;
 wire _08961_;
 wire _08962_;
 wire _08963_;
 wire _08964_;
 wire _08965_;
 wire _08966_;
 wire _08967_;
 wire _08968_;
 wire _08969_;
 wire _08970_;
 wire _08971_;
 wire _08972_;
 wire _08973_;
 wire _08974_;
 wire _08975_;
 wire _08976_;
 wire _08977_;
 wire _08978_;
 wire _08979_;
 wire _08980_;
 wire _08981_;
 wire _08982_;
 wire _08983_;
 wire _08984_;
 wire _08985_;
 wire _08986_;
 wire _08987_;
 wire _08988_;
 wire _08989_;
 wire _08990_;
 wire _08991_;
 wire _08992_;
 wire _08993_;
 wire _08994_;
 wire _08995_;
 wire _08996_;
 wire _08997_;
 wire _08998_;
 wire _08999_;
 wire _09000_;
 wire _09001_;
 wire _09002_;
 wire _09003_;
 wire _09004_;
 wire _09005_;
 wire _09006_;
 wire _09007_;
 wire _09008_;
 wire _09009_;
 wire _09010_;
 wire _09011_;
 wire _09012_;
 wire _09013_;
 wire _09014_;
 wire _09015_;
 wire _09016_;
 wire _09017_;
 wire _09018_;
 wire _09019_;
 wire _09020_;
 wire _09021_;
 wire _09022_;
 wire _09023_;
 wire _09024_;
 wire _09025_;
 wire _09026_;
 wire _09027_;
 wire _09028_;
 wire _09029_;
 wire _09030_;
 wire _09031_;
 wire _09032_;
 wire _09033_;
 wire _09034_;
 wire _09035_;
 wire _09036_;
 wire _09037_;
 wire _09038_;
 wire _09039_;
 wire _09040_;
 wire _09041_;
 wire _09042_;
 wire _09043_;
 wire _09044_;
 wire _09045_;
 wire _09046_;
 wire _09047_;
 wire _09048_;
 wire _09049_;
 wire _09050_;
 wire _09051_;
 wire _09052_;
 wire _09053_;
 wire _09054_;
 wire _09055_;
 wire _09056_;
 wire _09057_;
 wire _09058_;
 wire _09059_;
 wire _09060_;
 wire _09061_;
 wire _09062_;
 wire _09063_;
 wire _09064_;
 wire _09065_;
 wire _09066_;
 wire _09067_;
 wire _09068_;
 wire _09069_;
 wire _09070_;
 wire _09071_;
 wire _09072_;
 wire _09073_;
 wire _09074_;
 wire _09075_;
 wire _09076_;
 wire _09077_;
 wire _09078_;
 wire _09079_;
 wire _09080_;
 wire _09081_;
 wire _09082_;
 wire _09083_;
 wire _09084_;
 wire _09085_;
 wire _09086_;
 wire _09087_;
 wire _09088_;
 wire _09089_;
 wire _09090_;
 wire _09091_;
 wire _09092_;
 wire _09093_;
 wire _09094_;
 wire _09095_;
 wire _09096_;
 wire _09097_;
 wire _09098_;
 wire _09099_;
 wire _09100_;
 wire _09101_;
 wire _09102_;
 wire _09103_;
 wire _09104_;
 wire _09105_;
 wire _09106_;
 wire _09107_;
 wire _09108_;
 wire _09109_;
 wire _09110_;
 wire _09111_;
 wire _09112_;
 wire _09113_;
 wire _09114_;
 wire _09115_;
 wire _09116_;
 wire _09117_;
 wire _09118_;
 wire _09119_;
 wire _09120_;
 wire _09121_;
 wire _09122_;
 wire _09123_;
 wire _09124_;
 wire _09125_;
 wire _09126_;
 wire _09127_;
 wire _09128_;
 wire _09129_;
 wire _09130_;
 wire _09131_;
 wire _09132_;
 wire _09133_;
 wire _09134_;
 wire _09135_;
 wire _09136_;
 wire _09137_;
 wire _09138_;
 wire _09139_;
 wire _09140_;
 wire _09141_;
 wire _09142_;
 wire _09143_;
 wire _09144_;
 wire _09145_;
 wire _09146_;
 wire _09147_;
 wire _09148_;
 wire _09149_;
 wire _09150_;
 wire _09151_;
 wire _09152_;
 wire _09153_;
 wire _09154_;
 wire _09155_;
 wire _09156_;
 wire _09157_;
 wire _09158_;
 wire _09159_;
 wire _09160_;
 wire _09161_;
 wire _09162_;
 wire _09163_;
 wire _09164_;
 wire _09165_;
 wire _09166_;
 wire _09167_;
 wire _09168_;
 wire _09169_;
 wire _09170_;
 wire _09171_;
 wire _09172_;
 wire _09173_;
 wire _09174_;
 wire _09175_;
 wire _09176_;
 wire _09177_;
 wire _09178_;
 wire _09179_;
 wire _09180_;
 wire _09181_;
 wire _09182_;
 wire _09183_;
 wire _09184_;
 wire _09185_;
 wire _09186_;
 wire _09187_;
 wire _09188_;
 wire _09189_;
 wire _09190_;
 wire _09191_;
 wire _09192_;
 wire _09193_;
 wire _09194_;
 wire _09195_;
 wire _09196_;
 wire _09197_;
 wire _09198_;
 wire _09199_;
 wire _09200_;
 wire _09201_;
 wire _09202_;
 wire _09203_;
 wire _09204_;
 wire _09205_;
 wire _09206_;
 wire _09207_;
 wire _09208_;
 wire _09209_;
 wire _09210_;
 wire _09211_;
 wire _09212_;
 wire _09213_;
 wire _09214_;
 wire _09215_;
 wire _09216_;
 wire _09217_;
 wire _09218_;
 wire _09219_;
 wire _09220_;
 wire _09221_;
 wire _09222_;
 wire _09223_;
 wire _09224_;
 wire _09225_;
 wire _09226_;
 wire _09227_;
 wire _09228_;
 wire _09229_;
 wire _09230_;
 wire _09231_;
 wire _09232_;
 wire _09233_;
 wire _09234_;
 wire _09235_;
 wire _09236_;
 wire _09237_;
 wire _09238_;
 wire _09239_;
 wire _09240_;
 wire _09241_;
 wire _09242_;
 wire _09243_;
 wire _09244_;
 wire _09245_;
 wire _09246_;
 wire _09247_;
 wire _09248_;
 wire _09249_;
 wire _09250_;
 wire _09251_;
 wire _09252_;
 wire _09253_;
 wire _09254_;
 wire _09255_;
 wire _09256_;
 wire _09257_;
 wire _09258_;
 wire _09259_;
 wire _09260_;
 wire _09261_;
 wire _09262_;
 wire _09263_;
 wire _09264_;
 wire _09265_;
 wire _09266_;
 wire _09267_;
 wire _09268_;
 wire _09269_;
 wire _09270_;
 wire _09271_;
 wire _09272_;
 wire _09273_;
 wire _09274_;
 wire _09275_;
 wire _09276_;
 wire _09277_;
 wire _09278_;
 wire _09279_;
 wire _09280_;
 wire _09281_;
 wire _09282_;
 wire _09283_;
 wire _09284_;
 wire _09285_;
 wire _09286_;
 wire _09287_;
 wire _09288_;
 wire _09289_;
 wire _09290_;
 wire _09291_;
 wire _09292_;
 wire _09293_;
 wire _09294_;
 wire _09295_;
 wire _09296_;
 wire _09297_;
 wire _09298_;
 wire _09299_;
 wire _09300_;
 wire _09301_;
 wire _09302_;
 wire _09303_;
 wire _09304_;
 wire _09305_;
 wire _09306_;
 wire _09307_;
 wire _09308_;
 wire _09309_;
 wire _09310_;
 wire _09311_;
 wire _09312_;
 wire _09313_;
 wire _09314_;
 wire _09315_;
 wire _09316_;
 wire _09317_;
 wire _09318_;
 wire _09319_;
 wire _09320_;
 wire _09321_;
 wire _09322_;
 wire _09323_;
 wire _09324_;
 wire _09325_;
 wire _09326_;
 wire _09327_;
 wire _09328_;
 wire _09329_;
 wire _09330_;
 wire _09331_;
 wire _09332_;
 wire _09333_;
 wire _09334_;
 wire _09335_;
 wire _09336_;
 wire _09337_;
 wire _09338_;
 wire _09339_;
 wire _09340_;
 wire _09341_;
 wire _09342_;
 wire _09343_;
 wire _09344_;
 wire _09345_;
 wire _09346_;
 wire _09347_;
 wire _09348_;
 wire _09349_;
 wire _09350_;
 wire _09351_;
 wire _09352_;
 wire _09353_;
 wire _09354_;
 wire _09355_;
 wire _09356_;
 wire _09357_;
 wire _09358_;
 wire _09359_;
 wire _09360_;
 wire _09361_;
 wire _09362_;
 wire _09363_;
 wire _09364_;
 wire _09365_;
 wire _09366_;
 wire _09367_;
 wire _09368_;
 wire _09369_;
 wire _09370_;
 wire _09371_;
 wire _09372_;
 wire _09373_;
 wire _09374_;
 wire _09375_;
 wire _09376_;
 wire _09377_;
 wire _09378_;
 wire _09379_;
 wire _09380_;
 wire _09381_;
 wire _09382_;
 wire _09383_;
 wire _09384_;
 wire _09385_;
 wire _09386_;
 wire _09387_;
 wire _09388_;
 wire _09389_;
 wire _09390_;
 wire _09391_;
 wire _09392_;
 wire _09393_;
 wire _09394_;
 wire _09395_;
 wire _09396_;
 wire _09397_;
 wire _09398_;
 wire _09399_;
 wire _09400_;
 wire _09401_;
 wire _09402_;
 wire _09403_;
 wire _09404_;
 wire _09405_;
 wire _09406_;
 wire _09407_;
 wire _09408_;
 wire _09409_;
 wire _09410_;
 wire _09411_;
 wire _09412_;
 wire _09413_;
 wire _09414_;
 wire _09415_;
 wire _09416_;
 wire _09417_;
 wire _09418_;
 wire _09419_;
 wire _09420_;
 wire _09421_;
 wire _09422_;
 wire _09423_;
 wire _09424_;
 wire _09425_;
 wire _09426_;
 wire _09427_;
 wire _09428_;
 wire _09429_;
 wire _09430_;
 wire _09431_;
 wire _09432_;
 wire _09433_;
 wire _09434_;
 wire _09435_;
 wire _09436_;
 wire _09437_;
 wire _09438_;
 wire _09439_;
 wire _09440_;
 wire _09441_;
 wire _09442_;
 wire _09443_;
 wire _09444_;
 wire _09445_;
 wire _09446_;
 wire _09447_;
 wire _09448_;
 wire _09449_;
 wire _09450_;
 wire _09451_;
 wire _09452_;
 wire _09453_;
 wire _09454_;
 wire _09455_;
 wire _09456_;
 wire _09457_;
 wire _09458_;
 wire _09459_;
 wire _09460_;
 wire _09461_;
 wire _09462_;
 wire _09463_;
 wire _09464_;
 wire _09465_;
 wire _09466_;
 wire _09467_;
 wire _09468_;
 wire _09469_;
 wire _09470_;
 wire _09471_;
 wire _09472_;
 wire _09473_;
 wire _09474_;
 wire _09475_;
 wire _09476_;
 wire _09477_;
 wire _09478_;
 wire _09479_;
 wire _09480_;
 wire _09481_;
 wire _09482_;
 wire _09483_;
 wire _09484_;
 wire _09485_;
 wire _09486_;
 wire _09487_;
 wire _09488_;
 wire _09489_;
 wire _09490_;
 wire _09491_;
 wire _09492_;
 wire _09493_;
 wire _09494_;
 wire _09495_;
 wire _09496_;
 wire _09497_;
 wire _09498_;
 wire _09499_;
 wire _09500_;
 wire _09501_;
 wire _09502_;
 wire _09503_;
 wire _09504_;
 wire _09505_;
 wire _09506_;
 wire _09507_;
 wire _09508_;
 wire _09509_;
 wire _09510_;
 wire _09511_;
 wire _09512_;
 wire _09513_;
 wire _09514_;
 wire _09515_;
 wire _09516_;
 wire _09517_;
 wire _09518_;
 wire _09519_;
 wire _09520_;
 wire _09521_;
 wire _09522_;
 wire _09523_;
 wire _09524_;
 wire _09525_;
 wire _09526_;
 wire _09527_;
 wire _09528_;
 wire _09529_;
 wire _09530_;
 wire _09531_;
 wire _09532_;
 wire _09533_;
 wire _09534_;
 wire _09535_;
 wire _09536_;
 wire _09537_;
 wire _09538_;
 wire _09539_;
 wire _09540_;
 wire _09541_;
 wire _09542_;
 wire _09543_;
 wire _09544_;
 wire _09545_;
 wire _09546_;
 wire _09547_;
 wire _09548_;
 wire _09549_;
 wire _09550_;
 wire _09551_;
 wire _09552_;
 wire _09553_;
 wire _09554_;
 wire _09555_;
 wire _09556_;
 wire _09557_;
 wire _09558_;
 wire _09559_;
 wire _09560_;
 wire _09561_;
 wire _09562_;
 wire _09563_;
 wire _09564_;
 wire _09565_;
 wire _09566_;
 wire _09567_;
 wire _09568_;
 wire _09569_;
 wire _09570_;
 wire _09571_;
 wire _09572_;
 wire _09573_;
 wire _09574_;
 wire _09575_;
 wire _09576_;
 wire _09577_;
 wire _09578_;
 wire _09579_;
 wire _09580_;
 wire _09581_;
 wire _09582_;
 wire _09583_;
 wire _09584_;
 wire _09585_;
 wire _09586_;
 wire _09587_;
 wire _09588_;
 wire _09589_;
 wire _09590_;
 wire _09591_;
 wire _09592_;
 wire _09593_;
 wire _09594_;
 wire _09595_;
 wire _09596_;
 wire _09597_;
 wire _09598_;
 wire _09599_;
 wire _09600_;
 wire _09601_;
 wire _09602_;
 wire _09603_;
 wire _09604_;
 wire _09605_;
 wire _09606_;
 wire _09607_;
 wire _09608_;
 wire _09609_;
 wire _09610_;
 wire _09611_;
 wire _09612_;
 wire _09613_;
 wire _09614_;
 wire _09615_;
 wire _09616_;
 wire _09617_;
 wire _09618_;
 wire _09619_;
 wire _09620_;
 wire _09621_;
 wire _09622_;
 wire _09623_;
 wire _09624_;
 wire _09625_;
 wire _09626_;
 wire _09627_;
 wire _09628_;
 wire _09629_;
 wire _09630_;
 wire _09631_;
 wire _09632_;
 wire _09633_;
 wire _09634_;
 wire _09635_;
 wire _09636_;
 wire _09637_;
 wire _09638_;
 wire _09639_;
 wire _09640_;
 wire _09641_;
 wire _09642_;
 wire _09643_;
 wire _09644_;
 wire _09645_;
 wire _09646_;
 wire _09647_;
 wire _09648_;
 wire _09649_;
 wire _09650_;
 wire _09651_;
 wire _09652_;
 wire _09653_;
 wire _09654_;
 wire _09655_;
 wire _09656_;
 wire _09657_;
 wire _09658_;
 wire _09659_;
 wire _09660_;
 wire _09661_;
 wire _09662_;
 wire _09663_;
 wire _09664_;
 wire _09665_;
 wire _09666_;
 wire _09667_;
 wire _09668_;
 wire _09669_;
 wire _09670_;
 wire _09671_;
 wire _09672_;
 wire _09673_;
 wire _09674_;
 wire _09675_;
 wire _09676_;
 wire _09677_;
 wire _09678_;
 wire _09679_;
 wire _09680_;
 wire _09681_;
 wire _09682_;
 wire _09683_;
 wire _09684_;
 wire _09685_;
 wire _09686_;
 wire _09687_;
 wire _09688_;
 wire _09689_;
 wire _09690_;
 wire _09691_;
 wire _09692_;
 wire _09693_;
 wire _09694_;
 wire _09695_;
 wire _09696_;
 wire _09697_;
 wire _09698_;
 wire _09699_;
 wire _09700_;
 wire _09701_;
 wire _09702_;
 wire _09703_;
 wire _09704_;
 wire _09705_;
 wire _09706_;
 wire _09707_;
 wire _09708_;
 wire _09709_;
 wire _09710_;
 wire _09711_;
 wire _09712_;
 wire _09713_;
 wire _09714_;
 wire _09715_;
 wire _09716_;
 wire _09717_;
 wire _09718_;
 wire _09719_;
 wire _09720_;
 wire _09721_;
 wire _09722_;
 wire _09723_;
 wire _09724_;
 wire _09725_;
 wire _09726_;
 wire _09727_;
 wire _09728_;
 wire _09729_;
 wire _09730_;
 wire _09731_;
 wire _09732_;
 wire _09733_;
 wire _09734_;
 wire _09735_;
 wire _09736_;
 wire _09737_;
 wire _09738_;
 wire _09739_;
 wire _09740_;
 wire _09741_;
 wire _09742_;
 wire _09743_;
 wire _09744_;
 wire _09745_;
 wire _09746_;
 wire _09747_;
 wire _09748_;
 wire _09749_;
 wire _09750_;
 wire _09751_;
 wire _09752_;
 wire _09753_;
 wire _09754_;
 wire _09755_;
 wire _09756_;
 wire _09757_;
 wire _09758_;
 wire _09759_;
 wire _09760_;
 wire _09761_;
 wire _09762_;
 wire _09763_;
 wire _09764_;
 wire _09765_;
 wire _09766_;
 wire _09767_;
 wire _09768_;
 wire _09769_;
 wire _09770_;
 wire _09771_;
 wire _09772_;
 wire _09773_;
 wire _09774_;
 wire _09775_;
 wire _09776_;
 wire _09777_;
 wire _09778_;
 wire _09779_;
 wire _09780_;
 wire _09781_;
 wire _09782_;
 wire _09783_;
 wire _09784_;
 wire _09785_;
 wire _09786_;
 wire _09787_;
 wire _09788_;
 wire _09789_;
 wire _09790_;
 wire _09791_;
 wire _09792_;
 wire _09793_;
 wire _09794_;
 wire _09795_;
 wire _09796_;
 wire _09797_;
 wire _09798_;
 wire _09799_;
 wire _09800_;
 wire _09801_;
 wire _09802_;
 wire _09803_;
 wire _09804_;
 wire _09805_;
 wire _09806_;
 wire _09807_;
 wire _09808_;
 wire _09809_;
 wire _09810_;
 wire _09811_;
 wire _09812_;
 wire _09813_;
 wire _09814_;
 wire _09815_;
 wire _09816_;
 wire _09817_;
 wire _09818_;
 wire _09819_;
 wire _09820_;
 wire _09821_;
 wire _09822_;
 wire _09823_;
 wire _09824_;
 wire _09825_;
 wire _09826_;
 wire _09827_;
 wire _09828_;
 wire _09829_;
 wire _09830_;
 wire _09831_;
 wire _09832_;
 wire _09833_;
 wire _09834_;
 wire _09835_;
 wire _09836_;
 wire _09837_;
 wire _09838_;
 wire _09839_;
 wire _09840_;
 wire _09841_;
 wire _09842_;
 wire _09843_;
 wire _09844_;
 wire _09845_;
 wire _09846_;
 wire _09847_;
 wire _09848_;
 wire _09849_;
 wire _09850_;
 wire _09851_;
 wire _09852_;
 wire _09853_;
 wire _09854_;
 wire _09855_;
 wire _09856_;
 wire _09857_;
 wire _09858_;
 wire _09859_;
 wire _09860_;
 wire _09861_;
 wire _09862_;
 wire _09863_;
 wire _09864_;
 wire _09865_;
 wire _09866_;
 wire _09867_;
 wire _09868_;
 wire _09869_;
 wire _09870_;
 wire _09871_;
 wire _09872_;
 wire _09873_;
 wire _09874_;
 wire _09875_;
 wire _09876_;
 wire _09877_;
 wire _09878_;
 wire _09879_;
 wire _09880_;
 wire _09881_;
 wire _09882_;
 wire _09883_;
 wire _09884_;
 wire _09885_;
 wire _09886_;
 wire _09887_;
 wire _09888_;
 wire _09889_;
 wire _09890_;
 wire _09891_;
 wire _09892_;
 wire _09893_;
 wire _09894_;
 wire _09895_;
 wire _09896_;
 wire _09897_;
 wire _09898_;
 wire _09899_;
 wire _09900_;
 wire _09901_;
 wire _09902_;
 wire _09903_;
 wire _09904_;
 wire _09905_;
 wire _09906_;
 wire _09907_;
 wire _09908_;
 wire _09909_;
 wire _09910_;
 wire _09911_;
 wire _09912_;
 wire _09913_;
 wire _09914_;
 wire _09915_;
 wire _09916_;
 wire _09917_;
 wire _09918_;
 wire _09919_;
 wire _09920_;
 wire _09921_;
 wire _09922_;
 wire _09923_;
 wire _09924_;
 wire _09925_;
 wire _09926_;
 wire _09927_;
 wire _09928_;
 wire _09929_;
 wire _09930_;
 wire _09931_;
 wire _09932_;
 wire _09933_;
 wire _09934_;
 wire _09935_;
 wire _09936_;
 wire _09937_;
 wire _09938_;
 wire _09939_;
 wire _09940_;
 wire _09941_;
 wire _09942_;
 wire _09943_;
 wire _09944_;
 wire _09945_;
 wire _09946_;
 wire _09947_;
 wire _09948_;
 wire _09949_;
 wire _09950_;
 wire _09951_;
 wire _09952_;
 wire _09953_;
 wire _09954_;
 wire _09955_;
 wire _09956_;
 wire _09957_;
 wire _09958_;
 wire _09959_;
 wire _09960_;
 wire _09961_;
 wire _09962_;
 wire _09963_;
 wire _09964_;
 wire _09965_;
 wire _09966_;
 wire _09967_;
 wire _09968_;
 wire _09969_;
 wire _09970_;
 wire _09971_;
 wire _09972_;
 wire _09973_;
 wire _09974_;
 wire _09975_;
 wire _09976_;
 wire _09977_;
 wire _09978_;
 wire _09979_;
 wire _09980_;
 wire _09981_;
 wire _09982_;
 wire _09983_;
 wire _09984_;
 wire _09985_;
 wire _09986_;
 wire _09987_;
 wire _09988_;
 wire _09989_;
 wire _09990_;
 wire _09991_;
 wire _09992_;
 wire _09993_;
 wire _09994_;
 wire _09995_;
 wire _09996_;
 wire _09997_;
 wire _09998_;
 wire _09999_;
 wire _10000_;
 wire _10001_;
 wire _10002_;
 wire _10003_;
 wire _10004_;
 wire _10005_;
 wire _10006_;
 wire _10007_;
 wire _10008_;
 wire _10009_;
 wire _10010_;
 wire _10011_;
 wire _10012_;
 wire _10013_;
 wire _10014_;
 wire _10015_;
 wire _10016_;
 wire _10017_;
 wire _10018_;
 wire _10019_;
 wire _10020_;
 wire _10021_;
 wire _10022_;
 wire _10023_;
 wire _10024_;
 wire _10025_;
 wire _10026_;
 wire _10027_;
 wire _10028_;
 wire _10029_;
 wire _10030_;
 wire _10031_;
 wire _10032_;
 wire _10033_;
 wire _10034_;
 wire _10035_;
 wire _10036_;
 wire _10037_;
 wire _10038_;
 wire _10039_;
 wire _10040_;
 wire _10041_;
 wire _10042_;
 wire _10043_;
 wire _10044_;
 wire _10045_;
 wire _10046_;
 wire _10047_;
 wire _10048_;
 wire _10049_;
 wire _10050_;
 wire _10051_;
 wire _10052_;
 wire _10053_;
 wire _10054_;
 wire _10055_;
 wire _10056_;
 wire _10057_;
 wire _10058_;
 wire _10059_;
 wire _10060_;
 wire _10061_;
 wire _10062_;
 wire _10063_;
 wire _10064_;
 wire _10065_;
 wire _10066_;
 wire _10067_;
 wire _10068_;
 wire _10069_;
 wire _10070_;
 wire _10071_;
 wire _10072_;
 wire _10073_;
 wire _10074_;
 wire _10075_;
 wire _10076_;
 wire _10077_;
 wire _10078_;
 wire _10079_;
 wire _10080_;
 wire _10081_;
 wire _10082_;
 wire _10083_;
 wire _10084_;
 wire _10085_;
 wire _10086_;
 wire _10087_;
 wire _10088_;
 wire _10089_;
 wire _10090_;
 wire _10091_;
 wire _10092_;
 wire _10093_;
 wire _10094_;
 wire _10095_;
 wire _10096_;
 wire _10097_;
 wire _10098_;
 wire _10099_;
 wire _10100_;
 wire _10101_;
 wire _10102_;
 wire _10103_;
 wire _10104_;
 wire _10105_;
 wire _10106_;
 wire _10107_;
 wire _10108_;
 wire _10109_;
 wire _10110_;
 wire _10111_;
 wire _10112_;
 wire _10113_;
 wire _10114_;
 wire _10115_;
 wire _10116_;
 wire _10117_;
 wire _10118_;
 wire _10119_;
 wire _10120_;
 wire _10121_;
 wire _10122_;
 wire _10123_;
 wire _10124_;
 wire _10125_;
 wire _10126_;
 wire _10127_;
 wire _10128_;
 wire _10129_;
 wire _10130_;
 wire _10131_;
 wire _10132_;
 wire _10133_;
 wire _10134_;
 wire _10135_;
 wire _10136_;
 wire _10137_;
 wire _10138_;
 wire _10139_;
 wire _10140_;
 wire _10141_;
 wire _10142_;
 wire _10143_;
 wire _10144_;
 wire _10145_;
 wire _10146_;
 wire _10147_;
 wire _10148_;
 wire _10149_;
 wire _10150_;
 wire _10151_;
 wire _10152_;
 wire _10153_;
 wire _10154_;
 wire _10155_;
 wire _10156_;
 wire _10157_;
 wire _10158_;
 wire _10159_;
 wire _10160_;
 wire _10161_;
 wire _10162_;
 wire _10163_;
 wire _10164_;
 wire _10165_;
 wire _10166_;
 wire _10167_;
 wire _10168_;
 wire _10169_;
 wire _10170_;
 wire _10171_;
 wire _10172_;
 wire _10173_;
 wire _10174_;
 wire _10175_;
 wire _10176_;
 wire _10177_;
 wire _10178_;
 wire _10179_;
 wire _10180_;
 wire _10181_;
 wire _10182_;
 wire _10183_;
 wire _10184_;
 wire _10185_;
 wire _10186_;
 wire _10187_;
 wire _10188_;
 wire _10189_;
 wire _10190_;
 wire _10191_;
 wire _10192_;
 wire _10193_;
 wire _10194_;
 wire _10195_;
 wire _10196_;
 wire _10197_;
 wire _10198_;
 wire _10199_;
 wire _10200_;
 wire _10201_;
 wire _10202_;
 wire _10203_;
 wire _10204_;
 wire _10205_;
 wire _10206_;
 wire _10207_;
 wire _10208_;
 wire _10209_;
 wire _10210_;
 wire _10211_;
 wire _10212_;
 wire _10213_;
 wire _10214_;
 wire _10215_;
 wire _10216_;
 wire _10217_;
 wire _10218_;
 wire _10219_;
 wire _10220_;
 wire _10221_;
 wire _10222_;
 wire _10223_;
 wire _10224_;
 wire _10225_;
 wire _10226_;
 wire _10227_;
 wire _10228_;
 wire _10229_;
 wire _10230_;
 wire _10231_;
 wire _10232_;
 wire _10233_;
 wire _10234_;
 wire _10235_;
 wire _10236_;
 wire _10237_;
 wire _10238_;
 wire _10239_;
 wire _10240_;
 wire _10241_;
 wire _10242_;
 wire _10243_;
 wire _10244_;
 wire _10245_;
 wire _10246_;
 wire _10247_;
 wire _10248_;
 wire _10249_;
 wire _10250_;
 wire _10251_;
 wire _10252_;
 wire _10253_;
 wire _10254_;
 wire _10255_;
 wire _10256_;
 wire _10257_;
 wire _10258_;
 wire _10259_;
 wire _10260_;
 wire _10261_;
 wire _10262_;
 wire _10263_;
 wire _10264_;
 wire _10265_;
 wire _10266_;
 wire _10267_;
 wire _10268_;
 wire _10269_;
 wire _10270_;
 wire _10271_;
 wire _10272_;
 wire _10273_;
 wire _10274_;
 wire _10275_;
 wire _10276_;
 wire _10277_;
 wire _10278_;
 wire _10279_;
 wire _10280_;
 wire _10281_;
 wire _10282_;
 wire _10283_;
 wire _10284_;
 wire _10285_;
 wire _10286_;
 wire _10287_;
 wire _10288_;
 wire _10289_;
 wire _10290_;
 wire _10291_;
 wire _10292_;
 wire _10293_;
 wire _10294_;
 wire _10295_;
 wire _10296_;
 wire _10297_;
 wire _10298_;
 wire _10299_;
 wire _10300_;
 wire _10301_;
 wire _10302_;
 wire _10303_;
 wire _10304_;
 wire _10305_;
 wire _10306_;
 wire _10307_;
 wire _10308_;
 wire _10309_;
 wire _10310_;
 wire _10311_;
 wire _10312_;
 wire _10313_;
 wire _10314_;
 wire _10315_;
 wire _10316_;
 wire _10317_;
 wire _10318_;
 wire _10319_;
 wire _10320_;
 wire _10321_;
 wire _10322_;
 wire _10323_;
 wire _10324_;
 wire _10325_;
 wire _10326_;
 wire _10327_;
 wire _10328_;
 wire _10329_;
 wire _10330_;
 wire _10331_;
 wire _10332_;
 wire _10333_;
 wire _10334_;
 wire _10335_;
 wire _10336_;
 wire _10337_;
 wire _10338_;
 wire _10339_;
 wire _10340_;
 wire _10341_;
 wire _10342_;
 wire _10343_;
 wire _10344_;
 wire _10345_;
 wire _10346_;
 wire _10347_;
 wire _10348_;
 wire _10349_;
 wire _10350_;
 wire _10351_;
 wire _10352_;
 wire _10353_;
 wire _10354_;
 wire _10355_;
 wire _10356_;
 wire _10357_;
 wire _10358_;
 wire _10359_;
 wire _10360_;
 wire _10361_;
 wire _10362_;
 wire _10363_;
 wire _10364_;
 wire _10365_;
 wire _10366_;
 wire _10367_;
 wire _10368_;
 wire _10369_;
 wire _10370_;
 wire _10371_;
 wire _10372_;
 wire _10373_;
 wire _10374_;
 wire _10375_;
 wire _10376_;
 wire _10377_;
 wire _10378_;
 wire _10379_;
 wire _10380_;
 wire _10381_;
 wire _10382_;
 wire _10383_;
 wire _10384_;
 wire _10385_;
 wire _10386_;
 wire _10387_;
 wire _10388_;
 wire _10389_;
 wire _10390_;
 wire _10391_;
 wire _10392_;
 wire _10393_;
 wire _10394_;
 wire _10395_;
 wire _10396_;
 wire _10397_;
 wire _10398_;
 wire _10399_;
 wire _10400_;
 wire _10401_;
 wire _10402_;
 wire _10403_;
 wire _10404_;
 wire _10405_;
 wire _10406_;
 wire _10407_;
 wire _10408_;
 wire _10409_;
 wire _10410_;
 wire _10411_;
 wire _10412_;
 wire _10413_;
 wire _10414_;
 wire _10415_;
 wire _10416_;
 wire _10417_;
 wire _10418_;
 wire _10419_;
 wire _10420_;
 wire _10421_;
 wire _10422_;
 wire _10423_;
 wire _10424_;
 wire _10425_;
 wire _10426_;
 wire _10427_;
 wire _10428_;
 wire _10429_;
 wire _10430_;
 wire _10431_;
 wire _10432_;
 wire _10433_;
 wire _10434_;
 wire _10435_;
 wire _10436_;
 wire _10437_;
 wire _10438_;
 wire _10439_;
 wire _10440_;
 wire _10441_;
 wire _10442_;
 wire _10443_;
 wire _10444_;
 wire _10445_;
 wire _10446_;
 wire _10447_;
 wire _10448_;
 wire _10449_;
 wire _10450_;
 wire _10451_;
 wire _10452_;
 wire _10453_;
 wire _10454_;
 wire _10455_;
 wire _10456_;
 wire _10457_;
 wire _10458_;
 wire _10459_;
 wire _10460_;
 wire _10461_;
 wire _10462_;
 wire _10463_;
 wire _10464_;
 wire _10465_;
 wire _10466_;
 wire _10467_;
 wire _10468_;
 wire _10469_;
 wire _10470_;
 wire _10471_;
 wire _10472_;
 wire _10473_;
 wire _10474_;
 wire _10475_;
 wire _10476_;
 wire _10477_;
 wire _10478_;
 wire _10479_;
 wire _10480_;
 wire _10481_;
 wire _10482_;
 wire _10483_;
 wire _10484_;
 wire _10485_;
 wire _10486_;
 wire _10487_;
 wire _10488_;
 wire _10489_;
 wire _10490_;
 wire _10491_;
 wire _10492_;
 wire _10493_;
 wire _10494_;
 wire _10495_;
 wire _10496_;
 wire _10497_;
 wire _10498_;
 wire _10499_;
 wire _10500_;
 wire _10501_;
 wire _10502_;
 wire _10503_;
 wire _10504_;
 wire _10505_;
 wire _10506_;
 wire _10507_;
 wire _10508_;
 wire _10509_;
 wire _10510_;
 wire _10511_;
 wire _10512_;
 wire _10513_;
 wire _10514_;
 wire _10515_;
 wire _10516_;
 wire _10517_;
 wire _10518_;
 wire _10519_;
 wire _10520_;
 wire _10521_;
 wire _10522_;
 wire _10523_;
 wire _10524_;
 wire _10525_;
 wire _10526_;
 wire _10527_;
 wire _10528_;
 wire _10529_;
 wire _10530_;
 wire _10531_;
 wire _10532_;
 wire _10533_;
 wire _10534_;
 wire _10535_;
 wire _10536_;
 wire _10537_;
 wire _10538_;
 wire _10539_;
 wire _10540_;
 wire _10541_;
 wire _10542_;
 wire _10543_;
 wire _10544_;
 wire _10545_;
 wire _10546_;
 wire _10547_;
 wire _10548_;
 wire _10549_;
 wire _10550_;
 wire _10551_;
 wire _10552_;
 wire _10553_;
 wire _10554_;
 wire _10555_;
 wire _10556_;
 wire _10557_;
 wire _10558_;
 wire _10559_;
 wire _10560_;
 wire _10561_;
 wire _10562_;
 wire _10563_;
 wire _10564_;
 wire _10565_;
 wire _10566_;
 wire _10567_;
 wire _10568_;
 wire _10569_;
 wire _10570_;
 wire _10571_;
 wire _10572_;
 wire _10573_;
 wire _10574_;
 wire _10575_;
 wire _10576_;
 wire _10577_;
 wire _10578_;
 wire _10579_;
 wire _10580_;
 wire _10581_;
 wire _10582_;
 wire _10583_;
 wire _10584_;
 wire _10585_;
 wire _10586_;
 wire _10587_;
 wire _10588_;
 wire _10589_;
 wire _10590_;
 wire _10591_;
 wire _10592_;
 wire _10593_;
 wire _10594_;
 wire _10595_;
 wire _10596_;
 wire _10597_;
 wire _10598_;
 wire _10599_;
 wire _10600_;
 wire _10601_;
 wire _10602_;
 wire _10603_;
 wire _10604_;
 wire _10605_;
 wire _10606_;
 wire _10607_;
 wire _10608_;
 wire _10609_;
 wire _10610_;
 wire _10611_;
 wire _10612_;
 wire _10613_;
 wire _10614_;
 wire _10615_;
 wire _10616_;
 wire _10617_;
 wire _10618_;
 wire _10619_;
 wire _10620_;
 wire _10621_;
 wire _10622_;
 wire _10623_;
 wire _10624_;
 wire _10625_;
 wire _10626_;
 wire _10627_;
 wire _10628_;
 wire _10629_;
 wire _10630_;
 wire _10631_;
 wire _10632_;
 wire _10633_;
 wire _10634_;
 wire _10635_;
 wire _10636_;
 wire _10637_;
 wire _10638_;
 wire _10639_;
 wire _10640_;
 wire _10641_;
 wire _10642_;
 wire _10643_;
 wire _10644_;
 wire _10645_;
 wire _10646_;
 wire _10647_;
 wire _10648_;
 wire _10649_;
 wire _10650_;
 wire _10651_;
 wire _10652_;
 wire _10653_;
 wire _10654_;
 wire _10655_;
 wire _10656_;
 wire _10657_;
 wire _10658_;
 wire _10659_;
 wire _10660_;
 wire _10661_;
 wire _10662_;
 wire _10663_;
 wire _10664_;
 wire _10665_;
 wire _10666_;
 wire _10667_;
 wire _10668_;
 wire _10669_;
 wire _10670_;
 wire _10671_;
 wire _10672_;
 wire _10673_;
 wire _10674_;
 wire _10675_;
 wire _10676_;
 wire _10677_;
 wire _10678_;
 wire _10679_;
 wire _10680_;
 wire _10681_;
 wire _10682_;
 wire _10683_;
 wire _10684_;
 wire _10685_;
 wire _10686_;
 wire _10687_;
 wire _10688_;
 wire _10689_;
 wire _10690_;
 wire _10691_;
 wire _10692_;
 wire _10693_;
 wire _10694_;
 wire _10695_;
 wire _10696_;
 wire _10697_;
 wire _10698_;
 wire _10699_;
 wire _10700_;
 wire _10701_;
 wire _10702_;
 wire _10703_;
 wire _10704_;
 wire _10705_;
 wire _10706_;
 wire _10707_;
 wire _10708_;
 wire _10709_;
 wire _10710_;
 wire _10711_;
 wire _10712_;
 wire _10713_;
 wire _10714_;
 wire _10715_;
 wire _10716_;
 wire _10717_;
 wire _10718_;
 wire _10719_;
 wire _10720_;
 wire _10721_;
 wire _10722_;
 wire _10723_;
 wire _10724_;
 wire _10725_;
 wire _10726_;
 wire _10727_;
 wire _10728_;
 wire _10729_;
 wire _10730_;
 wire _10731_;
 wire _10732_;
 wire _10733_;
 wire _10734_;
 wire _10735_;
 wire _10736_;
 wire _10737_;
 wire _10738_;
 wire _10739_;
 wire _10740_;
 wire _10741_;
 wire _10742_;
 wire _10743_;
 wire _10744_;
 wire _10745_;
 wire _10746_;
 wire _10747_;
 wire _10748_;
 wire _10749_;
 wire _10750_;
 wire _10751_;
 wire _10752_;
 wire _10753_;
 wire _10754_;
 wire _10755_;
 wire _10756_;
 wire _10757_;
 wire _10758_;
 wire _10759_;
 wire _10760_;
 wire _10761_;
 wire _10762_;
 wire _10763_;
 wire _10764_;
 wire _10765_;
 wire _10766_;
 wire _10767_;
 wire _10768_;
 wire _10769_;
 wire _10770_;
 wire _10771_;
 wire _10772_;
 wire _10773_;
 wire _10774_;
 wire _10775_;
 wire _10776_;
 wire _10777_;
 wire _10778_;
 wire _10779_;
 wire _10780_;
 wire _10781_;
 wire _10782_;
 wire _10783_;
 wire _10784_;
 wire _10785_;
 wire _10786_;
 wire _10787_;
 wire _10788_;
 wire _10789_;
 wire _10790_;
 wire _10791_;
 wire _10792_;
 wire _10793_;
 wire _10794_;
 wire _10795_;
 wire _10796_;
 wire _10797_;
 wire _10798_;
 wire _10799_;
 wire _10800_;
 wire _10801_;
 wire _10802_;
 wire _10803_;
 wire _10804_;
 wire _10805_;
 wire _10806_;
 wire _10807_;
 wire _10808_;
 wire _10809_;
 wire _10810_;
 wire _10811_;
 wire _10812_;
 wire _10813_;
 wire _10814_;
 wire _10815_;
 wire _10816_;
 wire _10817_;
 wire _10818_;
 wire _10819_;
 wire _10820_;
 wire _10821_;
 wire _10822_;
 wire _10823_;
 wire _10824_;
 wire _10825_;
 wire _10826_;
 wire _10827_;
 wire _10828_;
 wire _10829_;
 wire _10830_;
 wire _10831_;
 wire _10832_;
 wire _10833_;
 wire _10834_;
 wire _10835_;
 wire _10836_;
 wire _10837_;
 wire _10838_;
 wire _10839_;
 wire _10840_;
 wire _10841_;
 wire _10842_;
 wire _10843_;
 wire _10844_;
 wire _10845_;
 wire _10846_;
 wire _10847_;
 wire _10848_;
 wire _10849_;
 wire _10850_;
 wire _10851_;
 wire _10852_;
 wire _10853_;
 wire _10854_;
 wire _10855_;
 wire _10856_;
 wire _10857_;
 wire _10858_;
 wire _10859_;
 wire _10860_;
 wire _10861_;
 wire _10862_;
 wire _10863_;
 wire _10864_;
 wire _10865_;
 wire _10866_;
 wire _10867_;
 wire _10868_;
 wire _10869_;
 wire _10870_;
 wire _10871_;
 wire _10872_;
 wire _10873_;
 wire _10874_;
 wire _10875_;
 wire _10876_;
 wire _10877_;
 wire _10878_;
 wire _10879_;
 wire _10880_;
 wire _10881_;
 wire _10882_;
 wire _10883_;
 wire _10884_;
 wire _10885_;
 wire _10886_;
 wire _10887_;
 wire _10888_;
 wire _10889_;
 wire _10890_;
 wire _10891_;
 wire _10892_;
 wire _10893_;
 wire _10894_;
 wire _10895_;
 wire _10896_;
 wire _10897_;
 wire _10898_;
 wire _10899_;
 wire _10900_;
 wire _10901_;
 wire _10902_;
 wire _10903_;
 wire _10904_;
 wire _10905_;
 wire _10906_;
 wire _10907_;
 wire _10908_;
 wire _10909_;
 wire _10910_;
 wire _10911_;
 wire _10912_;
 wire _10913_;
 wire _10914_;
 wire _10915_;
 wire _10916_;
 wire _10917_;
 wire _10918_;
 wire _10919_;
 wire _10920_;
 wire _10921_;
 wire _10922_;
 wire _10923_;
 wire _10924_;
 wire _10925_;
 wire _10926_;
 wire _10927_;
 wire _10928_;
 wire _10929_;
 wire _10930_;
 wire _10931_;
 wire _10932_;
 wire _10933_;
 wire _10934_;
 wire _10935_;
 wire _10936_;
 wire _10937_;
 wire _10938_;
 wire _10939_;
 wire _10940_;
 wire _10941_;
 wire _10942_;
 wire _10943_;
 wire _10944_;
 wire _10945_;
 wire _10946_;
 wire _10947_;
 wire _10948_;
 wire _10949_;
 wire _10950_;
 wire _10951_;
 wire _10952_;
 wire _10953_;
 wire _10954_;
 wire _10955_;
 wire _10956_;
 wire _10957_;
 wire _10958_;
 wire _10959_;
 wire _10960_;
 wire _10961_;
 wire _10962_;
 wire _10963_;
 wire _10964_;
 wire _10965_;
 wire _10966_;
 wire _10967_;
 wire _10968_;
 wire _10969_;
 wire _10970_;
 wire _10971_;
 wire _10972_;
 wire _10973_;
 wire _10974_;
 wire _10975_;
 wire _10976_;
 wire _10977_;
 wire _10978_;
 wire _10979_;
 wire _10980_;
 wire _10981_;
 wire _10982_;
 wire _10983_;
 wire _10984_;
 wire _10985_;
 wire _10986_;
 wire _10987_;
 wire _10988_;
 wire _10989_;
 wire _10990_;
 wire _10991_;
 wire _10992_;
 wire _10993_;
 wire _10994_;
 wire _10995_;
 wire _10996_;
 wire _10997_;
 wire _10998_;
 wire _10999_;
 wire _11000_;
 wire _11001_;
 wire _11002_;
 wire _11003_;
 wire _11004_;
 wire _11005_;
 wire _11006_;
 wire _11007_;
 wire _11008_;
 wire _11009_;
 wire _11010_;
 wire _11011_;
 wire _11012_;
 wire _11013_;
 wire _11014_;
 wire _11015_;
 wire _11016_;
 wire _11017_;
 wire _11018_;
 wire _11019_;
 wire _11020_;
 wire _11021_;
 wire _11022_;
 wire _11023_;
 wire _11024_;
 wire _11025_;
 wire _11026_;
 wire _11027_;
 wire _11028_;
 wire _11029_;
 wire _11030_;
 wire _11031_;
 wire _11032_;
 wire _11033_;
 wire _11034_;
 wire _11035_;
 wire _11036_;
 wire _11037_;
 wire _11038_;
 wire _11039_;
 wire _11040_;
 wire _11041_;
 wire _11042_;
 wire _11043_;
 wire _11044_;
 wire _11045_;
 wire _11046_;
 wire _11047_;
 wire _11048_;
 wire _11049_;
 wire _11050_;
 wire _11051_;
 wire _11052_;
 wire _11053_;
 wire _11054_;
 wire _11055_;
 wire _11056_;
 wire _11057_;
 wire _11058_;
 wire _11059_;
 wire _11060_;
 wire _11061_;
 wire _11062_;
 wire _11063_;
 wire _11064_;
 wire _11065_;
 wire _11066_;
 wire _11067_;
 wire _11068_;
 wire _11069_;
 wire _11070_;
 wire _11071_;
 wire _11072_;
 wire _11073_;
 wire _11074_;
 wire _11075_;
 wire _11076_;
 wire _11077_;
 wire _11078_;
 wire _11079_;
 wire _11080_;
 wire _11081_;
 wire _11082_;
 wire _11083_;
 wire _11084_;
 wire _11085_;
 wire _11086_;
 wire _11087_;
 wire _11088_;
 wire _11089_;
 wire _11090_;
 wire _11091_;
 wire _11092_;
 wire _11093_;
 wire _11094_;
 wire _11095_;
 wire _11096_;
 wire _11097_;
 wire _11098_;
 wire _11099_;
 wire _11100_;
 wire _11101_;
 wire _11102_;
 wire _11103_;
 wire _11104_;
 wire _11105_;
 wire _11106_;
 wire _11107_;
 wire _11108_;
 wire _11109_;
 wire _11110_;
 wire _11111_;
 wire _11112_;
 wire _11113_;
 wire _11114_;
 wire _11115_;
 wire _11116_;
 wire _11117_;
 wire _11118_;
 wire _11119_;
 wire _11120_;
 wire _11121_;
 wire _11122_;
 wire _11123_;
 wire _11124_;
 wire _11125_;
 wire _11126_;
 wire _11127_;
 wire _11128_;
 wire _11129_;
 wire _11130_;
 wire _11131_;
 wire _11132_;
 wire _11133_;
 wire _11134_;
 wire _11135_;
 wire _11136_;
 wire _11137_;
 wire _11138_;
 wire _11139_;
 wire _11140_;
 wire _11141_;
 wire _11142_;
 wire _11143_;
 wire _11144_;
 wire _11145_;
 wire _11146_;
 wire _11147_;
 wire _11148_;
 wire _11149_;
 wire _11150_;
 wire _11151_;
 wire _11152_;
 wire _11153_;
 wire _11154_;
 wire _11155_;
 wire _11156_;
 wire _11157_;
 wire _11158_;
 wire _11159_;
 wire _11160_;
 wire _11161_;
 wire _11162_;
 wire _11163_;
 wire _11164_;
 wire _11165_;
 wire _11166_;
 wire _11167_;
 wire _11168_;
 wire _11169_;
 wire _11170_;
 wire _11171_;
 wire _11172_;
 wire _11173_;
 wire _11174_;
 wire _11175_;
 wire _11176_;
 wire _11177_;
 wire _11178_;
 wire _11179_;
 wire _11180_;
 wire _11181_;
 wire _11182_;
 wire _11183_;
 wire _11184_;
 wire _11185_;
 wire _11186_;
 wire _11187_;
 wire _11188_;
 wire _11189_;
 wire _11190_;
 wire _11191_;
 wire _11192_;
 wire _11193_;
 wire _11194_;
 wire _11195_;
 wire _11196_;
 wire _11197_;
 wire _11198_;
 wire _11199_;
 wire _11200_;
 wire _11201_;
 wire _11202_;
 wire _11203_;
 wire _11204_;
 wire _11205_;
 wire _11206_;
 wire _11207_;
 wire _11208_;
 wire _11209_;
 wire _11210_;
 wire _11211_;
 wire _11212_;
 wire _11213_;
 wire _11214_;
 wire _11215_;
 wire _11216_;
 wire _11217_;
 wire _11218_;
 wire _11219_;
 wire _11220_;
 wire _11221_;
 wire _11222_;
 wire _11223_;
 wire _11224_;
 wire _11225_;
 wire _11226_;
 wire _11227_;
 wire _11228_;
 wire _11229_;
 wire _11230_;
 wire _11231_;
 wire _11232_;
 wire _11233_;
 wire _11234_;
 wire _11235_;
 wire _11236_;
 wire _11237_;
 wire _11238_;
 wire _11239_;
 wire _11240_;
 wire _11241_;
 wire _11242_;
 wire _11243_;
 wire _11244_;
 wire _11245_;
 wire _11246_;
 wire _11247_;
 wire _11248_;
 wire _11249_;
 wire _11250_;
 wire _11251_;
 wire _11252_;
 wire _11253_;
 wire _11254_;
 wire _11255_;
 wire _11256_;
 wire _11257_;
 wire _11258_;
 wire _11259_;
 wire _11260_;
 wire _11261_;
 wire _11262_;
 wire _11263_;
 wire _11264_;
 wire _11265_;
 wire _11266_;
 wire _11267_;
 wire _11268_;
 wire _11269_;
 wire _11270_;
 wire _11271_;
 wire _11272_;
 wire _11273_;
 wire _11274_;
 wire _11275_;
 wire _11276_;
 wire _11277_;
 wire _11278_;
 wire _11279_;
 wire _11280_;
 wire _11281_;
 wire _11282_;
 wire _11283_;
 wire _11284_;
 wire _11285_;
 wire _11286_;
 wire _11287_;
 wire _11288_;
 wire _11289_;
 wire _11290_;
 wire _11291_;
 wire _11292_;
 wire _11293_;
 wire _11294_;
 wire _11295_;
 wire _11296_;
 wire _11297_;
 wire _11298_;
 wire _11299_;
 wire _11300_;
 wire _11301_;
 wire _11302_;
 wire _11303_;
 wire _11304_;
 wire _11305_;
 wire _11306_;
 wire _11307_;
 wire _11308_;
 wire _11309_;
 wire _11310_;
 wire _11311_;
 wire _11312_;
 wire _11313_;
 wire _11314_;
 wire _11315_;
 wire _11316_;
 wire _11317_;
 wire _11318_;
 wire _11319_;
 wire _11320_;
 wire _11321_;
 wire _11322_;
 wire _11323_;
 wire _11324_;
 wire _11325_;
 wire _11326_;
 wire _11327_;
 wire _11328_;
 wire _11329_;
 wire _11330_;
 wire _11331_;
 wire _11332_;
 wire _11333_;
 wire _11334_;
 wire _11335_;
 wire _11336_;
 wire _11337_;
 wire _11338_;
 wire _11339_;
 wire _11340_;
 wire _11341_;
 wire _11342_;
 wire _11343_;
 wire _11344_;
 wire _11345_;
 wire _11346_;
 wire _11347_;
 wire _11348_;
 wire _11349_;
 wire _11350_;
 wire _11351_;
 wire _11352_;
 wire _11353_;
 wire _11354_;
 wire _11355_;
 wire _11356_;
 wire _11357_;
 wire _11358_;
 wire _11359_;
 wire _11360_;
 wire _11361_;
 wire _11362_;
 wire _11363_;
 wire _11364_;
 wire _11365_;
 wire _11366_;
 wire _11367_;
 wire _11368_;
 wire _11369_;
 wire _11370_;
 wire _11371_;
 wire _11372_;
 wire _11373_;
 wire _11374_;
 wire _11375_;
 wire _11376_;
 wire _11377_;
 wire _11378_;
 wire _11379_;
 wire _11380_;
 wire _11381_;
 wire _11382_;
 wire _11383_;
 wire _11384_;
 wire _11385_;
 wire _11386_;
 wire _11387_;
 wire _11388_;
 wire _11389_;
 wire _11390_;
 wire _11391_;
 wire _11392_;
 wire _11393_;
 wire _11394_;
 wire _11395_;
 wire _11396_;
 wire _11397_;
 wire _11398_;
 wire _11399_;
 wire _11400_;
 wire _11401_;
 wire _11402_;
 wire _11403_;
 wire _11404_;
 wire _11405_;
 wire _11406_;
 wire _11407_;
 wire _11408_;
 wire _11409_;
 wire _11410_;
 wire _11411_;
 wire _11412_;
 wire _11413_;
 wire _11414_;
 wire _11415_;
 wire _11416_;
 wire _11417_;
 wire _11418_;
 wire _11419_;
 wire _11420_;
 wire _11421_;
 wire _11422_;
 wire _11423_;
 wire _11424_;
 wire _11425_;
 wire _11426_;
 wire _11427_;
 wire _11428_;
 wire _11429_;
 wire _11430_;
 wire _11431_;
 wire _11432_;
 wire _11433_;
 wire _11434_;
 wire _11435_;
 wire _11436_;
 wire _11437_;
 wire _11438_;
 wire _11439_;
 wire _11440_;
 wire _11441_;
 wire _11442_;
 wire _11443_;
 wire _11444_;
 wire _11445_;
 wire _11446_;
 wire _11447_;
 wire _11448_;
 wire _11449_;
 wire _11450_;
 wire _11451_;
 wire _11452_;
 wire _11453_;
 wire _11454_;
 wire _11455_;
 wire _11456_;
 wire _11457_;
 wire _11458_;
 wire _11459_;
 wire _11460_;
 wire _11461_;
 wire _11462_;
 wire _11463_;
 wire _11464_;
 wire _11465_;
 wire _11466_;
 wire _11467_;
 wire _11468_;
 wire _11469_;
 wire _11470_;
 wire _11471_;
 wire _11472_;
 wire _11473_;
 wire _11474_;
 wire _11475_;
 wire _11476_;
 wire _11477_;
 wire _11478_;
 wire _11479_;
 wire _11480_;
 wire _11481_;
 wire _11482_;
 wire _11483_;
 wire _11484_;
 wire _11485_;
 wire _11486_;
 wire _11487_;
 wire _11488_;
 wire _11489_;
 wire _11490_;
 wire _11491_;
 wire _11492_;
 wire _11493_;
 wire _11494_;
 wire _11495_;
 wire _11496_;
 wire _11497_;
 wire _11498_;
 wire _11499_;
 wire _11500_;
 wire _11501_;
 wire _11502_;
 wire _11503_;
 wire _11504_;
 wire _11505_;
 wire _11506_;
 wire _11507_;
 wire _11508_;
 wire _11509_;
 wire _11510_;
 wire _11511_;
 wire _11512_;
 wire _11513_;
 wire _11514_;
 wire _11515_;
 wire _11516_;
 wire _11517_;
 wire _11518_;
 wire _11519_;
 wire _11520_;
 wire _11521_;
 wire _11522_;
 wire _11523_;
 wire _11524_;
 wire _11525_;
 wire _11526_;
 wire _11527_;
 wire _11528_;
 wire _11529_;
 wire _11530_;
 wire _11531_;
 wire _11532_;
 wire _11533_;
 wire _11534_;
 wire _11535_;
 wire _11536_;
 wire _11537_;
 wire _11538_;
 wire _11539_;
 wire _11540_;
 wire _11541_;
 wire _11542_;
 wire _11543_;
 wire _11544_;
 wire _11545_;
 wire _11546_;
 wire _11547_;
 wire _11548_;
 wire _11549_;
 wire _11550_;
 wire _11551_;
 wire _11552_;
 wire _11553_;
 wire _11554_;
 wire _11555_;
 wire _11556_;
 wire _11557_;
 wire _11558_;
 wire _11559_;
 wire _11560_;
 wire _11561_;
 wire _11562_;
 wire _11563_;
 wire _11564_;
 wire _11565_;
 wire _11566_;
 wire _11567_;
 wire _11568_;
 wire _11569_;
 wire _11570_;
 wire _11571_;
 wire _11572_;
 wire _11573_;
 wire _11574_;
 wire _11575_;
 wire _11576_;
 wire _11577_;
 wire _11578_;
 wire _11579_;
 wire _11580_;
 wire _11581_;
 wire _11582_;
 wire _11583_;
 wire _11584_;
 wire _11585_;
 wire _11586_;
 wire _11587_;
 wire _11588_;
 wire _11589_;
 wire _11590_;
 wire _11591_;
 wire _11592_;
 wire _11593_;
 wire _11594_;
 wire _11595_;
 wire _11596_;
 wire _11597_;
 wire _11598_;
 wire _11599_;
 wire _11600_;
 wire _11601_;
 wire _11602_;
 wire _11603_;
 wire _11604_;
 wire _11605_;
 wire _11606_;
 wire _11607_;
 wire _11608_;
 wire _11609_;
 wire _11610_;
 wire _11611_;
 wire _11612_;
 wire _11613_;
 wire _11614_;
 wire _11615_;
 wire _11616_;
 wire _11617_;
 wire _11618_;
 wire _11619_;
 wire _11620_;
 wire _11621_;
 wire _11622_;
 wire _11623_;
 wire _11624_;
 wire _11625_;
 wire _11626_;
 wire _11627_;
 wire _11628_;
 wire _11629_;
 wire _11630_;
 wire _11631_;
 wire _11632_;
 wire _11633_;
 wire _11634_;
 wire _11635_;
 wire _11636_;
 wire _11637_;
 wire _11638_;
 wire _11639_;
 wire _11640_;
 wire _11641_;
 wire _11642_;
 wire _11643_;
 wire _11644_;
 wire _11645_;
 wire _11646_;
 wire _11647_;
 wire _11648_;
 wire _11649_;
 wire _11650_;
 wire _11651_;
 wire _11652_;
 wire _11653_;
 wire _11654_;
 wire _11655_;
 wire _11656_;
 wire _11657_;
 wire _11658_;
 wire _11659_;
 wire _11660_;
 wire _11661_;
 wire _11662_;
 wire _11663_;
 wire _11664_;
 wire _11665_;
 wire _11666_;
 wire _11667_;
 wire _11668_;
 wire _11669_;
 wire _11670_;
 wire _11671_;
 wire _11672_;
 wire _11673_;
 wire _11674_;
 wire _11675_;
 wire _11676_;
 wire _11677_;
 wire _11678_;
 wire _11679_;
 wire _11680_;
 wire _11681_;
 wire _11682_;
 wire _11683_;
 wire _11684_;
 wire _11685_;
 wire _11686_;
 wire _11687_;
 wire _11688_;
 wire _11689_;
 wire _11690_;
 wire _11691_;
 wire _11692_;
 wire _11693_;
 wire _11694_;
 wire _11695_;
 wire _11696_;
 wire _11697_;
 wire _11698_;
 wire _11699_;
 wire _11700_;
 wire _11701_;
 wire _11702_;
 wire _11703_;
 wire _11704_;
 wire _11705_;
 wire _11706_;
 wire _11707_;
 wire _11708_;
 wire _11709_;
 wire _11710_;
 wire _11711_;
 wire _11712_;
 wire _11713_;
 wire _11714_;
 wire _11715_;
 wire _11716_;
 wire _11717_;
 wire _11718_;
 wire _11719_;
 wire _11720_;
 wire _11721_;
 wire _11722_;
 wire _11723_;
 wire _11724_;
 wire _11725_;
 wire _11726_;
 wire _11727_;
 wire _11728_;
 wire _11729_;
 wire _11730_;
 wire _11731_;
 wire _11732_;
 wire _11733_;
 wire _11734_;
 wire _11735_;
 wire _11736_;
 wire _11737_;
 wire _11738_;
 wire _11739_;
 wire _11740_;
 wire _11741_;
 wire _11742_;
 wire _11743_;
 wire _11744_;
 wire _11745_;
 wire _11746_;
 wire _11747_;
 wire _11748_;
 wire _11749_;
 wire _11750_;
 wire _11751_;
 wire _11752_;
 wire _11753_;
 wire _11754_;
 wire _11755_;
 wire _11756_;
 wire _11757_;
 wire _11758_;
 wire _11759_;
 wire _11760_;
 wire _11761_;
 wire _11762_;
 wire _11763_;
 wire _11764_;
 wire _11765_;
 wire _11766_;
 wire _11767_;
 wire _11768_;
 wire _11769_;
 wire _11770_;
 wire _11771_;
 wire _11772_;
 wire _11773_;
 wire _11774_;
 wire _11775_;
 wire _11776_;
 wire _11777_;
 wire _11778_;
 wire _11779_;
 wire _11780_;
 wire _11781_;
 wire _11782_;
 wire _11783_;
 wire _11784_;
 wire _11785_;
 wire _11786_;
 wire _11787_;
 wire _11788_;
 wire _11789_;
 wire _11790_;
 wire _11791_;
 wire _11792_;
 wire _11793_;
 wire _11794_;
 wire _11795_;
 wire _11796_;
 wire _11797_;
 wire _11798_;
 wire _11799_;
 wire _11800_;
 wire _11801_;
 wire _11802_;
 wire _11803_;
 wire _11804_;
 wire _11805_;
 wire _11806_;
 wire _11807_;
 wire _11808_;
 wire _11809_;
 wire _11810_;
 wire _11811_;
 wire _11812_;
 wire _11813_;
 wire _11814_;
 wire _11815_;
 wire _11816_;
 wire _11817_;
 wire _11818_;
 wire _11819_;
 wire _11820_;
 wire _11821_;
 wire _11822_;
 wire _11823_;
 wire _11824_;
 wire _11825_;
 wire _11826_;
 wire _11827_;
 wire _11828_;
 wire _11829_;
 wire _11830_;
 wire _11831_;
 wire _11832_;
 wire _11833_;
 wire _11834_;
 wire _11835_;
 wire _11836_;
 wire _11837_;
 wire _11838_;
 wire _11839_;
 wire _11840_;
 wire _11841_;
 wire _11842_;
 wire _11843_;
 wire _11844_;
 wire _11845_;
 wire _11846_;
 wire _11847_;
 wire _11848_;
 wire _11849_;
 wire _11850_;
 wire _11851_;
 wire _11852_;
 wire _11853_;
 wire _11854_;
 wire _11855_;
 wire _11856_;
 wire _11857_;
 wire _11858_;
 wire _11859_;
 wire _11860_;
 wire _11861_;
 wire _11862_;
 wire _11863_;
 wire _11864_;
 wire _11865_;
 wire _11866_;
 wire _11867_;
 wire _11868_;
 wire _11869_;
 wire _11870_;
 wire _11871_;
 wire _11872_;
 wire _11873_;
 wire _11874_;
 wire _11875_;
 wire _11876_;
 wire _11877_;
 wire _11878_;
 wire _11879_;
 wire _11880_;
 wire _11881_;
 wire _11882_;
 wire _11883_;
 wire _11884_;
 wire _11885_;
 wire _11886_;
 wire _11887_;
 wire _11888_;
 wire _11889_;
 wire _11890_;
 wire _11891_;
 wire _11892_;
 wire _11893_;
 wire _11894_;
 wire _11895_;
 wire _11896_;
 wire _11897_;
 wire _11898_;
 wire _11899_;
 wire _11900_;
 wire _11901_;
 wire _11902_;
 wire _11903_;
 wire _11904_;
 wire _11905_;
 wire _11906_;
 wire _11907_;
 wire _11908_;
 wire _11909_;
 wire _11910_;
 wire _11911_;
 wire _11912_;
 wire _11913_;
 wire _11914_;
 wire _11915_;
 wire _11916_;
 wire _11917_;
 wire _11918_;
 wire _11919_;
 wire _11920_;
 wire _11921_;
 wire _11922_;
 wire _11923_;
 wire _11924_;
 wire _11925_;
 wire _11926_;
 wire _11927_;
 wire _11928_;
 wire _11929_;
 wire _11930_;
 wire _11931_;
 wire _11932_;
 wire _11933_;
 wire _11934_;
 wire _11935_;
 wire _11936_;
 wire _11937_;
 wire _11938_;
 wire _11939_;
 wire _11940_;
 wire _11941_;
 wire _11942_;
 wire _11943_;
 wire _11944_;
 wire _11945_;
 wire _11946_;
 wire _11947_;
 wire _11948_;
 wire _11949_;
 wire _11950_;
 wire _11951_;
 wire _11952_;
 wire _11953_;
 wire _11954_;
 wire _11955_;
 wire _11956_;
 wire _11957_;
 wire _11958_;
 wire _11959_;
 wire _11960_;
 wire _11961_;
 wire _11962_;
 wire _11963_;
 wire _11964_;
 wire _11965_;
 wire _11966_;
 wire _11967_;
 wire _11968_;
 wire _11969_;
 wire _11970_;
 wire _11971_;
 wire _11972_;
 wire _11973_;
 wire _11974_;
 wire _11975_;
 wire _11976_;
 wire _11977_;
 wire _11978_;
 wire _11979_;
 wire _11980_;
 wire _11981_;
 wire _11982_;
 wire _11983_;
 wire _11984_;
 wire _11985_;
 wire _11986_;
 wire _11987_;
 wire _11988_;
 wire _11989_;
 wire _11990_;
 wire _11991_;
 wire _11992_;
 wire _11993_;
 wire _11994_;
 wire _11995_;
 wire _11996_;
 wire _11997_;
 wire _11998_;
 wire _11999_;
 wire _12000_;
 wire _12001_;
 wire _12002_;
 wire _12003_;
 wire _12004_;
 wire _12005_;
 wire _12006_;
 wire _12007_;
 wire _12008_;
 wire _12009_;
 wire _12010_;
 wire _12011_;
 wire _12012_;
 wire _12013_;
 wire _12014_;
 wire _12015_;
 wire _12016_;
 wire _12017_;
 wire _12018_;
 wire _12019_;
 wire _12020_;
 wire _12021_;
 wire _12022_;
 wire _12023_;
 wire _12024_;
 wire _12025_;
 wire _12026_;
 wire _12027_;
 wire _12028_;
 wire _12029_;
 wire _12030_;
 wire _12031_;
 wire _12032_;
 wire _12033_;
 wire _12034_;
 wire _12035_;
 wire _12036_;
 wire _12037_;
 wire _12038_;
 wire _12039_;
 wire _12040_;
 wire _12041_;
 wire _12042_;
 wire _12043_;
 wire _12044_;
 wire _12045_;
 wire _12046_;
 wire _12047_;
 wire _12048_;
 wire _12049_;
 wire _12050_;
 wire _12051_;
 wire _12052_;
 wire _12053_;
 wire _12054_;
 wire _12055_;
 wire _12056_;
 wire _12057_;
 wire _12058_;
 wire _12059_;
 wire _12060_;
 wire _12061_;
 wire _12062_;
 wire _12063_;
 wire _12064_;
 wire _12065_;
 wire _12066_;
 wire _12067_;
 wire _12068_;
 wire _12069_;
 wire _12070_;
 wire _12071_;
 wire _12072_;
 wire _12073_;
 wire _12074_;
 wire _12075_;
 wire _12076_;
 wire _12077_;
 wire _12078_;
 wire _12079_;
 wire _12080_;
 wire _12081_;
 wire _12082_;
 wire _12083_;
 wire _12084_;
 wire _12085_;
 wire _12086_;
 wire _12087_;
 wire _12088_;
 wire _12089_;
 wire _12090_;
 wire _12091_;
 wire _12092_;
 wire _12093_;
 wire _12094_;
 wire _12095_;
 wire _12096_;
 wire _12097_;
 wire _12098_;
 wire _12099_;
 wire _12100_;
 wire _12101_;
 wire _12102_;
 wire _12103_;
 wire _12104_;
 wire _12105_;
 wire _12106_;
 wire _12107_;
 wire _12108_;
 wire _12109_;
 wire _12110_;
 wire _12111_;
 wire _12112_;
 wire _12113_;
 wire _12114_;
 wire _12115_;
 wire _12116_;
 wire _12117_;
 wire _12118_;
 wire _12119_;
 wire _12120_;
 wire _12121_;
 wire _12122_;
 wire _12123_;
 wire _12124_;
 wire _12125_;
 wire _12126_;
 wire _12127_;
 wire _12128_;
 wire _12129_;
 wire _12130_;
 wire _12131_;
 wire _12132_;
 wire _12133_;
 wire _12134_;
 wire _12135_;
 wire _12136_;
 wire _12137_;
 wire _12138_;
 wire _12139_;
 wire _12140_;
 wire _12141_;
 wire _12142_;
 wire _12143_;
 wire _12144_;
 wire _12145_;
 wire _12146_;
 wire _12147_;
 wire _12148_;
 wire _12149_;
 wire _12150_;
 wire _12151_;
 wire _12152_;
 wire _12153_;
 wire _12154_;
 wire _12155_;
 wire _12156_;
 wire _12157_;
 wire _12158_;
 wire _12159_;
 wire _12160_;
 wire _12161_;
 wire _12162_;
 wire _12163_;
 wire _12164_;
 wire _12165_;
 wire _12166_;
 wire _12167_;
 wire _12168_;
 wire _12169_;
 wire _12170_;
 wire _12171_;
 wire _12172_;
 wire _12173_;
 wire _12174_;
 wire _12175_;
 wire _12176_;
 wire _12177_;
 wire _12178_;
 wire _12179_;
 wire _12180_;
 wire _12181_;
 wire _12182_;
 wire _12183_;
 wire _12184_;
 wire _12185_;
 wire _12186_;
 wire _12187_;
 wire _12188_;
 wire _12189_;
 wire _12190_;
 wire _12191_;
 wire _12192_;
 wire _12193_;
 wire _12194_;
 wire _12195_;
 wire _12196_;
 wire _12197_;
 wire _12198_;
 wire _12199_;
 wire _12200_;
 wire _12201_;
 wire _12202_;
 wire _12203_;
 wire _12204_;
 wire _12205_;
 wire _12206_;
 wire _12207_;
 wire _12208_;
 wire _12209_;
 wire _12210_;
 wire _12211_;
 wire _12212_;
 wire _12213_;
 wire _12214_;
 wire _12215_;
 wire _12216_;
 wire _12217_;
 wire _12218_;
 wire _12219_;
 wire _12220_;
 wire _12221_;
 wire _12222_;
 wire _12223_;
 wire _12224_;
 wire _12225_;
 wire _12226_;
 wire _12227_;
 wire _12228_;
 wire _12229_;
 wire _12230_;
 wire _12231_;
 wire _12232_;
 wire _12233_;
 wire _12234_;
 wire _12235_;
 wire _12236_;
 wire _12237_;
 wire _12238_;
 wire _12239_;
 wire _12240_;
 wire _12241_;
 wire _12242_;
 wire _12243_;
 wire _12244_;
 wire _12245_;
 wire _12246_;
 wire _12247_;
 wire _12248_;
 wire _12249_;
 wire _12250_;
 wire _12251_;
 wire _12252_;
 wire _12253_;
 wire _12254_;
 wire _12255_;
 wire _12256_;
 wire _12257_;
 wire _12258_;
 wire _12259_;
 wire _12260_;
 wire _12261_;
 wire _12262_;
 wire _12263_;
 wire _12264_;
 wire _12265_;
 wire _12266_;
 wire _12267_;
 wire _12268_;
 wire _12269_;
 wire _12270_;
 wire _12271_;
 wire _12272_;
 wire _12273_;
 wire _12274_;
 wire _12275_;
 wire _12276_;
 wire _12277_;
 wire _12278_;
 wire _12279_;
 wire _12280_;
 wire _12281_;
 wire _12282_;
 wire _12283_;
 wire _12284_;
 wire _12285_;
 wire _12286_;
 wire _12287_;
 wire _12288_;
 wire _12289_;
 wire _12290_;
 wire _12291_;
 wire _12292_;
 wire _12293_;
 wire _12294_;
 wire _12295_;
 wire _12296_;
 wire _12297_;
 wire _12298_;
 wire _12299_;
 wire _12300_;
 wire _12301_;
 wire _12302_;
 wire _12303_;
 wire _12304_;
 wire _12305_;
 wire _12306_;
 wire _12307_;
 wire _12308_;
 wire _12309_;
 wire _12310_;
 wire _12311_;
 wire _12312_;
 wire _12313_;
 wire _12314_;
 wire _12315_;
 wire _12316_;
 wire _12317_;
 wire _12318_;
 wire _12319_;
 wire _12320_;
 wire _12321_;
 wire _12322_;
 wire _12323_;
 wire _12324_;
 wire _12325_;
 wire _12326_;
 wire _12327_;
 wire _12328_;
 wire _12329_;
 wire _12330_;
 wire _12331_;
 wire _12332_;
 wire _12333_;
 wire _12334_;
 wire _12335_;
 wire _12336_;
 wire _12337_;
 wire _12338_;
 wire _12339_;
 wire _12340_;
 wire _12341_;
 wire _12342_;
 wire _12343_;
 wire _12344_;
 wire _12345_;
 wire _12346_;
 wire _12347_;
 wire _12348_;
 wire _12349_;
 wire _12350_;
 wire _12351_;
 wire _12352_;
 wire _12353_;
 wire _12354_;
 wire _12355_;
 wire _12356_;
 wire _12357_;
 wire _12358_;
 wire _12359_;
 wire _12360_;
 wire _12361_;
 wire _12362_;
 wire _12363_;
 wire _12364_;
 wire _12365_;
 wire _12366_;
 wire _12367_;
 wire _12368_;
 wire _12369_;
 wire _12370_;
 wire _12371_;
 wire _12372_;
 wire _12373_;
 wire _12374_;
 wire _12375_;
 wire _12376_;
 wire _12377_;
 wire _12378_;
 wire _12379_;
 wire _12380_;
 wire _12381_;
 wire _12382_;
 wire _12383_;
 wire _12384_;
 wire _12385_;
 wire _12386_;
 wire _12387_;
 wire _12388_;
 wire _12389_;
 wire _12390_;
 wire _12391_;
 wire _12392_;
 wire _12393_;
 wire _12394_;
 wire _12395_;
 wire _12396_;
 wire _12397_;
 wire _12398_;
 wire _12399_;
 wire _12400_;
 wire _12401_;
 wire _12402_;
 wire _12403_;
 wire _12404_;
 wire _12405_;
 wire _12406_;
 wire _12407_;
 wire _12408_;
 wire _12409_;
 wire _12410_;
 wire _12411_;
 wire _12412_;
 wire _12413_;
 wire _12414_;
 wire _12415_;
 wire _12416_;
 wire _12417_;
 wire _12418_;
 wire _12419_;
 wire _12420_;
 wire _12421_;
 wire _12422_;
 wire _12423_;
 wire _12424_;
 wire _12425_;
 wire _12426_;
 wire _12427_;
 wire _12428_;
 wire _12429_;
 wire _12430_;
 wire _12431_;
 wire _12432_;
 wire _12433_;
 wire _12434_;
 wire _12435_;
 wire _12436_;
 wire _12437_;
 wire _12438_;
 wire _12439_;
 wire _12440_;
 wire _12441_;
 wire _12442_;
 wire _12443_;
 wire _12444_;
 wire _12445_;
 wire _12446_;
 wire _12447_;
 wire _12448_;
 wire _12449_;
 wire _12450_;
 wire _12451_;
 wire _12452_;
 wire _12453_;
 wire _12454_;
 wire _12455_;
 wire _12456_;
 wire _12457_;
 wire _12458_;
 wire _12459_;
 wire _12460_;
 wire _12461_;
 wire _12462_;
 wire _12463_;
 wire _12464_;
 wire _12465_;
 wire _12466_;
 wire _12467_;
 wire _12468_;
 wire _12469_;
 wire _12470_;
 wire _12471_;
 wire _12472_;
 wire _12473_;
 wire _12474_;
 wire _12475_;
 wire _12476_;
 wire _12477_;
 wire _12478_;
 wire _12479_;
 wire _12480_;
 wire _12481_;
 wire _12482_;
 wire _12483_;
 wire _12484_;
 wire _12485_;
 wire _12486_;
 wire _12487_;
 wire _12488_;
 wire _12489_;
 wire _12490_;
 wire _12491_;
 wire _12492_;
 wire _12493_;
 wire _12494_;
 wire _12495_;
 wire _12496_;
 wire _12497_;
 wire _12498_;
 wire _12499_;
 wire _12500_;
 wire _12501_;
 wire _12502_;
 wire _12503_;
 wire _12504_;
 wire _12505_;
 wire _12506_;
 wire _12507_;
 wire _12508_;
 wire _12509_;
 wire _12510_;
 wire _12511_;
 wire _12512_;
 wire _12513_;
 wire _12514_;
 wire _12515_;
 wire _12516_;
 wire _12517_;
 wire _12518_;
 wire _12519_;
 wire _12520_;
 wire _12521_;
 wire _12522_;
 wire _12523_;
 wire _12524_;
 wire _12525_;
 wire _12526_;
 wire _12527_;
 wire _12528_;
 wire _12529_;
 wire _12530_;
 wire _12531_;
 wire _12532_;
 wire _12533_;
 wire _12534_;
 wire _12535_;
 wire _12536_;
 wire _12537_;
 wire _12538_;
 wire _12539_;
 wire _12540_;
 wire _12541_;
 wire _12542_;
 wire _12543_;
 wire _12544_;
 wire _12545_;
 wire _12546_;
 wire _12547_;
 wire _12548_;
 wire _12549_;
 wire _12550_;
 wire _12551_;
 wire _12552_;
 wire _12553_;
 wire _12554_;
 wire _12555_;
 wire _12556_;
 wire _12557_;
 wire _12558_;
 wire _12559_;
 wire _12560_;
 wire _12561_;
 wire _12562_;
 wire _12563_;
 wire _12564_;
 wire _12565_;
 wire _12566_;
 wire _12567_;
 wire _12568_;
 wire _12569_;
 wire _12570_;
 wire _12571_;
 wire _12572_;
 wire _12573_;
 wire _12574_;
 wire _12575_;
 wire _12576_;
 wire _12577_;
 wire _12578_;
 wire _12579_;
 wire _12580_;
 wire _12581_;
 wire _12582_;
 wire _12583_;
 wire _12584_;
 wire _12585_;
 wire _12586_;
 wire _12587_;
 wire _12588_;
 wire _12589_;
 wire _12590_;
 wire _12591_;
 wire _12592_;
 wire _12593_;
 wire _12594_;
 wire _12595_;
 wire _12596_;
 wire _12597_;
 wire _12598_;
 wire _12599_;
 wire _12600_;
 wire _12601_;
 wire _12602_;
 wire _12603_;
 wire _12604_;
 wire _12605_;
 wire _12606_;
 wire _12607_;
 wire _12608_;
 wire _12609_;
 wire _12610_;
 wire _12611_;
 wire _12612_;
 wire _12613_;
 wire _12614_;
 wire _12615_;
 wire _12616_;
 wire _12617_;
 wire _12618_;
 wire _12619_;
 wire _12620_;
 wire _12621_;
 wire _12622_;
 wire _12623_;
 wire _12624_;
 wire _12625_;
 wire _12626_;
 wire _12627_;
 wire _12628_;
 wire _12629_;
 wire _12630_;
 wire _12631_;
 wire _12632_;
 wire _12633_;
 wire _12634_;
 wire _12635_;
 wire _12636_;
 wire _12637_;
 wire _12638_;
 wire _12639_;
 wire _12640_;
 wire _12641_;
 wire _12642_;
 wire _12643_;
 wire _12644_;
 wire _12645_;
 wire _12646_;
 wire _12647_;
 wire _12648_;
 wire _12649_;
 wire _12650_;
 wire _12651_;
 wire _12652_;
 wire _12653_;
 wire _12654_;
 wire _12655_;
 wire _12656_;
 wire _12657_;
 wire _12658_;
 wire _12659_;
 wire _12660_;
 wire _12661_;
 wire _12662_;
 wire _12663_;
 wire _12664_;
 wire _12665_;
 wire _12666_;
 wire _12667_;
 wire _12668_;
 wire _12669_;
 wire _12670_;
 wire _12671_;
 wire _12672_;
 wire _12673_;
 wire _12674_;
 wire _12675_;
 wire _12676_;
 wire _12677_;
 wire _12678_;
 wire _12679_;
 wire _12680_;
 wire _12681_;
 wire _12682_;
 wire _12683_;
 wire _12684_;
 wire _12685_;
 wire _12686_;
 wire _12687_;
 wire _12688_;
 wire _12689_;
 wire _12690_;
 wire _12691_;
 wire _12692_;
 wire _12693_;
 wire _12694_;
 wire _12695_;
 wire _12696_;
 wire _12697_;
 wire _12698_;
 wire _12699_;
 wire _12700_;
 wire _12701_;
 wire _12702_;
 wire _12703_;
 wire _12704_;
 wire _12705_;
 wire _12706_;
 wire _12707_;
 wire _12708_;
 wire _12709_;
 wire _12710_;
 wire _12711_;
 wire _12712_;
 wire _12713_;
 wire _12714_;
 wire _12715_;
 wire _12716_;
 wire _12717_;
 wire _12718_;
 wire _12719_;
 wire _12720_;
 wire _12721_;
 wire _12722_;
 wire _12723_;
 wire _12724_;
 wire _12725_;
 wire _12726_;
 wire _12727_;
 wire _12728_;
 wire _12729_;
 wire _12730_;
 wire _12731_;
 wire _12732_;
 wire _12733_;
 wire _12734_;
 wire _12735_;
 wire _12736_;
 wire _12737_;
 wire _12738_;
 wire _12739_;
 wire _12740_;
 wire _12741_;
 wire _12742_;
 wire _12743_;
 wire _12744_;
 wire _12745_;
 wire _12746_;
 wire _12747_;
 wire _12748_;
 wire _12749_;
 wire _12750_;
 wire _12751_;
 wire _12752_;
 wire _12753_;
 wire _12754_;
 wire _12755_;
 wire _12756_;
 wire _12757_;
 wire _12758_;
 wire _12759_;
 wire _12760_;
 wire _12761_;
 wire _12762_;
 wire _12763_;
 wire _12764_;
 wire _12765_;
 wire _12766_;
 wire _12767_;
 wire _12768_;
 wire _12769_;
 wire _12770_;
 wire _12771_;
 wire _12772_;
 wire _12773_;
 wire _12774_;
 wire _12775_;
 wire _12776_;
 wire _12777_;
 wire _12778_;
 wire _12779_;
 wire _12780_;
 wire _12781_;
 wire _12782_;
 wire _12783_;
 wire _12784_;
 wire _12785_;
 wire _12786_;
 wire _12787_;
 wire _12788_;
 wire _12789_;
 wire _12790_;
 wire _12791_;
 wire _12792_;
 wire _12793_;
 wire _12794_;
 wire _12795_;
 wire _12796_;
 wire _12797_;
 wire _12798_;
 wire _12799_;
 wire _12800_;
 wire _12801_;
 wire _12802_;
 wire _12803_;
 wire _12804_;
 wire _12805_;
 wire _12806_;
 wire _12807_;
 wire _12808_;
 wire _12809_;
 wire _12810_;
 wire _12811_;
 wire _12812_;
 wire _12813_;
 wire _12814_;
 wire _12815_;
 wire _12816_;
 wire _12817_;
 wire _12818_;
 wire _12819_;
 wire _12820_;
 wire _12821_;
 wire _12822_;
 wire _12823_;
 wire _12824_;
 wire _12825_;
 wire _12826_;
 wire _12827_;
 wire _12828_;
 wire _12829_;
 wire _12830_;
 wire _12831_;
 wire _12832_;
 wire _12833_;
 wire _12834_;
 wire _12835_;
 wire _12836_;
 wire _12837_;
 wire _12838_;
 wire _12839_;
 wire _12840_;
 wire _12841_;
 wire _12842_;
 wire _12843_;
 wire _12844_;
 wire _12845_;
 wire _12846_;
 wire _12847_;
 wire _12848_;
 wire _12849_;
 wire _12850_;
 wire _12851_;
 wire _12852_;
 wire _12853_;
 wire _12854_;
 wire _12855_;
 wire _12856_;
 wire _12857_;
 wire _12858_;
 wire _12859_;
 wire _12860_;
 wire _12861_;
 wire _12862_;
 wire _12863_;
 wire _12864_;
 wire _12865_;
 wire _12866_;
 wire _12867_;
 wire _12868_;
 wire _12869_;
 wire _12870_;
 wire _12871_;
 wire _12872_;
 wire _12873_;
 wire _12874_;
 wire _12875_;
 wire _12876_;
 wire _12877_;
 wire _12878_;
 wire _12879_;
 wire _12880_;
 wire _12881_;
 wire _12882_;
 wire _12883_;
 wire _12884_;
 wire _12885_;
 wire _12886_;
 wire _12887_;
 wire _12888_;
 wire _12889_;
 wire _12890_;
 wire _12891_;
 wire _12892_;
 wire _12893_;
 wire _12894_;
 wire _12895_;
 wire _12896_;
 wire _12897_;
 wire _12898_;
 wire _12899_;
 wire _12900_;
 wire _12901_;
 wire _12902_;
 wire _12903_;
 wire _12904_;
 wire _12905_;
 wire _12906_;
 wire _12907_;
 wire _12908_;
 wire _12909_;
 wire _12910_;
 wire _12911_;
 wire _12912_;
 wire _12913_;
 wire _12914_;
 wire _12915_;
 wire _12916_;
 wire _12917_;
 wire _12918_;
 wire _12919_;
 wire _12920_;
 wire _12921_;
 wire _12922_;
 wire _12923_;
 wire _12924_;
 wire _12925_;
 wire _12926_;
 wire _12927_;
 wire _12928_;
 wire _12929_;
 wire _12930_;
 wire _12931_;
 wire _12932_;
 wire _12933_;
 wire _12934_;
 wire _12935_;
 wire _12936_;
 wire _12937_;
 wire _12938_;
 wire _12939_;
 wire _12940_;
 wire _12941_;
 wire _12942_;
 wire _12943_;
 wire _12944_;
 wire _12945_;
 wire _12946_;
 wire _12947_;
 wire _12948_;
 wire _12949_;
 wire _12950_;
 wire _12951_;
 wire _12952_;
 wire _12953_;
 wire _12954_;
 wire _12955_;
 wire _12956_;
 wire _12957_;
 wire _12958_;
 wire _12959_;
 wire _12960_;
 wire _12961_;
 wire _12962_;
 wire _12963_;
 wire _12964_;
 wire _12965_;
 wire _12966_;
 wire _12967_;
 wire _12968_;
 wire _12969_;
 wire _12970_;
 wire _12971_;
 wire _12972_;
 wire _12973_;
 wire _12974_;
 wire _12975_;
 wire _12976_;
 wire _12977_;
 wire _12978_;
 wire _12979_;
 wire _12980_;
 wire _12981_;
 wire _12982_;
 wire _12983_;
 wire _12984_;
 wire _12985_;
 wire _12986_;
 wire _12987_;
 wire _12988_;
 wire _12989_;
 wire _12990_;
 wire _12991_;
 wire _12992_;
 wire _12993_;
 wire _12994_;
 wire _12995_;
 wire _12996_;
 wire _12997_;
 wire _12998_;
 wire _12999_;
 wire _13000_;
 wire _13001_;
 wire _13002_;
 wire _13003_;
 wire _13004_;
 wire _13005_;
 wire _13006_;
 wire _13007_;
 wire _13008_;
 wire _13009_;
 wire _13010_;
 wire _13011_;
 wire _13012_;
 wire _13013_;
 wire _13014_;
 wire _13015_;
 wire _13016_;
 wire _13017_;
 wire _13018_;
 wire _13019_;
 wire _13020_;
 wire _13021_;
 wire _13022_;
 wire _13023_;
 wire _13024_;
 wire _13025_;
 wire _13026_;
 wire _13027_;
 wire _13028_;
 wire _13029_;
 wire _13030_;
 wire _13031_;
 wire _13032_;
 wire _13033_;
 wire _13034_;
 wire _13035_;
 wire _13036_;
 wire _13037_;
 wire _13038_;
 wire _13039_;
 wire _13040_;
 wire _13041_;
 wire _13042_;
 wire _13043_;
 wire _13044_;
 wire _13045_;
 wire _13046_;
 wire _13047_;
 wire _13048_;
 wire _13049_;
 wire _13050_;
 wire _13051_;
 wire _13052_;
 wire _13053_;
 wire _13054_;
 wire _13055_;
 wire _13056_;
 wire _13057_;
 wire _13058_;
 wire _13059_;
 wire _13060_;
 wire _13061_;
 wire _13062_;
 wire _13063_;
 wire _13064_;
 wire _13065_;
 wire _13066_;
 wire _13067_;
 wire _13068_;
 wire _13069_;
 wire _13070_;
 wire _13071_;
 wire _13072_;
 wire _13073_;
 wire _13074_;
 wire _13075_;
 wire _13076_;
 wire _13077_;
 wire _13078_;
 wire _13079_;
 wire _13080_;
 wire _13081_;
 wire _13082_;
 wire _13083_;
 wire _13084_;
 wire _13085_;
 wire _13086_;
 wire _13087_;
 wire _13088_;
 wire _13089_;
 wire _13090_;
 wire _13091_;
 wire _13092_;
 wire _13093_;
 wire _13094_;
 wire _13095_;
 wire _13096_;
 wire _13097_;
 wire _13098_;
 wire _13099_;
 wire _13100_;
 wire _13101_;
 wire _13102_;
 wire _13103_;
 wire _13104_;
 wire _13105_;
 wire _13106_;
 wire _13107_;
 wire _13108_;
 wire _13109_;
 wire _13110_;
 wire _13111_;
 wire _13112_;
 wire _13113_;
 wire _13114_;
 wire _13115_;
 wire _13116_;
 wire _13117_;
 wire _13118_;
 wire _13119_;
 wire _13120_;
 wire _13121_;
 wire _13122_;
 wire _13123_;
 wire _13124_;
 wire _13125_;
 wire _13126_;
 wire _13127_;
 wire _13128_;
 wire _13129_;
 wire _13130_;
 wire _13131_;
 wire _13132_;
 wire _13133_;
 wire _13134_;
 wire _13135_;
 wire _13136_;
 wire _13137_;
 wire _13138_;
 wire _13139_;
 wire _13140_;
 wire _13141_;
 wire _13142_;
 wire _13143_;
 wire _13144_;
 wire _13145_;
 wire _13146_;
 wire _13147_;
 wire _13148_;
 wire _13149_;
 wire _13150_;
 wire _13151_;
 wire _13152_;
 wire _13153_;
 wire _13154_;
 wire _13155_;
 wire _13156_;
 wire _13157_;
 wire _13158_;
 wire _13159_;
 wire _13160_;
 wire _13161_;
 wire _13162_;
 wire _13163_;
 wire _13164_;
 wire _13165_;
 wire _13166_;
 wire _13167_;
 wire _13168_;
 wire _13169_;
 wire _13170_;
 wire _13171_;
 wire _13172_;
 wire _13173_;
 wire _13174_;
 wire _13175_;
 wire _13176_;
 wire _13177_;
 wire _13178_;
 wire _13179_;
 wire _13180_;
 wire _13181_;
 wire _13182_;
 wire _13183_;
 wire _13184_;
 wire _13185_;
 wire _13186_;
 wire _13187_;
 wire _13188_;
 wire _13189_;
 wire _13190_;
 wire _13191_;
 wire _13192_;
 wire _13193_;
 wire _13194_;
 wire _13195_;
 wire _13196_;
 wire _13197_;
 wire _13198_;
 wire _13199_;
 wire _13200_;
 wire _13201_;
 wire _13202_;
 wire _13203_;
 wire _13204_;
 wire _13205_;
 wire _13206_;
 wire _13207_;
 wire _13208_;
 wire _13209_;
 wire _13210_;
 wire _13211_;
 wire _13212_;
 wire _13213_;
 wire _13214_;
 wire _13215_;
 wire _13216_;
 wire _13217_;
 wire _13218_;
 wire _13219_;
 wire _13220_;
 wire _13221_;
 wire _13222_;
 wire _13223_;
 wire _13224_;
 wire _13225_;
 wire _13226_;
 wire _13227_;
 wire _13228_;
 wire _13229_;
 wire _13230_;
 wire _13231_;
 wire _13232_;
 wire _13233_;
 wire _13234_;
 wire _13235_;
 wire _13236_;
 wire _13237_;
 wire _13238_;
 wire _13239_;
 wire _13240_;
 wire _13241_;
 wire _13242_;
 wire _13243_;
 wire _13244_;
 wire _13245_;
 wire _13246_;
 wire _13247_;
 wire _13248_;
 wire _13249_;
 wire _13250_;
 wire _13251_;
 wire _13252_;
 wire _13253_;
 wire _13254_;
 wire _13255_;
 wire _13256_;
 wire _13257_;
 wire _13258_;
 wire _13259_;
 wire _13260_;
 wire _13261_;
 wire _13262_;
 wire _13263_;
 wire _13264_;
 wire _13265_;
 wire _13266_;
 wire _13267_;
 wire _13268_;
 wire _13269_;
 wire _13270_;
 wire _13271_;
 wire _13272_;
 wire _13273_;
 wire _13274_;
 wire _13275_;
 wire _13276_;
 wire _13277_;
 wire _13278_;
 wire _13279_;
 wire _13280_;
 wire _13281_;
 wire _13282_;
 wire _13283_;
 wire _13284_;
 wire _13285_;
 wire _13286_;
 wire _13287_;
 wire _13288_;
 wire _13289_;
 wire _13290_;
 wire _13291_;
 wire _13292_;
 wire _13293_;
 wire _13294_;
 wire _13295_;
 wire _13296_;
 wire _13297_;
 wire _13298_;
 wire _13299_;
 wire _13300_;
 wire _13301_;
 wire _13302_;
 wire _13303_;
 wire _13304_;
 wire _13305_;
 wire _13306_;
 wire _13307_;
 wire _13308_;
 wire _13309_;
 wire _13310_;
 wire _13311_;
 wire _13312_;
 wire _13313_;
 wire _13314_;
 wire _13315_;
 wire _13316_;
 wire _13317_;
 wire _13318_;
 wire _13319_;
 wire _13320_;
 wire _13321_;
 wire _13322_;
 wire _13323_;
 wire _13324_;
 wire _13325_;
 wire _13326_;
 wire _13327_;
 wire _13328_;
 wire _13329_;
 wire _13330_;
 wire _13331_;
 wire _13332_;
 wire _13333_;
 wire _13334_;
 wire _13335_;
 wire _13336_;
 wire _13337_;
 wire _13338_;
 wire _13339_;
 wire _13340_;
 wire _13341_;
 wire _13342_;
 wire _13343_;
 wire _13344_;
 wire _13345_;
 wire _13346_;
 wire _13347_;
 wire _13348_;
 wire _13349_;
 wire _13350_;
 wire _13351_;
 wire _13352_;
 wire _13353_;
 wire _13354_;
 wire _13355_;
 wire _13356_;
 wire _13357_;
 wire _13358_;
 wire _13359_;
 wire _13360_;
 wire _13361_;
 wire _13362_;
 wire _13363_;
 wire _13364_;
 wire _13365_;
 wire _13366_;
 wire _13367_;
 wire _13368_;
 wire _13369_;
 wire _13370_;
 wire _13371_;
 wire _13372_;
 wire _13373_;
 wire _13374_;
 wire _13375_;
 wire _13376_;
 wire _13377_;
 wire _13378_;
 wire _13379_;
 wire _13380_;
 wire _13381_;
 wire _13382_;
 wire _13383_;
 wire _13384_;
 wire _13385_;
 wire _13386_;
 wire _13387_;
 wire _13388_;
 wire _13389_;
 wire _13390_;
 wire _13391_;
 wire _13392_;
 wire _13393_;
 wire _13394_;
 wire _13395_;
 wire _13396_;
 wire _13397_;
 wire _13398_;
 wire _13399_;
 wire _13400_;
 wire _13401_;
 wire _13402_;
 wire _13403_;
 wire _13404_;
 wire _13405_;
 wire _13406_;
 wire _13407_;
 wire _13408_;
 wire _13409_;
 wire _13410_;
 wire _13411_;
 wire _13412_;
 wire _13413_;
 wire _13414_;
 wire _13415_;
 wire _13416_;
 wire _13417_;
 wire _13418_;
 wire _13419_;
 wire _13420_;
 wire _13421_;
 wire _13422_;
 wire _13423_;
 wire _13424_;
 wire _13425_;
 wire _13426_;
 wire _13427_;
 wire _13428_;
 wire _13429_;
 wire _13430_;
 wire _13431_;
 wire _13432_;
 wire _13433_;
 wire _13434_;
 wire _13435_;
 wire _13436_;
 wire _13437_;
 wire _13438_;
 wire _13439_;
 wire _13440_;
 wire _13441_;
 wire _13442_;
 wire _13443_;
 wire _13444_;
 wire _13445_;
 wire _13446_;
 wire _13447_;
 wire _13448_;
 wire _13449_;
 wire _13450_;
 wire _13451_;
 wire _13452_;
 wire _13453_;
 wire _13454_;
 wire _13455_;
 wire _13456_;
 wire _13457_;
 wire _13458_;
 wire _13459_;
 wire _13460_;
 wire _13461_;
 wire _13462_;
 wire _13463_;
 wire _13464_;
 wire _13465_;
 wire _13466_;
 wire _13467_;
 wire _13468_;
 wire _13469_;
 wire _13470_;
 wire _13471_;
 wire _13472_;
 wire _13473_;
 wire _13474_;
 wire _13475_;
 wire _13476_;
 wire _13477_;
 wire _13478_;
 wire _13479_;
 wire _13480_;
 wire _13481_;
 wire _13482_;
 wire _13483_;
 wire _13484_;
 wire _13485_;
 wire _13486_;
 wire _13487_;
 wire _13488_;
 wire _13489_;
 wire _13490_;
 wire _13491_;
 wire _13492_;
 wire _13493_;
 wire _13494_;
 wire _13495_;
 wire _13496_;
 wire _13497_;
 wire _13498_;
 wire _13499_;
 wire _13500_;
 wire _13501_;
 wire _13502_;
 wire _13503_;
 wire _13504_;
 wire _13505_;
 wire _13506_;
 wire _13507_;
 wire _13508_;
 wire _13509_;
 wire _13510_;
 wire _13511_;
 wire _13512_;
 wire _13513_;
 wire _13514_;
 wire _13515_;
 wire _13516_;
 wire _13517_;
 wire _13518_;
 wire _13519_;
 wire _13520_;
 wire _13521_;
 wire _13522_;
 wire _13523_;
 wire _13524_;
 wire _13525_;
 wire _13526_;
 wire _13527_;
 wire _13528_;
 wire _13529_;
 wire _13530_;
 wire _13531_;
 wire _13532_;
 wire _13533_;
 wire _13534_;
 wire _13535_;
 wire _13536_;
 wire _13537_;
 wire _13538_;
 wire _13539_;
 wire _13540_;
 wire _13541_;
 wire _13542_;
 wire _13543_;
 wire _13544_;
 wire _13545_;
 wire _13546_;
 wire _13547_;
 wire _13548_;
 wire _13549_;
 wire _13550_;
 wire _13551_;
 wire _13552_;
 wire _13553_;
 wire _13554_;
 wire _13555_;
 wire _13556_;
 wire _13557_;
 wire _13558_;
 wire _13559_;
 wire _13560_;
 wire _13561_;
 wire _13562_;
 wire _13563_;
 wire _13564_;
 wire _13565_;
 wire _13566_;
 wire _13567_;
 wire _13568_;
 wire _13569_;
 wire _13570_;
 wire _13571_;
 wire _13572_;
 wire _13573_;
 wire _13574_;
 wire _13575_;
 wire _13576_;
 wire _13577_;
 wire _13578_;
 wire _13579_;
 wire _13580_;
 wire _13581_;
 wire _13582_;
 wire _13583_;
 wire _13584_;
 wire _13585_;
 wire _13586_;
 wire _13587_;
 wire _13588_;
 wire _13589_;
 wire _13590_;
 wire _13591_;
 wire _13592_;
 wire _13593_;
 wire _13594_;
 wire _13595_;
 wire _13596_;
 wire _13597_;
 wire _13598_;
 wire _13599_;
 wire _13600_;
 wire _13601_;
 wire _13602_;
 wire _13603_;
 wire _13604_;
 wire _13605_;
 wire _13606_;
 wire _13607_;
 wire _13608_;
 wire _13609_;
 wire _13610_;
 wire _13611_;
 wire _13612_;
 wire _13613_;
 wire _13614_;
 wire _13615_;
 wire _13616_;
 wire _13617_;
 wire _13618_;
 wire _13619_;
 wire _13620_;
 wire _13621_;
 wire _13622_;
 wire _13623_;
 wire _13624_;
 wire _13625_;
 wire _13626_;
 wire _13627_;
 wire _13628_;
 wire _13629_;
 wire _13630_;
 wire _13631_;
 wire _13632_;
 wire _13633_;
 wire _13634_;
 wire _13635_;
 wire _13636_;
 wire _13637_;
 wire _13638_;
 wire _13639_;
 wire _13640_;
 wire _13641_;
 wire _13642_;
 wire _13643_;
 wire _13644_;
 wire _13645_;
 wire _13646_;
 wire _13647_;
 wire _13648_;
 wire _13649_;
 wire _13650_;
 wire _13651_;
 wire _13652_;
 wire _13653_;
 wire _13654_;
 wire _13655_;
 wire _13656_;
 wire _13657_;
 wire _13658_;
 wire _13659_;
 wire _13660_;
 wire _13661_;
 wire _13662_;
 wire _13663_;
 wire _13664_;
 wire _13665_;
 wire _13666_;
 wire _13667_;
 wire _13668_;
 wire _13669_;
 wire _13670_;
 wire _13671_;
 wire _13672_;
 wire _13673_;
 wire _13674_;
 wire _13675_;
 wire _13676_;
 wire _13677_;
 wire _13678_;
 wire _13679_;
 wire _13680_;
 wire _13681_;
 wire _13682_;
 wire _13683_;
 wire _13684_;
 wire _13685_;
 wire _13686_;
 wire _13687_;
 wire _13688_;
 wire _13689_;
 wire _13690_;
 wire _13691_;
 wire _13692_;
 wire _13693_;
 wire _13694_;
 wire _13695_;
 wire _13696_;
 wire _13697_;
 wire _13698_;
 wire _13699_;
 wire _13700_;
 wire _13701_;
 wire _13702_;
 wire _13703_;
 wire _13704_;
 wire _13705_;
 wire _13706_;
 wire _13707_;
 wire _13708_;
 wire _13709_;
 wire _13710_;
 wire _13711_;
 wire _13712_;
 wire _13713_;
 wire _13714_;
 wire _13715_;
 wire _13716_;
 wire _13717_;
 wire _13718_;
 wire _13719_;
 wire _13720_;
 wire _13721_;
 wire _13722_;
 wire _13723_;
 wire _13724_;
 wire _13725_;
 wire _13726_;
 wire _13727_;
 wire _13728_;
 wire _13729_;
 wire _13730_;
 wire _13731_;
 wire _13732_;
 wire _13733_;
 wire _13734_;
 wire _13735_;
 wire _13736_;
 wire _13737_;
 wire _13738_;
 wire _13739_;
 wire _13740_;
 wire _13741_;
 wire _13742_;
 wire _13743_;
 wire _13744_;
 wire _13745_;
 wire _13746_;
 wire _13747_;
 wire _13748_;
 wire _13749_;
 wire _13750_;
 wire _13751_;
 wire _13752_;
 wire _13753_;
 wire _13754_;
 wire _13755_;
 wire _13756_;
 wire _13757_;
 wire _13758_;
 wire _13759_;
 wire _13760_;
 wire _13761_;
 wire _13762_;
 wire _13763_;
 wire _13764_;
 wire _13765_;
 wire _13766_;
 wire _13767_;
 wire _13768_;
 wire _13769_;
 wire _13770_;
 wire _13771_;
 wire _13772_;
 wire _13773_;
 wire _13774_;
 wire _13775_;
 wire _13776_;
 wire _13777_;
 wire _13778_;
 wire _13779_;
 wire _13780_;
 wire _13781_;
 wire _13782_;
 wire _13783_;
 wire _13784_;
 wire _13785_;
 wire _13786_;
 wire _13787_;
 wire _13788_;
 wire _13789_;
 wire _13790_;
 wire _13791_;
 wire _13792_;
 wire _13793_;
 wire _13794_;
 wire _13795_;
 wire _13796_;
 wire _13797_;
 wire _13798_;
 wire _13799_;
 wire _13800_;
 wire _13801_;
 wire _13802_;
 wire _13803_;
 wire _13804_;
 wire _13805_;
 wire _13806_;
 wire _13807_;
 wire _13808_;
 wire _13809_;
 wire _13810_;
 wire _13811_;
 wire _13812_;
 wire _13813_;
 wire _13814_;
 wire _13815_;
 wire _13816_;
 wire _13817_;
 wire _13818_;
 wire _13819_;
 wire _13820_;
 wire _13821_;
 wire _13822_;
 wire _13823_;
 wire _13824_;
 wire _13825_;
 wire _13826_;
 wire _13827_;
 wire _13828_;
 wire _13829_;
 wire _13830_;
 wire _13831_;
 wire _13832_;
 wire _13833_;
 wire _13834_;
 wire _13835_;
 wire _13836_;
 wire _13837_;
 wire _13838_;
 wire _13839_;
 wire _13840_;
 wire _13841_;
 wire _13842_;
 wire _13843_;
 wire _13844_;
 wire _13845_;
 wire _13846_;
 wire _13847_;
 wire _13848_;
 wire _13849_;
 wire _13850_;
 wire _13851_;
 wire _13852_;
 wire _13853_;
 wire _13854_;
 wire _13855_;
 wire _13856_;
 wire _13857_;
 wire _13858_;
 wire _13859_;
 wire _13860_;
 wire _13861_;
 wire _13862_;
 wire _13863_;
 wire _13864_;
 wire _13865_;
 wire _13866_;
 wire _13867_;
 wire _13868_;
 wire _13869_;
 wire _13870_;
 wire _13871_;
 wire _13872_;
 wire _13873_;
 wire _13874_;
 wire _13875_;
 wire _13876_;
 wire _13877_;
 wire _13878_;
 wire _13879_;
 wire _13880_;
 wire _13881_;
 wire _13882_;
 wire _13883_;
 wire _13884_;
 wire _13885_;
 wire _13886_;
 wire _13887_;
 wire _13888_;
 wire _13889_;
 wire _13890_;
 wire _13891_;
 wire _13892_;
 wire _13893_;
 wire _13894_;
 wire _13895_;
 wire _13896_;
 wire _13897_;
 wire _13898_;
 wire _13899_;
 wire _13900_;
 wire _13901_;
 wire _13902_;
 wire _13903_;
 wire _13904_;
 wire _13905_;
 wire _13906_;
 wire _13907_;
 wire _13908_;
 wire _13909_;
 wire _13910_;
 wire _13911_;
 wire _13912_;
 wire _13913_;
 wire _13914_;
 wire _13915_;
 wire _13916_;
 wire _13917_;
 wire _13918_;
 wire _13919_;
 wire _13920_;
 wire _13921_;
 wire _13922_;
 wire _13923_;
 wire _13924_;
 wire _13925_;
 wire _13926_;
 wire _13927_;
 wire _13928_;
 wire _13929_;
 wire _13930_;
 wire _13931_;
 wire _13932_;
 wire _13933_;
 wire _13934_;
 wire _13935_;
 wire _13936_;
 wire _13937_;
 wire _13938_;
 wire _13939_;
 wire _13940_;
 wire _13941_;
 wire _13942_;
 wire _13943_;
 wire _13944_;
 wire _13945_;
 wire _13946_;
 wire _13947_;
 wire _13948_;
 wire _13949_;
 wire _13950_;
 wire _13951_;
 wire _13952_;
 wire _13953_;
 wire _13954_;
 wire _13955_;
 wire _13956_;
 wire _13957_;
 wire _13958_;
 wire _13959_;
 wire _13960_;
 wire _13961_;
 wire _13962_;
 wire _13963_;
 wire _13964_;
 wire _13965_;
 wire _13966_;
 wire _13967_;
 wire _13968_;
 wire _13969_;
 wire _13970_;
 wire _13971_;
 wire _13972_;
 wire _13973_;
 wire _13974_;
 wire _13975_;
 wire _13976_;
 wire _13977_;
 wire _13978_;
 wire _13979_;
 wire _13980_;
 wire _13981_;
 wire _13982_;
 wire _13983_;
 wire _13984_;
 wire _13985_;
 wire _13986_;
 wire _13987_;
 wire _13988_;
 wire _13989_;
 wire _13990_;
 wire _13991_;
 wire _13992_;
 wire _13993_;
 wire _13994_;
 wire _13995_;
 wire _13996_;
 wire _13997_;
 wire _13998_;
 wire _13999_;
 wire _14000_;
 wire _14001_;
 wire _14002_;
 wire _14003_;
 wire _14004_;
 wire _14005_;
 wire _14006_;
 wire _14007_;
 wire _14008_;
 wire _14009_;
 wire _14010_;
 wire _14011_;
 wire _14012_;
 wire _14013_;
 wire _14014_;
 wire _14015_;
 wire _14016_;
 wire _14017_;
 wire _14018_;
 wire _14019_;
 wire _14020_;
 wire _14021_;
 wire _14022_;
 wire _14023_;
 wire _14024_;
 wire _14025_;
 wire _14026_;
 wire _14027_;
 wire _14028_;
 wire _14029_;
 wire _14030_;
 wire _14031_;
 wire _14032_;
 wire _14033_;
 wire _14034_;
 wire _14035_;
 wire _14036_;
 wire _14037_;
 wire _14038_;
 wire _14039_;
 wire _14040_;
 wire _14041_;
 wire _14042_;
 wire _14043_;
 wire _14044_;
 wire _14045_;
 wire _14046_;
 wire _14047_;
 wire _14048_;
 wire _14049_;
 wire _14050_;
 wire _14051_;
 wire _14052_;
 wire _14053_;
 wire _14054_;
 wire _14055_;
 wire _14056_;
 wire _14057_;
 wire _14058_;
 wire _14059_;
 wire _14060_;
 wire _14061_;
 wire _14062_;
 wire _14063_;
 wire _14064_;
 wire _14065_;
 wire _14066_;
 wire _14067_;
 wire _14068_;
 wire _14069_;
 wire _14070_;
 wire _14071_;
 wire _14072_;
 wire _14073_;
 wire _14074_;
 wire _14075_;
 wire _14076_;
 wire _14077_;
 wire _14078_;
 wire _14079_;
 wire _14080_;
 wire _14081_;
 wire _14082_;
 wire _14083_;
 wire _14084_;
 wire _14085_;
 wire _14086_;
 wire _14087_;
 wire _14088_;
 wire _14089_;
 wire _14090_;
 wire _14091_;
 wire _14092_;
 wire _14093_;
 wire _14094_;
 wire _14095_;
 wire _14096_;
 wire _14097_;
 wire _14098_;
 wire _14099_;
 wire _14100_;
 wire _14101_;
 wire _14102_;
 wire _14103_;
 wire _14104_;
 wire _14105_;
 wire _14106_;
 wire _14107_;
 wire _14108_;
 wire _14109_;
 wire _14110_;
 wire _14111_;
 wire _14112_;
 wire _14113_;
 wire _14114_;
 wire _14115_;
 wire _14116_;
 wire _14117_;
 wire _14118_;
 wire _14119_;
 wire _14120_;
 wire _14121_;
 wire _14122_;
 wire _14123_;
 wire _14124_;
 wire _14125_;
 wire _14126_;
 wire _14127_;
 wire _14128_;
 wire _14129_;
 wire _14130_;
 wire _14131_;
 wire _14132_;
 wire _14133_;
 wire _14134_;
 wire _14135_;
 wire _14136_;
 wire _14137_;
 wire _14138_;
 wire _14139_;
 wire _14140_;
 wire _14141_;
 wire _14142_;
 wire _14143_;
 wire _14144_;
 wire _14145_;
 wire _14146_;
 wire _14147_;
 wire _14148_;
 wire _14149_;
 wire _14150_;
 wire _14151_;
 wire _14152_;
 wire _14153_;
 wire _14154_;
 wire _14155_;
 wire _14156_;
 wire _14157_;
 wire _14158_;
 wire _14159_;
 wire _14160_;
 wire _14161_;
 wire _14162_;
 wire _14163_;
 wire _14164_;
 wire _14165_;
 wire _14166_;
 wire _14167_;
 wire _14168_;
 wire _14169_;
 wire _14170_;
 wire _14171_;
 wire _14172_;
 wire _14173_;
 wire _14174_;
 wire _14175_;
 wire _14176_;
 wire _14177_;
 wire _14178_;
 wire _14179_;
 wire _14180_;
 wire _14181_;
 wire _14182_;
 wire _14183_;
 wire _14184_;
 wire _14185_;
 wire _14186_;
 wire _14187_;
 wire _14188_;
 wire _14189_;
 wire _14190_;
 wire _14191_;
 wire _14192_;
 wire _14193_;
 wire _14194_;
 wire _14195_;
 wire _14196_;
 wire _14197_;
 wire _14198_;
 wire _14199_;
 wire _14200_;
 wire _14201_;
 wire _14202_;
 wire _14203_;
 wire _14204_;
 wire _14205_;
 wire _14206_;
 wire _14207_;
 wire _14208_;
 wire _14209_;
 wire _14210_;
 wire _14211_;
 wire _14212_;
 wire _14213_;
 wire _14214_;
 wire _14215_;
 wire _14216_;
 wire _14217_;
 wire _14218_;
 wire _14219_;
 wire _14220_;
 wire _14221_;
 wire _14222_;
 wire _14223_;
 wire _14224_;
 wire _14225_;
 wire _14226_;
 wire _14227_;
 wire _14228_;
 wire _14229_;
 wire _14230_;
 wire _14231_;
 wire _14232_;
 wire _14233_;
 wire _14234_;
 wire _14235_;
 wire _14236_;
 wire _14237_;
 wire _14238_;
 wire _14239_;
 wire _14240_;
 wire _14241_;
 wire _14242_;
 wire _14243_;
 wire _14244_;
 wire _14245_;
 wire _14246_;
 wire _14247_;
 wire _14248_;
 wire _14249_;
 wire _14250_;
 wire _14251_;
 wire _14252_;
 wire _14253_;
 wire _14254_;
 wire _14255_;
 wire _14256_;
 wire _14257_;
 wire _14258_;
 wire _14259_;
 wire _14260_;
 wire _14261_;
 wire _14262_;
 wire _14263_;
 wire _14264_;
 wire _14265_;
 wire _14266_;
 wire _14267_;
 wire _14268_;
 wire _14269_;
 wire _14270_;
 wire _14271_;
 wire _14272_;
 wire _14273_;
 wire _14274_;
 wire _14275_;
 wire _14276_;
 wire _14277_;
 wire _14278_;
 wire _14279_;
 wire _14280_;
 wire _14281_;
 wire _14282_;
 wire _14283_;
 wire _14284_;
 wire _14285_;
 wire _14286_;
 wire _14287_;
 wire _14288_;
 wire _14289_;
 wire _14290_;
 wire _14291_;
 wire _14292_;
 wire _14293_;
 wire _14294_;
 wire _14295_;
 wire _14296_;
 wire _14297_;
 wire _14298_;
 wire _14299_;
 wire _14300_;
 wire _14301_;
 wire _14302_;
 wire _14303_;
 wire _14304_;
 wire _14305_;
 wire _14306_;
 wire _14307_;
 wire _14308_;
 wire _14309_;
 wire _14310_;
 wire _14311_;
 wire _14312_;
 wire _14313_;
 wire _14314_;
 wire _14315_;
 wire _14316_;
 wire _14317_;
 wire _14318_;
 wire _14319_;
 wire _14320_;
 wire _14321_;
 wire _14322_;
 wire _14323_;
 wire _14324_;
 wire _14325_;
 wire _14326_;
 wire _14327_;
 wire _14328_;
 wire _14329_;
 wire _14330_;
 wire _14331_;
 wire _14332_;
 wire _14333_;
 wire _14334_;
 wire _14335_;
 wire _14336_;
 wire _14337_;
 wire _14338_;
 wire _14339_;
 wire _14340_;
 wire _14341_;
 wire _14342_;
 wire _14343_;
 wire _14344_;
 wire _14345_;
 wire _14346_;
 wire _14347_;
 wire _14348_;
 wire _14349_;
 wire _14350_;
 wire _14351_;
 wire _14352_;
 wire _14353_;
 wire _14354_;
 wire _14355_;
 wire _14356_;
 wire _14357_;
 wire _14358_;
 wire _14359_;
 wire _14360_;
 wire _14361_;
 wire _14362_;
 wire _14363_;
 wire _14364_;
 wire _14365_;
 wire _14366_;
 wire _14367_;
 wire _14368_;
 wire _14369_;
 wire _14370_;
 wire _14371_;
 wire _14372_;
 wire _14373_;
 wire _14374_;
 wire _14375_;
 wire _14376_;
 wire _14377_;
 wire _14378_;
 wire _14379_;
 wire _14380_;
 wire _14381_;
 wire _14382_;
 wire _14383_;
 wire _14384_;
 wire _14385_;
 wire _14386_;
 wire _14387_;
 wire _14388_;
 wire _14389_;
 wire _14390_;
 wire _14391_;
 wire _14392_;
 wire _14393_;
 wire _14394_;
 wire _14395_;
 wire _14396_;
 wire _14397_;
 wire _14398_;
 wire _14399_;
 wire _14400_;
 wire _14401_;
 wire _14402_;
 wire _14403_;
 wire _14404_;
 wire _14405_;
 wire _14406_;
 wire _14407_;
 wire _14408_;
 wire _14409_;
 wire _14410_;
 wire _14411_;
 wire _14412_;
 wire _14413_;
 wire _14414_;
 wire _14415_;
 wire _14416_;
 wire _14417_;
 wire _14418_;
 wire _14419_;
 wire _14420_;
 wire _14421_;
 wire _14422_;
 wire _14423_;
 wire _14424_;
 wire _14425_;
 wire _14426_;
 wire _14427_;
 wire _14428_;
 wire _14429_;
 wire _14430_;
 wire _14431_;
 wire _14432_;
 wire _14433_;
 wire _14434_;
 wire _14435_;
 wire _14436_;
 wire _14437_;
 wire _14438_;
 wire _14439_;
 wire _14440_;
 wire _14441_;
 wire _14442_;
 wire _14443_;
 wire _14444_;
 wire _14445_;
 wire _14446_;
 wire _14447_;
 wire _14448_;
 wire _14449_;
 wire _14450_;
 wire _14451_;
 wire _14452_;
 wire _14453_;
 wire _14454_;
 wire _14455_;
 wire _14456_;
 wire _14457_;
 wire _14458_;
 wire _14459_;
 wire _14460_;
 wire _14461_;
 wire _14462_;
 wire _14463_;
 wire _14464_;
 wire _14465_;
 wire _14466_;
 wire _14467_;
 wire _14468_;
 wire _14469_;
 wire _14470_;
 wire _14471_;
 wire _14472_;
 wire _14473_;
 wire _14474_;
 wire _14475_;
 wire _14476_;
 wire _14477_;
 wire _14478_;
 wire _14479_;
 wire _14480_;
 wire _14481_;
 wire _14482_;
 wire _14483_;
 wire _14484_;
 wire _14485_;
 wire _14486_;
 wire _14487_;
 wire _14488_;
 wire _14489_;
 wire _14490_;
 wire _14491_;
 wire _14492_;
 wire _14493_;
 wire _14494_;
 wire _14495_;
 wire _14496_;
 wire _14497_;
 wire _14498_;
 wire _14499_;
 wire _14500_;
 wire _14501_;
 wire _14502_;
 wire _14503_;
 wire _14504_;
 wire _14505_;
 wire _14506_;
 wire _14507_;
 wire _14508_;
 wire _14509_;
 wire _14510_;
 wire _14511_;
 wire _14512_;
 wire _14513_;
 wire _14514_;
 wire _14515_;
 wire _14516_;
 wire _14517_;
 wire _14518_;
 wire _14519_;
 wire _14520_;
 wire _14521_;
 wire _14522_;
 wire _14523_;
 wire _14524_;
 wire _14525_;
 wire _14526_;
 wire _14527_;
 wire _14528_;
 wire _14529_;
 wire _14530_;
 wire _14531_;
 wire _14532_;
 wire _14533_;
 wire _14534_;
 wire _14535_;
 wire _14536_;
 wire _14537_;
 wire _14538_;
 wire _14539_;
 wire _14540_;
 wire _14541_;
 wire _14542_;
 wire _14543_;
 wire _14544_;
 wire _14545_;
 wire _14546_;
 wire _14547_;
 wire _14548_;
 wire _14549_;
 wire _14550_;
 wire _14551_;
 wire _14552_;
 wire _14553_;
 wire _14554_;
 wire _14555_;
 wire _14556_;
 wire _14557_;
 wire _14558_;
 wire _14559_;
 wire _14560_;
 wire _14561_;
 wire _14562_;
 wire _14563_;
 wire _14564_;
 wire _14565_;
 wire _14566_;
 wire _14567_;
 wire _14568_;
 wire _14569_;
 wire _14570_;
 wire _14571_;
 wire _14572_;
 wire _14573_;
 wire _14574_;
 wire _14575_;
 wire _14576_;
 wire _14577_;
 wire _14578_;
 wire _14579_;
 wire _14580_;
 wire _14581_;
 wire _14582_;
 wire _14583_;
 wire _14584_;
 wire _14585_;
 wire _14586_;
 wire _14587_;
 wire _14588_;
 wire _14589_;
 wire _14590_;
 wire _14591_;
 wire _14592_;
 wire _14593_;
 wire _14594_;
 wire _14595_;
 wire _14596_;
 wire _14597_;
 wire _14598_;
 wire _14599_;
 wire _14600_;
 wire _14601_;
 wire _14602_;
 wire _14603_;
 wire _14604_;
 wire _14605_;
 wire _14606_;
 wire _14607_;
 wire _14608_;
 wire _14609_;
 wire _14610_;
 wire _14611_;
 wire _14612_;
 wire _14613_;
 wire _14614_;
 wire _14615_;
 wire _14616_;
 wire _14617_;
 wire _14618_;
 wire _14619_;
 wire _14620_;
 wire _14621_;
 wire _14622_;
 wire _14623_;
 wire _14624_;
 wire _14625_;
 wire _14626_;
 wire _14627_;
 wire _14628_;
 wire _14629_;
 wire _14630_;
 wire _14631_;
 wire _14632_;
 wire _14633_;
 wire _14634_;
 wire _14635_;
 wire _14636_;
 wire _14637_;
 wire _14638_;
 wire _14639_;
 wire _14640_;
 wire _14641_;
 wire _14642_;
 wire _14643_;
 wire _14644_;
 wire _14645_;
 wire _14646_;
 wire _14647_;
 wire _14648_;
 wire _14649_;
 wire _14650_;
 wire _14651_;
 wire _14652_;
 wire _14653_;
 wire _14654_;
 wire _14655_;
 wire _14656_;
 wire _14657_;
 wire _14658_;
 wire _14659_;
 wire _14660_;
 wire _14661_;
 wire _14662_;
 wire _14663_;
 wire _14664_;
 wire _14665_;
 wire _14666_;
 wire _14667_;
 wire _14668_;
 wire _14669_;
 wire _14670_;
 wire _14671_;
 wire _14672_;
 wire _14673_;
 wire _14674_;
 wire _14675_;
 wire _14676_;
 wire _14677_;
 wire _14678_;
 wire _14679_;
 wire _14680_;
 wire _14681_;
 wire _14682_;
 wire _14683_;
 wire _14684_;
 wire _14685_;
 wire _14686_;
 wire _14687_;
 wire _14688_;
 wire _14689_;
 wire _14690_;
 wire _14691_;
 wire _14692_;
 wire _14693_;
 wire _14694_;
 wire _14695_;
 wire _14696_;
 wire _14697_;
 wire _14698_;
 wire _14699_;
 wire _14700_;
 wire _14701_;
 wire _14702_;
 wire _14703_;
 wire _14704_;
 wire _14705_;
 wire _14706_;
 wire _14707_;
 wire _14708_;
 wire _14709_;
 wire _14710_;
 wire _14711_;
 wire _14712_;
 wire _14713_;
 wire _14714_;
 wire _14715_;
 wire _14716_;
 wire _14717_;
 wire _14718_;
 wire _14719_;
 wire _14720_;
 wire _14721_;
 wire _14722_;
 wire _14723_;
 wire _14724_;
 wire _14725_;
 wire _14726_;
 wire _14727_;
 wire _14728_;
 wire _14729_;
 wire _14730_;
 wire _14731_;
 wire _14732_;
 wire _14733_;
 wire _14734_;
 wire _14735_;
 wire _14736_;
 wire _14737_;
 wire _14738_;
 wire _14739_;
 wire _14740_;
 wire _14741_;
 wire _14742_;
 wire _14743_;
 wire _14744_;
 wire _14745_;
 wire _14746_;
 wire _14747_;
 wire _14748_;
 wire _14749_;
 wire _14750_;
 wire _14751_;
 wire _14752_;
 wire _14753_;
 wire _14754_;
 wire _14755_;
 wire _14756_;
 wire _14757_;
 wire _14758_;
 wire _14759_;
 wire _14760_;
 wire _14761_;
 wire _14762_;
 wire _14763_;
 wire _14764_;
 wire _14765_;
 wire _14766_;
 wire _14767_;
 wire _14768_;
 wire _14769_;
 wire _14770_;
 wire _14771_;
 wire _14772_;
 wire _14773_;
 wire _14774_;
 wire _14775_;
 wire _14776_;
 wire _14777_;
 wire _14778_;
 wire _14779_;
 wire _14780_;
 wire _14781_;
 wire _14782_;
 wire _14783_;
 wire _14784_;
 wire _14785_;
 wire _14786_;
 wire _14787_;
 wire _14788_;
 wire _14789_;
 wire _14790_;
 wire _14791_;
 wire _14792_;
 wire _14793_;
 wire _14794_;
 wire _14795_;
 wire _14796_;
 wire _14797_;
 wire _14798_;
 wire _14799_;
 wire _14800_;
 wire _14801_;
 wire _14802_;
 wire _14803_;
 wire _14804_;
 wire _14805_;
 wire _14806_;
 wire _14807_;
 wire _14808_;
 wire _14809_;
 wire _14810_;
 wire _14811_;
 wire _14812_;
 wire _14813_;
 wire _14814_;
 wire _14815_;
 wire _14816_;
 wire _14817_;
 wire _14818_;
 wire _14819_;
 wire _14820_;
 wire _14821_;
 wire _14822_;
 wire _14823_;
 wire _14824_;
 wire _14825_;
 wire _14826_;
 wire _14827_;
 wire _14828_;
 wire _14829_;
 wire _14830_;
 wire _14831_;
 wire _14832_;
 wire _14833_;
 wire _14834_;
 wire _14835_;
 wire _14836_;
 wire _14837_;
 wire _14838_;
 wire _14839_;
 wire _14840_;
 wire _14841_;
 wire _14842_;
 wire _14843_;
 wire _14844_;
 wire _14845_;
 wire _14846_;
 wire _14847_;
 wire _14848_;
 wire _14849_;
 wire _14850_;
 wire _14851_;
 wire _14852_;
 wire _14853_;
 wire _14854_;
 wire _14855_;
 wire _14856_;
 wire _14857_;
 wire _14858_;
 wire _14859_;
 wire _14860_;
 wire _14861_;
 wire _14862_;
 wire _14863_;
 wire _14864_;
 wire _14865_;
 wire _14866_;
 wire _14867_;
 wire _14868_;
 wire _14869_;
 wire _14870_;
 wire _14871_;
 wire _14872_;
 wire _14873_;
 wire _14874_;
 wire _14875_;
 wire _14876_;
 wire _14877_;
 wire _14878_;
 wire _14879_;
 wire _14880_;
 wire _14881_;
 wire _14882_;
 wire _14883_;
 wire _14884_;
 wire _14885_;
 wire _14886_;
 wire _14887_;
 wire _14888_;
 wire _14889_;
 wire _14890_;
 wire _14891_;
 wire _14892_;
 wire _14893_;
 wire _14894_;
 wire _14895_;
 wire _14896_;
 wire _14897_;
 wire _14898_;
 wire _14899_;
 wire _14900_;
 wire _14901_;
 wire _14902_;
 wire _14903_;
 wire _14904_;
 wire _14905_;
 wire _14906_;
 wire _14907_;
 wire _14908_;
 wire _14909_;
 wire _14910_;
 wire _14911_;
 wire _14912_;
 wire _14913_;
 wire _14914_;
 wire _14915_;
 wire _14916_;
 wire _14917_;
 wire _14918_;
 wire _14919_;
 wire _14920_;
 wire _14921_;
 wire _14922_;
 wire _14923_;
 wire _14924_;
 wire _14925_;
 wire _14926_;
 wire _14927_;
 wire _14928_;
 wire _14929_;
 wire _14930_;
 wire _14931_;
 wire _14932_;
 wire _14933_;
 wire _14934_;
 wire _14935_;
 wire _14936_;
 wire _14937_;
 wire _14938_;
 wire _14939_;
 wire _14940_;
 wire _14941_;
 wire _14942_;
 wire _14943_;
 wire _14944_;
 wire _14945_;
 wire _14946_;
 wire _14947_;
 wire _14948_;
 wire _14949_;
 wire _14950_;
 wire _14951_;
 wire _14952_;
 wire _14953_;
 wire _14954_;
 wire _14955_;
 wire _14956_;
 wire _14957_;
 wire _14958_;
 wire _14959_;
 wire _14960_;
 wire _14961_;
 wire _14962_;
 wire _14963_;
 wire _14964_;
 wire _14965_;
 wire _14966_;
 wire _14967_;
 wire _14968_;
 wire _14969_;
 wire _14970_;
 wire _14971_;
 wire _14972_;
 wire _14973_;
 wire _14974_;
 wire _14975_;
 wire _14976_;
 wire _14977_;
 wire _14978_;
 wire _14979_;
 wire _14980_;
 wire _14981_;
 wire _14982_;
 wire _14983_;
 wire _14984_;
 wire _14985_;
 wire _14986_;
 wire _14987_;
 wire _14988_;
 wire _14989_;
 wire _14990_;
 wire _14991_;
 wire _14992_;
 wire _14993_;
 wire _14994_;
 wire _14995_;
 wire _14996_;
 wire _14997_;
 wire _14998_;
 wire _14999_;
 wire _15000_;
 wire _15001_;
 wire _15002_;
 wire _15003_;
 wire _15004_;
 wire _15005_;
 wire _15006_;
 wire _15007_;
 wire _15008_;
 wire _15009_;
 wire _15010_;
 wire _15011_;
 wire _15012_;
 wire _15013_;
 wire _15014_;
 wire _15015_;
 wire _15016_;
 wire _15017_;
 wire _15018_;
 wire _15019_;
 wire _15020_;
 wire _15021_;
 wire _15022_;
 wire _15023_;
 wire _15024_;
 wire _15025_;
 wire _15026_;
 wire _15027_;
 wire _15028_;
 wire _15029_;
 wire _15030_;
 wire _15031_;
 wire _15032_;
 wire _15033_;
 wire _15034_;
 wire _15035_;
 wire _15036_;
 wire _15037_;
 wire _15038_;
 wire _15039_;
 wire _15040_;
 wire _15041_;
 wire _15042_;
 wire _15043_;
 wire _15044_;
 wire _15045_;
 wire _15046_;
 wire _15047_;
 wire _15048_;
 wire _15049_;
 wire _15050_;
 wire _15051_;
 wire _15052_;
 wire _15053_;
 wire _15054_;
 wire _15055_;
 wire _15056_;
 wire _15057_;
 wire _15058_;
 wire _15059_;
 wire _15060_;
 wire _15061_;
 wire _15062_;
 wire _15063_;
 wire _15064_;
 wire _15065_;
 wire _15066_;
 wire _15067_;
 wire _15068_;
 wire _15069_;
 wire _15070_;
 wire _15071_;
 wire _15072_;
 wire _15073_;
 wire _15074_;
 wire _15075_;
 wire _15076_;
 wire _15077_;
 wire _15078_;
 wire _15079_;
 wire _15080_;
 wire _15081_;
 wire _15082_;
 wire _15083_;
 wire _15084_;
 wire _15085_;
 wire _15086_;
 wire _15087_;
 wire _15088_;
 wire _15089_;
 wire _15090_;
 wire _15091_;
 wire _15092_;
 wire _15093_;
 wire _15094_;
 wire _15095_;
 wire _15096_;
 wire _15097_;
 wire _15098_;
 wire _15099_;
 wire _15100_;
 wire _15101_;
 wire _15102_;
 wire _15103_;
 wire _15104_;
 wire _15105_;
 wire _15106_;
 wire _15107_;
 wire _15108_;
 wire _15109_;
 wire _15110_;
 wire _15111_;
 wire _15112_;
 wire _15113_;
 wire _15114_;
 wire _15115_;
 wire _15116_;
 wire _15117_;
 wire _15118_;
 wire _15119_;
 wire _15120_;
 wire _15121_;
 wire _15122_;
 wire _15123_;
 wire _15124_;
 wire _15125_;
 wire _15126_;
 wire _15127_;
 wire _15128_;
 wire _15129_;
 wire _15130_;
 wire _15131_;
 wire _15132_;
 wire _15133_;
 wire _15134_;
 wire _15135_;
 wire _15136_;
 wire _15137_;
 wire _15138_;
 wire _15139_;
 wire _15140_;
 wire _15141_;
 wire _15142_;
 wire _15143_;
 wire _15144_;
 wire _15145_;
 wire _15146_;
 wire _15147_;
 wire _15148_;
 wire _15149_;
 wire _15150_;
 wire _15151_;
 wire _15152_;
 wire _15153_;
 wire _15154_;
 wire _15155_;
 wire _15156_;
 wire _15157_;
 wire _15158_;
 wire _15159_;
 wire _15160_;
 wire _15161_;
 wire _15162_;
 wire _15163_;
 wire _15164_;
 wire _15165_;
 wire _15166_;
 wire _15167_;
 wire _15168_;
 wire _15169_;
 wire _15170_;
 wire _15171_;
 wire _15172_;
 wire _15173_;
 wire _15174_;
 wire _15175_;
 wire _15176_;
 wire _15177_;
 wire _15178_;
 wire _15179_;
 wire _15180_;
 wire _15181_;
 wire _15182_;
 wire _15183_;
 wire _15184_;
 wire _15185_;
 wire _15186_;
 wire _15187_;
 wire _15188_;
 wire _15189_;
 wire _15190_;
 wire _15191_;
 wire _15192_;
 wire _15193_;
 wire _15194_;
 wire _15195_;
 wire _15196_;
 wire _15197_;
 wire _15198_;
 wire _15199_;
 wire _15200_;
 wire _15201_;
 wire _15202_;
 wire _15203_;
 wire _15204_;
 wire _15205_;
 wire _15206_;
 wire _15207_;
 wire _15208_;
 wire _15209_;
 wire _15210_;
 wire _15211_;
 wire _15212_;
 wire _15213_;
 wire _15214_;
 wire _15215_;
 wire _15216_;
 wire _15217_;
 wire _15218_;
 wire _15219_;
 wire _15220_;
 wire _15221_;
 wire _15222_;
 wire _15223_;
 wire _15224_;
 wire _15225_;
 wire _15226_;
 wire _15227_;
 wire _15228_;
 wire _15229_;
 wire _15230_;
 wire _15231_;
 wire _15232_;
 wire _15233_;
 wire _15234_;
 wire _15235_;
 wire _15236_;
 wire _15237_;
 wire _15238_;
 wire _15239_;
 wire _15240_;
 wire _15241_;
 wire _15242_;
 wire _15243_;
 wire _15244_;
 wire _15245_;
 wire _15246_;
 wire _15247_;
 wire _15248_;
 wire _15249_;
 wire _15250_;
 wire _15251_;
 wire _15252_;
 wire _15253_;
 wire _15254_;
 wire _15255_;
 wire _15256_;
 wire _15257_;
 wire _15258_;
 wire _15259_;
 wire _15260_;
 wire _15261_;
 wire _15262_;
 wire _15263_;
 wire _15264_;
 wire _15265_;
 wire _15266_;
 wire _15267_;
 wire _15268_;
 wire _15269_;
 wire _15270_;
 wire _15271_;
 wire _15272_;
 wire _15273_;
 wire _15274_;
 wire _15275_;
 wire _15276_;
 wire _15277_;
 wire _15278_;
 wire _15279_;
 wire _15280_;
 wire _15281_;
 wire _15282_;
 wire _15283_;
 wire _15284_;
 wire _15285_;
 wire _15286_;
 wire _15287_;
 wire _15288_;
 wire _15289_;
 wire _15290_;
 wire _15291_;
 wire _15292_;
 wire _15293_;
 wire _15294_;
 wire _15295_;
 wire _15296_;
 wire _15297_;
 wire _15298_;
 wire _15299_;
 wire _15300_;
 wire _15301_;
 wire _15302_;
 wire _15303_;
 wire _15304_;
 wire _15305_;
 wire _15306_;
 wire _15307_;
 wire _15308_;
 wire _15309_;
 wire _15310_;
 wire _15311_;
 wire _15312_;
 wire _15313_;
 wire _15314_;
 wire _15315_;
 wire _15316_;
 wire _15317_;
 wire _15318_;
 wire _15319_;
 wire _15320_;
 wire _15321_;
 wire _15322_;
 wire _15323_;
 wire _15324_;
 wire _15325_;
 wire _15326_;
 wire _15327_;
 wire _15328_;
 wire _15329_;
 wire _15330_;
 wire _15331_;
 wire _15332_;
 wire _15333_;
 wire _15334_;
 wire _15335_;
 wire _15336_;
 wire _15337_;
 wire _15338_;
 wire _15339_;
 wire _15340_;
 wire _15341_;
 wire _15342_;
 wire _15343_;
 wire _15344_;
 wire _15345_;
 wire _15346_;
 wire _15347_;
 wire _15348_;
 wire _15349_;
 wire _15350_;
 wire _15351_;
 wire _15352_;
 wire _15353_;
 wire _15354_;
 wire _15355_;
 wire _15356_;
 wire _15357_;
 wire _15358_;
 wire _15359_;
 wire _15360_;
 wire _15361_;
 wire _15362_;
 wire _15363_;
 wire _15364_;
 wire _15365_;
 wire _15366_;
 wire _15367_;
 wire _15368_;
 wire _15369_;
 wire _15370_;
 wire _15371_;
 wire _15372_;
 wire _15373_;
 wire _15374_;
 wire _15375_;
 wire _15376_;
 wire _15377_;
 wire _15378_;
 wire _15379_;
 wire _15380_;
 wire _15381_;
 wire _15382_;
 wire _15383_;
 wire _15384_;
 wire _15385_;
 wire _15386_;
 wire _15387_;
 wire _15388_;
 wire _15389_;
 wire _15390_;
 wire _15391_;
 wire _15392_;
 wire _15393_;
 wire _15394_;
 wire _15395_;
 wire _15396_;
 wire _15397_;
 wire _15398_;
 wire _15399_;
 wire _15400_;
 wire _15401_;
 wire _15402_;
 wire _15403_;
 wire _15404_;
 wire _15405_;
 wire _15406_;
 wire _15407_;
 wire _15408_;
 wire _15409_;
 wire _15410_;
 wire _15411_;
 wire _15412_;
 wire _15413_;
 wire _15414_;
 wire _15415_;
 wire _15416_;
 wire _15417_;
 wire _15418_;
 wire _15419_;
 wire _15420_;
 wire _15421_;
 wire _15422_;
 wire _15423_;
 wire _15424_;
 wire _15425_;
 wire _15426_;
 wire _15427_;
 wire _15428_;
 wire _15429_;
 wire _15430_;
 wire _15431_;
 wire _15432_;
 wire _15433_;
 wire _15434_;
 wire _15435_;
 wire _15436_;
 wire _15437_;
 wire _15438_;
 wire _15439_;
 wire _15440_;
 wire _15441_;
 wire _15442_;
 wire _15443_;
 wire _15444_;
 wire _15445_;
 wire _15446_;
 wire _15447_;
 wire _15448_;
 wire _15449_;
 wire _15450_;
 wire _15451_;
 wire _15452_;
 wire _15453_;
 wire _15454_;
 wire _15455_;
 wire _15456_;
 wire _15457_;
 wire _15458_;
 wire _15459_;
 wire _15460_;
 wire _15461_;
 wire _15462_;
 wire _15463_;
 wire _15464_;
 wire _15465_;
 wire _15466_;
 wire _15467_;
 wire _15468_;
 wire _15469_;
 wire _15470_;
 wire _15471_;
 wire _15472_;
 wire _15473_;
 wire _15474_;
 wire _15475_;
 wire _15476_;
 wire _15477_;
 wire _15478_;
 wire _15479_;
 wire _15480_;
 wire _15481_;
 wire _15482_;
 wire _15483_;
 wire _15484_;
 wire _15485_;
 wire _15486_;
 wire _15487_;
 wire _15488_;
 wire _15489_;
 wire _15490_;
 wire _15491_;
 wire _15492_;
 wire _15493_;
 wire _15494_;
 wire _15495_;
 wire _15496_;
 wire _15497_;
 wire _15498_;
 wire _15499_;
 wire _15500_;
 wire _15501_;
 wire _15502_;
 wire _15503_;
 wire _15504_;
 wire _15505_;
 wire _15506_;
 wire _15507_;
 wire _15508_;
 wire _15509_;
 wire _15510_;
 wire _15511_;
 wire _15512_;
 wire _15513_;
 wire _15514_;
 wire _15515_;
 wire _15516_;
 wire _15517_;
 wire _15518_;
 wire _15519_;
 wire _15520_;
 wire _15521_;
 wire _15522_;
 wire _15523_;
 wire _15524_;
 wire _15525_;
 wire _15526_;
 wire _15527_;
 wire _15528_;
 wire _15529_;
 wire _15530_;
 wire _15531_;
 wire _15532_;
 wire _15533_;
 wire _15534_;
 wire _15535_;
 wire _15536_;
 wire _15537_;
 wire _15538_;
 wire _15539_;
 wire _15540_;
 wire _15541_;
 wire _15542_;
 wire _15543_;
 wire _15544_;
 wire _15545_;
 wire _15546_;
 wire _15547_;
 wire _15548_;
 wire _15549_;
 wire _15550_;
 wire _15551_;
 wire _15552_;
 wire _15553_;
 wire _15554_;
 wire _15555_;
 wire _15556_;
 wire _15557_;
 wire _15558_;
 wire _15559_;
 wire _15560_;
 wire _15561_;
 wire _15562_;
 wire _15563_;
 wire _15564_;
 wire _15565_;
 wire _15566_;
 wire _15567_;
 wire _15568_;
 wire _15569_;
 wire _15570_;
 wire _15571_;
 wire _15572_;
 wire _15573_;
 wire _15574_;
 wire _15575_;
 wire _15576_;
 wire _15577_;
 wire _15578_;
 wire _15579_;
 wire _15580_;
 wire _15581_;
 wire _15582_;
 wire _15583_;
 wire _15584_;
 wire _15585_;
 wire _15586_;
 wire _15587_;
 wire _15588_;
 wire _15589_;
 wire _15590_;
 wire _15591_;
 wire _15592_;
 wire _15593_;
 wire _15594_;
 wire _15595_;
 wire _15596_;
 wire _15597_;
 wire _15598_;
 wire _15599_;
 wire _15600_;
 wire _15601_;
 wire _15602_;
 wire _15603_;
 wire _15604_;
 wire _15605_;
 wire _15606_;
 wire _15607_;
 wire _15608_;
 wire _15609_;
 wire _15610_;
 wire _15611_;
 wire _15612_;
 wire _15613_;
 wire _15614_;
 wire _15615_;
 wire _15616_;
 wire _15617_;
 wire _15618_;
 wire _15619_;
 wire _15620_;
 wire _15621_;
 wire _15622_;
 wire _15623_;
 wire _15624_;
 wire _15625_;
 wire _15626_;
 wire _15627_;
 wire _15628_;
 wire _15629_;
 wire _15630_;
 wire _15631_;
 wire _15632_;
 wire _15633_;
 wire _15634_;
 wire _15635_;
 wire _15636_;
 wire _15637_;
 wire _15638_;
 wire _15639_;
 wire _15640_;
 wire _15641_;
 wire _15642_;
 wire _15643_;
 wire _15644_;
 wire _15645_;
 wire _15646_;
 wire _15647_;
 wire _15648_;
 wire _15649_;
 wire _15650_;
 wire _15651_;
 wire _15652_;
 wire _15653_;
 wire _15654_;
 wire _15655_;
 wire _15656_;
 wire _15657_;
 wire _15658_;
 wire _15659_;
 wire _15660_;
 wire _15661_;
 wire _15662_;
 wire _15663_;
 wire _15664_;
 wire _15665_;
 wire _15666_;
 wire _15667_;
 wire _15668_;
 wire _15669_;
 wire _15670_;
 wire _15671_;
 wire _15672_;
 wire _15673_;
 wire _15674_;
 wire _15675_;
 wire _15676_;
 wire _15677_;
 wire _15678_;
 wire _15679_;
 wire _15680_;
 wire _15681_;
 wire _15682_;
 wire _15683_;
 wire _15684_;
 wire _15685_;
 wire _15686_;
 wire _15687_;
 wire _15688_;
 wire _15689_;
 wire _15690_;
 wire _15691_;
 wire _15692_;
 wire _15693_;
 wire _15694_;
 wire _15695_;
 wire _15696_;
 wire _15697_;
 wire _15698_;
 wire _15699_;
 wire _15700_;
 wire _15701_;
 wire _15702_;
 wire _15703_;
 wire _15704_;
 wire _15705_;
 wire _15706_;
 wire _15707_;
 wire _15708_;
 wire _15709_;
 wire _15710_;
 wire _15711_;
 wire _15712_;
 wire _15713_;
 wire _15714_;
 wire _15715_;
 wire _15716_;
 wire _15717_;
 wire _15718_;
 wire _15719_;
 wire _15720_;
 wire _15721_;
 wire _15722_;
 wire _15723_;
 wire _15724_;
 wire _15725_;
 wire _15726_;
 wire _15727_;
 wire _15728_;
 wire _15729_;
 wire _15730_;
 wire _15731_;
 wire _15732_;
 wire _15733_;
 wire _15734_;
 wire _15735_;
 wire _15736_;
 wire _15737_;
 wire _15738_;
 wire _15739_;
 wire _15740_;
 wire _15741_;
 wire _15742_;
 wire _15743_;
 wire _15744_;
 wire _15745_;
 wire _15746_;
 wire _15747_;
 wire _15748_;
 wire _15749_;
 wire _15750_;
 wire _15751_;
 wire _15752_;
 wire _15753_;
 wire _15754_;
 wire _15755_;
 wire _15756_;
 wire _15757_;
 wire _15758_;
 wire _15759_;
 wire _15760_;
 wire _15761_;
 wire _15762_;
 wire _15763_;
 wire _15764_;
 wire _15765_;
 wire _15766_;
 wire _15767_;
 wire _15768_;
 wire _15769_;
 wire _15770_;
 wire _15771_;
 wire _15772_;
 wire _15773_;
 wire _15774_;
 wire _15775_;
 wire _15776_;
 wire _15777_;
 wire _15778_;
 wire _15779_;
 wire _15780_;
 wire _15781_;
 wire _15782_;
 wire _15783_;
 wire _15784_;
 wire _15785_;
 wire _15786_;
 wire _15787_;
 wire _15788_;
 wire _15789_;
 wire _15790_;
 wire _15791_;
 wire _15792_;
 wire _15793_;
 wire _15794_;
 wire _15795_;
 wire _15796_;
 wire _15797_;
 wire _15798_;
 wire _15799_;
 wire _15800_;
 wire _15801_;
 wire _15802_;
 wire _15803_;
 wire _15804_;
 wire _15805_;
 wire _15806_;
 wire _15807_;
 wire _15808_;
 wire _15809_;
 wire _15810_;
 wire _15811_;
 wire _15812_;
 wire _15813_;
 wire _15814_;
 wire _15815_;
 wire _15816_;
 wire _15817_;
 wire _15818_;
 wire _15819_;
 wire _15820_;
 wire _15821_;
 wire _15822_;
 wire _15823_;
 wire _15824_;
 wire _15825_;
 wire _15826_;
 wire _15827_;
 wire _15828_;
 wire _15829_;
 wire _15830_;
 wire _15831_;
 wire _15832_;
 wire _15833_;
 wire _15834_;
 wire _15835_;
 wire _15836_;
 wire _15837_;
 wire _15838_;
 wire _15839_;
 wire _15840_;
 wire _15841_;
 wire _15842_;
 wire _15843_;
 wire _15844_;
 wire _15845_;
 wire _15846_;
 wire _15847_;
 wire _15848_;
 wire _15849_;
 wire _15850_;
 wire _15851_;
 wire _15852_;
 wire _15853_;
 wire _15854_;
 wire _15855_;
 wire _15856_;
 wire _15857_;
 wire _15858_;
 wire _15859_;
 wire _15860_;
 wire _15861_;
 wire _15862_;
 wire _15863_;
 wire _15864_;
 wire _15865_;
 wire _15866_;
 wire _15867_;
 wire _15868_;
 wire _15869_;
 wire _15870_;
 wire _15871_;
 wire _15872_;
 wire _15873_;
 wire _15874_;
 wire _15875_;
 wire _15876_;
 wire _15877_;
 wire _15878_;
 wire _15879_;
 wire _15880_;
 wire _15881_;
 wire _15882_;
 wire _15883_;
 wire _15884_;
 wire _15885_;
 wire _15886_;
 wire _15887_;
 wire _15888_;
 wire _15889_;
 wire _15890_;
 wire _15891_;
 wire _15892_;
 wire _15893_;
 wire _15894_;
 wire _15895_;
 wire _15896_;
 wire _15897_;
 wire _15898_;
 wire _15899_;
 wire _15900_;
 wire _15901_;
 wire _15902_;
 wire _15903_;
 wire _15904_;
 wire _15905_;
 wire _15906_;
 wire _15907_;
 wire _15908_;
 wire _15909_;
 wire _15910_;
 wire _15911_;
 wire _15912_;
 wire _15913_;
 wire _15914_;
 wire _15915_;
 wire _15916_;
 wire _15917_;
 wire _15918_;
 wire _15919_;
 wire _15920_;
 wire _15921_;
 wire _15922_;
 wire _15923_;
 wire _15924_;
 wire _15925_;
 wire _15926_;
 wire _15927_;
 wire _15928_;
 wire _15929_;
 wire _15930_;
 wire _15931_;
 wire _15932_;
 wire _15933_;
 wire _15934_;
 wire _15935_;
 wire _15936_;
 wire _15937_;
 wire _15938_;
 wire _15939_;
 wire _15940_;
 wire _15941_;
 wire _15942_;
 wire _15943_;
 wire _15944_;
 wire _15945_;
 wire _15946_;
 wire _15947_;
 wire _15948_;
 wire _15949_;
 wire _15950_;
 wire _15951_;
 wire _15952_;
 wire _15953_;
 wire _15954_;
 wire _15955_;
 wire _15956_;
 wire _15957_;
 wire _15958_;
 wire _15959_;
 wire _15960_;
 wire _15961_;
 wire _15962_;
 wire _15963_;
 wire _15964_;
 wire _15965_;
 wire _15966_;
 wire _15967_;
 wire _15968_;
 wire _15969_;
 wire _15970_;
 wire _15971_;
 wire _15972_;
 wire _15973_;
 wire _15974_;
 wire _15975_;
 wire _15976_;
 wire _15977_;
 wire _15978_;
 wire _15979_;
 wire _15980_;
 wire _15981_;
 wire _15982_;
 wire _15983_;
 wire _15984_;
 wire _15985_;
 wire _15986_;
 wire _15987_;
 wire _15988_;
 wire _15989_;
 wire _15990_;
 wire _15991_;
 wire _15992_;
 wire _15993_;
 wire _15994_;
 wire _15995_;
 wire _15996_;
 wire _15997_;
 wire _15998_;
 wire _15999_;
 wire _16000_;
 wire _16001_;
 wire _16002_;
 wire _16003_;
 wire _16004_;
 wire _16005_;
 wire _16006_;
 wire _16007_;
 wire _16008_;
 wire _16009_;
 wire _16010_;
 wire _16011_;
 wire _16012_;
 wire _16013_;
 wire _16014_;
 wire _16015_;
 wire _16016_;
 wire _16017_;
 wire _16018_;
 wire _16019_;
 wire _16020_;
 wire _16021_;
 wire _16022_;
 wire _16023_;
 wire _16024_;
 wire _16025_;
 wire _16026_;
 wire _16027_;
 wire _16028_;
 wire _16029_;
 wire _16030_;
 wire _16031_;
 wire _16032_;
 wire _16033_;
 wire _16034_;
 wire _16035_;
 wire _16036_;
 wire _16037_;
 wire _16038_;
 wire _16039_;
 wire _16040_;
 wire _16041_;
 wire _16042_;
 wire _16043_;
 wire _16044_;
 wire _16045_;
 wire _16046_;
 wire _16047_;
 wire _16048_;
 wire _16049_;
 wire _16050_;
 wire _16051_;
 wire _16052_;
 wire _16053_;
 wire _16054_;
 wire _16055_;
 wire _16056_;
 wire _16057_;
 wire _16058_;
 wire _16059_;
 wire _16060_;
 wire _16061_;
 wire _16062_;
 wire _16063_;
 wire _16064_;
 wire _16065_;
 wire _16066_;
 wire _16067_;
 wire _16068_;
 wire _16069_;
 wire _16070_;
 wire _16071_;
 wire _16072_;
 wire _16073_;
 wire _16074_;
 wire _16075_;
 wire _16076_;
 wire _16077_;
 wire _16078_;
 wire _16079_;
 wire _16080_;
 wire _16081_;
 wire _16082_;
 wire _16083_;
 wire _16084_;
 wire _16085_;
 wire _16086_;
 wire _16087_;
 wire _16088_;
 wire _16089_;
 wire _16090_;
 wire _16091_;
 wire _16092_;
 wire _16093_;
 wire _16094_;
 wire _16095_;
 wire _16096_;
 wire _16097_;
 wire _16098_;
 wire _16099_;
 wire _16100_;
 wire _16101_;
 wire _16102_;
 wire _16103_;
 wire _16104_;
 wire _16105_;
 wire _16106_;
 wire _16107_;
 wire _16108_;
 wire _16109_;
 wire _16110_;
 wire _16111_;
 wire _16112_;
 wire _16113_;
 wire _16114_;
 wire _16115_;
 wire _16116_;
 wire _16117_;
 wire _16118_;
 wire _16119_;
 wire _16120_;
 wire _16121_;
 wire _16122_;
 wire _16123_;
 wire _16124_;
 wire _16125_;
 wire _16126_;
 wire _16127_;
 wire _16128_;
 wire _16129_;
 wire _16130_;
 wire _16131_;
 wire _16132_;
 wire _16133_;
 wire _16134_;
 wire _16135_;
 wire _16136_;
 wire _16137_;
 wire _16138_;
 wire _16139_;
 wire _16140_;
 wire _16141_;
 wire _16142_;
 wire _16143_;
 wire _16144_;
 wire _16145_;
 wire _16146_;
 wire _16147_;
 wire _16148_;
 wire _16149_;
 wire _16150_;
 wire _16151_;
 wire _16152_;
 wire _16153_;
 wire _16154_;
 wire _16155_;
 wire _16156_;
 wire _16157_;
 wire _16158_;
 wire _16159_;
 wire _16160_;
 wire _16161_;
 wire _16162_;
 wire _16163_;
 wire _16164_;
 wire _16165_;
 wire _16166_;
 wire _16167_;
 wire _16168_;
 wire _16169_;
 wire _16170_;
 wire _16171_;
 wire _16172_;
 wire _16173_;
 wire _16174_;
 wire _16175_;
 wire _16176_;
 wire _16177_;
 wire _16178_;
 wire _16179_;
 wire _16180_;
 wire _16181_;
 wire _16182_;
 wire _16183_;
 wire _16184_;
 wire _16185_;
 wire _16186_;
 wire _16187_;
 wire _16188_;
 wire _16189_;
 wire _16190_;
 wire _16191_;
 wire _16192_;
 wire _16193_;
 wire _16194_;
 wire _16195_;
 wire _16196_;
 wire _16197_;
 wire _16198_;
 wire _16199_;
 wire _16200_;
 wire _16201_;
 wire _16202_;
 wire _16203_;
 wire _16204_;
 wire _16205_;
 wire _16206_;
 wire _16207_;
 wire _16208_;
 wire _16209_;
 wire _16210_;
 wire _16211_;
 wire _16212_;
 wire _16213_;
 wire _16214_;
 wire _16215_;
 wire _16216_;
 wire _16217_;
 wire _16218_;
 wire _16219_;
 wire _16220_;
 wire _16221_;
 wire _16222_;
 wire _16223_;
 wire _16224_;
 wire _16225_;
 wire _16226_;
 wire _16227_;
 wire _16228_;
 wire _16229_;
 wire _16230_;
 wire _16231_;
 wire _16232_;
 wire _16233_;
 wire _16234_;
 wire _16235_;
 wire _16236_;
 wire _16237_;
 wire _16238_;
 wire _16239_;
 wire _16240_;
 wire _16241_;
 wire _16242_;
 wire _16243_;
 wire _16244_;
 wire _16245_;
 wire _16246_;
 wire _16247_;
 wire _16248_;
 wire _16249_;
 wire _16250_;
 wire _16251_;
 wire _16252_;
 wire _16253_;
 wire _16254_;
 wire _16255_;
 wire _16256_;
 wire _16257_;
 wire _16258_;
 wire _16259_;
 wire _16260_;
 wire _16261_;
 wire _16262_;
 wire _16263_;
 wire _16264_;
 wire _16265_;
 wire _16266_;
 wire _16267_;
 wire _16268_;
 wire _16269_;
 wire _16270_;
 wire _16271_;
 wire _16272_;
 wire _16273_;
 wire _16274_;
 wire _16275_;
 wire _16276_;
 wire _16277_;
 wire _16278_;
 wire _16279_;
 wire _16280_;
 wire _16281_;
 wire _16282_;
 wire _16283_;
 wire _16284_;
 wire _16285_;
 wire _16286_;
 wire _16287_;
 wire _16288_;
 wire _16289_;
 wire _16290_;
 wire _16291_;
 wire _16292_;
 wire _16293_;
 wire _16294_;
 wire _16295_;
 wire _16296_;
 wire _16297_;
 wire _16298_;
 wire _16299_;
 wire _16300_;
 wire _16301_;
 wire _16302_;
 wire _16303_;
 wire _16304_;
 wire _16305_;
 wire _16306_;
 wire _16307_;
 wire _16308_;
 wire _16309_;
 wire _16310_;
 wire _16311_;
 wire _16312_;
 wire _16313_;
 wire _16314_;
 wire _16315_;
 wire _16316_;
 wire _16317_;
 wire _16318_;
 wire _16319_;
 wire _16320_;
 wire _16321_;
 wire _16322_;
 wire _16323_;
 wire _16324_;
 wire _16325_;
 wire _16326_;
 wire _16327_;
 wire _16328_;
 wire _16329_;
 wire _16330_;
 wire _16331_;
 wire _16332_;
 wire _16333_;
 wire _16334_;
 wire _16335_;
 wire _16336_;
 wire _16337_;
 wire _16338_;
 wire _16339_;
 wire _16340_;
 wire _16341_;
 wire _16342_;
 wire _16343_;
 wire _16344_;
 wire _16345_;
 wire _16346_;
 wire _16347_;
 wire _16348_;
 wire _16349_;
 wire _16350_;
 wire _16351_;
 wire _16352_;
 wire _16353_;
 wire _16354_;
 wire _16355_;
 wire _16356_;
 wire _16357_;
 wire _16358_;
 wire _16359_;
 wire _16360_;
 wire _16361_;
 wire _16362_;
 wire _16363_;
 wire _16364_;
 wire _16365_;
 wire _16366_;
 wire _16367_;
 wire _16368_;
 wire _16369_;
 wire _16370_;
 wire _16371_;
 wire _16372_;
 wire _16373_;
 wire _16374_;
 wire _16375_;
 wire _16376_;
 wire _16377_;
 wire _16378_;
 wire _16379_;
 wire _16380_;
 wire _16381_;
 wire _16382_;
 wire _16383_;
 wire _16384_;
 wire _16385_;
 wire _16386_;
 wire _16387_;
 wire _16388_;
 wire _16389_;
 wire _16390_;
 wire _16391_;
 wire _16392_;
 wire _16393_;
 wire _16394_;
 wire _16395_;
 wire _16396_;
 wire _16397_;
 wire _16398_;
 wire _16399_;
 wire _16400_;
 wire _16401_;
 wire _16402_;
 wire _16403_;
 wire _16404_;
 wire _16405_;
 wire _16406_;
 wire _16407_;
 wire _16408_;
 wire _16409_;
 wire _16410_;
 wire _16411_;
 wire _16412_;
 wire _16413_;
 wire _16414_;
 wire _16415_;
 wire _16416_;
 wire _16417_;
 wire _16418_;
 wire _16419_;
 wire _16420_;
 wire _16421_;
 wire _16422_;
 wire _16423_;
 wire _16424_;
 wire _16425_;
 wire _16426_;
 wire _16427_;
 wire _16428_;
 wire _16429_;
 wire _16430_;
 wire _16431_;
 wire _16432_;
 wire _16433_;
 wire _16434_;
 wire _16435_;
 wire _16436_;
 wire _16437_;
 wire _16438_;
 wire _16439_;
 wire _16440_;
 wire _16441_;
 wire _16442_;
 wire _16443_;
 wire _16444_;
 wire _16445_;
 wire _16446_;
 wire _16447_;
 wire _16448_;
 wire _16449_;
 wire _16450_;
 wire _16451_;
 wire _16452_;
 wire _16453_;
 wire _16454_;
 wire _16455_;
 wire _16456_;
 wire _16457_;
 wire _16458_;
 wire _16459_;
 wire _16460_;
 wire _16461_;
 wire _16462_;
 wire _16463_;
 wire _16464_;
 wire _16465_;
 wire _16466_;
 wire _16467_;
 wire _16468_;
 wire _16469_;
 wire _16470_;
 wire _16471_;
 wire _16472_;
 wire _16473_;
 wire _16474_;
 wire _16475_;
 wire _16476_;
 wire _16477_;
 wire _16478_;
 wire _16479_;
 wire _16480_;
 wire _16481_;
 wire _16482_;
 wire _16483_;
 wire _16484_;
 wire _16485_;
 wire _16486_;
 wire _16487_;
 wire _16488_;
 wire _16489_;
 wire _16490_;
 wire _16491_;
 wire _16492_;
 wire _16493_;
 wire _16494_;
 wire _16495_;
 wire _16496_;
 wire _16497_;
 wire _16498_;
 wire _16499_;
 wire _16500_;
 wire _16501_;
 wire _16502_;
 wire _16503_;
 wire _16504_;
 wire _16505_;
 wire _16506_;
 wire _16507_;
 wire _16508_;
 wire _16509_;
 wire _16510_;
 wire _16511_;
 wire _16512_;
 wire _16513_;
 wire _16514_;
 wire _16515_;
 wire _16516_;
 wire _16517_;
 wire _16518_;
 wire _16519_;
 wire _16520_;
 wire _16521_;
 wire _16522_;
 wire _16523_;
 wire _16524_;
 wire _16525_;
 wire _16526_;
 wire _16527_;
 wire _16528_;
 wire _16529_;
 wire _16530_;
 wire _16531_;
 wire _16532_;
 wire _16533_;
 wire _16534_;
 wire _16535_;
 wire _16536_;
 wire _16537_;
 wire _16538_;
 wire _16539_;
 wire _16540_;
 wire _16541_;
 wire _16542_;
 wire _16543_;
 wire _16544_;
 wire _16545_;
 wire _16546_;
 wire _16547_;
 wire _16548_;
 wire _16549_;
 wire _16550_;
 wire _16551_;
 wire _16552_;
 wire _16553_;
 wire _16554_;
 wire _16555_;
 wire _16556_;
 wire _16557_;
 wire _16558_;
 wire _16559_;
 wire _16560_;
 wire _16561_;
 wire _16562_;
 wire _16563_;
 wire _16564_;
 wire _16565_;
 wire _16566_;
 wire _16567_;
 wire _16568_;
 wire _16569_;
 wire _16570_;
 wire _16571_;
 wire _16572_;
 wire _16573_;
 wire _16574_;
 wire _16575_;
 wire _16576_;
 wire _16577_;
 wire _16578_;
 wire _16579_;
 wire _16580_;
 wire _16581_;
 wire _16582_;
 wire _16583_;
 wire _16584_;
 wire _16585_;
 wire _16586_;
 wire _16587_;
 wire _16588_;
 wire _16589_;
 wire _16590_;
 wire _16591_;
 wire _16592_;
 wire _16593_;
 wire _16594_;
 wire _16595_;
 wire _16596_;
 wire _16597_;
 wire _16598_;
 wire _16599_;
 wire _16600_;
 wire _16601_;
 wire _16602_;
 wire _16603_;
 wire _16604_;
 wire _16605_;
 wire _16606_;
 wire _16607_;
 wire _16608_;
 wire _16609_;
 wire _16610_;
 wire _16611_;
 wire _16612_;
 wire _16613_;
 wire _16614_;
 wire _16615_;
 wire _16616_;
 wire _16617_;
 wire _16618_;
 wire _16619_;
 wire _16620_;
 wire _16621_;
 wire _16622_;
 wire _16623_;
 wire _16624_;
 wire _16625_;
 wire _16626_;
 wire _16627_;
 wire _16628_;
 wire _16629_;
 wire _16630_;
 wire _16631_;
 wire _16632_;
 wire _16633_;
 wire _16634_;
 wire _16635_;
 wire _16636_;
 wire _16637_;
 wire _16638_;
 wire _16639_;
 wire _16640_;
 wire _16641_;
 wire _16642_;
 wire _16643_;
 wire _16644_;
 wire _16645_;
 wire _16646_;
 wire _16647_;
 wire _16648_;
 wire _16649_;
 wire _16650_;
 wire _16651_;
 wire _16652_;
 wire _16653_;
 wire _16654_;
 wire _16655_;
 wire _16656_;
 wire _16657_;
 wire _16658_;
 wire _16659_;
 wire _16660_;
 wire _16661_;
 wire _16662_;
 wire _16663_;
 wire _16664_;
 wire _16665_;
 wire _16666_;
 wire _16667_;
 wire _16668_;
 wire _16669_;
 wire _16670_;
 wire _16671_;
 wire _16672_;
 wire _16673_;
 wire _16674_;
 wire _16675_;
 wire _16676_;
 wire _16677_;
 wire _16678_;
 wire _16679_;
 wire _16680_;
 wire _16681_;
 wire _16682_;
 wire _16683_;
 wire _16684_;
 wire _16685_;
 wire _16686_;
 wire _16687_;
 wire _16688_;
 wire _16689_;
 wire _16690_;
 wire _16691_;
 wire _16692_;
 wire _16693_;
 wire _16694_;
 wire _16695_;
 wire _16696_;
 wire _16697_;
 wire _16698_;
 wire _16699_;
 wire _16700_;
 wire _16701_;
 wire _16702_;
 wire _16703_;
 wire _16704_;
 wire _16705_;
 wire _16706_;
 wire _16707_;
 wire _16708_;
 wire _16709_;
 wire _16710_;
 wire _16711_;
 wire _16712_;
 wire _16713_;
 wire _16714_;
 wire _16715_;
 wire _16716_;
 wire _16717_;
 wire _16718_;
 wire _16719_;
 wire _16720_;
 wire _16721_;
 wire _16722_;
 wire _16723_;
 wire _16724_;
 wire _16725_;
 wire _16726_;
 wire _16727_;
 wire _16728_;
 wire _16729_;
 wire _16730_;
 wire _16731_;
 wire _16732_;
 wire _16733_;
 wire _16734_;
 wire _16735_;
 wire _16736_;
 wire _16737_;
 wire _16738_;
 wire _16739_;
 wire _16740_;
 wire _16741_;
 wire _16742_;
 wire _16743_;
 wire _16744_;
 wire _16745_;
 wire _16746_;
 wire _16747_;
 wire _16748_;
 wire _16749_;
 wire _16750_;
 wire _16751_;
 wire _16752_;
 wire _16753_;
 wire _16754_;
 wire _16755_;
 wire _16756_;
 wire _16757_;
 wire _16758_;
 wire _16759_;
 wire _16760_;
 wire _16761_;
 wire _16762_;
 wire _16763_;
 wire _16764_;
 wire _16765_;
 wire _16766_;
 wire _16767_;
 wire _16768_;
 wire _16769_;
 wire _16770_;
 wire _16771_;
 wire _16772_;
 wire _16773_;
 wire _16774_;
 wire _16775_;
 wire _16776_;
 wire _16777_;
 wire _16778_;
 wire _16779_;
 wire _16780_;
 wire _16781_;
 wire _16782_;
 wire _16783_;
 wire _16784_;
 wire _16785_;
 wire _16786_;
 wire _16787_;
 wire _16788_;
 wire _16789_;
 wire _16790_;
 wire _16791_;
 wire _16792_;
 wire _16793_;
 wire _16794_;
 wire _16795_;
 wire _16796_;
 wire _16797_;
 wire _16798_;
 wire _16799_;
 wire _16800_;
 wire _16801_;
 wire _16802_;
 wire _16803_;
 wire _16804_;
 wire _16805_;
 wire _16806_;
 wire _16807_;
 wire _16808_;
 wire _16809_;
 wire _16810_;
 wire _16811_;
 wire _16812_;
 wire _16813_;
 wire _16814_;
 wire _16815_;
 wire _16816_;
 wire _16817_;
 wire _16818_;
 wire _16819_;
 wire _16820_;
 wire _16821_;
 wire _16822_;
 wire _16823_;
 wire _16824_;
 wire _16825_;
 wire _16826_;
 wire _16827_;
 wire _16828_;
 wire _16829_;
 wire _16830_;
 wire _16831_;
 wire _16832_;
 wire _16833_;
 wire _16834_;
 wire _16835_;
 wire _16836_;
 wire _16837_;
 wire _16838_;
 wire _16839_;
 wire _16840_;
 wire _16841_;
 wire _16842_;
 wire _16843_;
 wire _16844_;
 wire _16845_;
 wire _16846_;
 wire _16847_;
 wire _16848_;
 wire _16849_;
 wire _16850_;
 wire _16851_;
 wire _16852_;
 wire _16853_;
 wire _16854_;
 wire _16855_;
 wire _16856_;
 wire _16857_;
 wire _16858_;
 wire _16859_;
 wire _16860_;
 wire _16861_;
 wire _16862_;
 wire _16863_;
 wire _16864_;
 wire _16865_;
 wire _16866_;
 wire _16867_;
 wire _16868_;
 wire _16869_;
 wire _16870_;
 wire _16871_;
 wire _16872_;
 wire _16873_;
 wire _16874_;
 wire _16875_;
 wire _16876_;
 wire _16877_;
 wire _16878_;
 wire _16879_;
 wire _16880_;
 wire _16881_;
 wire _16882_;
 wire _16883_;
 wire _16884_;
 wire _16885_;
 wire _16886_;
 wire _16887_;
 wire _16888_;
 wire _16889_;
 wire _16890_;
 wire _16891_;
 wire _16892_;
 wire _16893_;
 wire _16894_;
 wire _16895_;
 wire _16896_;
 wire _16897_;
 wire _16898_;
 wire _16899_;
 wire _16900_;
 wire _16901_;
 wire _16902_;
 wire _16903_;
 wire _16904_;
 wire _16905_;
 wire _16906_;
 wire _16907_;
 wire _16908_;
 wire _16909_;
 wire _16910_;
 wire _16911_;
 wire _16912_;
 wire _16913_;
 wire _16914_;
 wire _16915_;
 wire _16916_;
 wire _16917_;
 wire _16918_;
 wire _16919_;
 wire _16920_;
 wire _16921_;
 wire _16922_;
 wire _16923_;
 wire _16924_;
 wire _16925_;
 wire _16926_;
 wire _16927_;
 wire _16928_;
 wire _16929_;
 wire _16930_;
 wire _16931_;
 wire _16932_;
 wire _16933_;
 wire _16934_;
 wire _16935_;
 wire _16936_;
 wire _16937_;
 wire _16938_;
 wire _16939_;
 wire _16940_;
 wire _16941_;
 wire _16942_;
 wire _16943_;
 wire _16944_;
 wire _16945_;
 wire _16946_;
 wire _16947_;
 wire _16948_;
 wire _16949_;
 wire _16950_;
 wire _16951_;
 wire _16952_;
 wire _16953_;
 wire _16954_;
 wire _16955_;
 wire _16956_;
 wire _16957_;
 wire _16958_;
 wire _16959_;
 wire _16960_;
 wire _16961_;
 wire _16962_;
 wire _16963_;
 wire _16964_;
 wire _16965_;
 wire _16966_;
 wire _16967_;
 wire _16968_;
 wire _16969_;
 wire _16970_;
 wire _16971_;
 wire _16972_;
 wire _16973_;
 wire _16974_;
 wire _16975_;
 wire _16976_;
 wire _16977_;
 wire _16978_;
 wire _16979_;
 wire _16980_;
 wire _16981_;
 wire _16982_;
 wire _16983_;
 wire _16984_;
 wire _16985_;
 wire _16986_;
 wire _16987_;
 wire _16988_;
 wire _16989_;
 wire _16990_;
 wire _16991_;
 wire _16992_;
 wire _16993_;
 wire _16994_;
 wire _16995_;
 wire _16996_;
 wire _16997_;
 wire _16998_;
 wire _16999_;
 wire _17000_;
 wire _17001_;
 wire _17002_;
 wire _17003_;
 wire _17004_;
 wire _17005_;
 wire _17006_;
 wire _17007_;
 wire _17008_;
 wire _17009_;
 wire _17010_;
 wire _17011_;
 wire _17012_;
 wire _17013_;
 wire _17014_;
 wire _17015_;
 wire _17016_;
 wire _17017_;
 wire _17018_;
 wire _17019_;
 wire _17020_;
 wire _17021_;
 wire _17022_;
 wire _17023_;
 wire _17024_;
 wire _17025_;
 wire _17026_;
 wire _17027_;
 wire _17028_;
 wire _17029_;
 wire _17030_;
 wire _17031_;
 wire _17032_;
 wire _17033_;
 wire _17034_;
 wire _17035_;
 wire _17036_;
 wire _17037_;
 wire _17038_;
 wire _17039_;
 wire _17040_;
 wire _17041_;
 wire _17042_;
 wire _17043_;
 wire _17044_;
 wire _17045_;
 wire _17046_;
 wire _17047_;
 wire _17048_;
 wire _17049_;
 wire _17050_;
 wire _17051_;
 wire _17052_;
 wire _17053_;
 wire _17054_;
 wire _17055_;
 wire _17056_;
 wire _17057_;
 wire _17058_;
 wire _17059_;
 wire _17060_;
 wire _17061_;
 wire _17062_;
 wire _17063_;
 wire _17064_;
 wire _17065_;
 wire _17066_;
 wire _17067_;
 wire _17068_;
 wire _17069_;
 wire _17070_;
 wire _17071_;
 wire _17072_;
 wire _17073_;
 wire _17074_;
 wire _17075_;
 wire _17076_;
 wire _17077_;
 wire _17078_;
 wire _17079_;
 wire _17080_;
 wire _17081_;
 wire _17082_;
 wire _17083_;
 wire _17084_;
 wire _17085_;
 wire _17086_;
 wire _17087_;
 wire _17088_;
 wire _17089_;
 wire _17090_;
 wire _17091_;
 wire _17092_;
 wire _17093_;
 wire _17094_;
 wire _17095_;
 wire _17096_;
 wire _17097_;
 wire _17098_;
 wire _17099_;
 wire _17100_;
 wire _17101_;
 wire _17102_;
 wire _17103_;
 wire _17104_;
 wire _17105_;
 wire _17106_;
 wire _17107_;
 wire _17108_;
 wire _17109_;
 wire _17110_;
 wire _17111_;
 wire _17112_;
 wire _17113_;
 wire _17114_;
 wire _17115_;
 wire _17116_;
 wire _17117_;
 wire _17118_;
 wire _17119_;
 wire _17120_;
 wire _17121_;
 wire _17122_;
 wire _17123_;
 wire _17124_;
 wire _17125_;
 wire _17126_;
 wire _17127_;
 wire _17128_;
 wire _17129_;
 wire _17130_;
 wire _17131_;
 wire _17132_;
 wire _17133_;
 wire _17134_;
 wire _17135_;
 wire _17136_;
 wire _17137_;
 wire _17138_;
 wire _17139_;
 wire _17140_;
 wire _17141_;
 wire _17142_;
 wire _17143_;
 wire _17144_;
 wire _17145_;
 wire _17146_;
 wire _17147_;
 wire _17148_;
 wire _17149_;
 wire _17150_;
 wire _17151_;
 wire _17152_;
 wire _17153_;
 wire _17154_;
 wire _17155_;
 wire _17156_;
 wire _17157_;
 wire _17158_;
 wire _17159_;
 wire _17160_;
 wire _17161_;
 wire _17162_;
 wire _17163_;
 wire _17164_;
 wire _17165_;
 wire _17166_;
 wire _17167_;
 wire _17168_;
 wire _17169_;
 wire _17170_;
 wire _17171_;
 wire _17172_;
 wire _17173_;
 wire _17174_;
 wire _17175_;
 wire _17176_;
 wire _17177_;
 wire _17178_;
 wire _17179_;
 wire _17180_;
 wire _17181_;
 wire _17182_;
 wire _17183_;
 wire _17184_;
 wire _17185_;
 wire _17186_;
 wire _17187_;
 wire _17188_;
 wire _17189_;
 wire _17190_;
 wire _17191_;
 wire _17192_;
 wire _17193_;
 wire _17194_;
 wire _17195_;
 wire _17196_;
 wire _17197_;
 wire _17198_;
 wire _17199_;
 wire _17200_;
 wire _17201_;
 wire _17202_;
 wire _17203_;
 wire _17204_;
 wire _17205_;
 wire _17206_;
 wire _17207_;
 wire _17208_;
 wire _17209_;
 wire _17210_;
 wire _17211_;
 wire _17212_;
 wire _17213_;
 wire _17214_;
 wire _17215_;
 wire _17216_;
 wire _17217_;
 wire _17218_;
 wire _17219_;
 wire _17220_;
 wire _17221_;
 wire _17222_;
 wire _17223_;
 wire _17224_;
 wire _17225_;
 wire _17226_;
 wire _17227_;
 wire _17228_;
 wire _17229_;
 wire _17230_;
 wire _17231_;
 wire _17232_;
 wire _17233_;
 wire _17234_;
 wire _17235_;
 wire _17236_;
 wire _17237_;
 wire _17238_;
 wire _17239_;
 wire _17240_;
 wire _17241_;
 wire _17242_;
 wire _17243_;
 wire _17244_;
 wire _17245_;
 wire _17246_;
 wire _17247_;
 wire _17248_;
 wire _17249_;
 wire _17250_;
 wire _17251_;
 wire _17252_;
 wire _17253_;
 wire _17254_;
 wire _17255_;
 wire _17256_;
 wire _17257_;
 wire _17258_;
 wire _17259_;
 wire _17260_;
 wire _17261_;
 wire _17262_;
 wire _17263_;
 wire _17264_;
 wire _17265_;
 wire _17266_;
 wire _17267_;
 wire _17268_;
 wire _17269_;
 wire _17270_;
 wire _17271_;
 wire _17272_;
 wire _17273_;
 wire _17274_;
 wire _17275_;
 wire _17276_;
 wire _17277_;
 wire _17278_;
 wire _17279_;
 wire _17280_;
 wire _17281_;
 wire _17282_;
 wire _17283_;
 wire _17284_;
 wire _17285_;
 wire _17286_;
 wire _17287_;
 wire _17288_;
 wire _17289_;
 wire _17290_;
 wire _17291_;
 wire _17292_;
 wire _17293_;
 wire _17294_;
 wire _17295_;
 wire _17296_;
 wire _17297_;
 wire _17298_;
 wire _17299_;
 wire _17300_;
 wire _17301_;
 wire _17302_;
 wire _17303_;
 wire _17304_;
 wire _17305_;
 wire _17306_;
 wire _17307_;
 wire _17308_;
 wire _17309_;
 wire _17310_;
 wire _17311_;
 wire _17312_;
 wire _17313_;
 wire _17314_;
 wire _17315_;
 wire _17316_;
 wire _17317_;
 wire _17318_;
 wire _17319_;
 wire _17320_;
 wire _17321_;
 wire _17322_;
 wire _17323_;
 wire _17324_;
 wire _17325_;
 wire _17326_;
 wire _17327_;
 wire _17328_;
 wire _17329_;
 wire _17330_;
 wire _17331_;
 wire _17332_;
 wire _17333_;
 wire _17334_;
 wire _17335_;
 wire _17336_;
 wire _17337_;
 wire _17338_;
 wire _17339_;
 wire _17340_;
 wire _17341_;
 wire _17342_;
 wire _17343_;
 wire _17344_;
 wire _17345_;
 wire _17346_;
 wire _17347_;
 wire _17348_;
 wire _17349_;
 wire _17350_;
 wire _17351_;
 wire _17352_;
 wire _17353_;
 wire _17354_;
 wire _17355_;
 wire _17356_;
 wire _17357_;
 wire _17358_;
 wire _17359_;
 wire _17360_;
 wire _17361_;
 wire _17362_;
 wire _17363_;
 wire _17364_;
 wire _17365_;
 wire _17366_;
 wire _17367_;
 wire _17368_;
 wire _17369_;
 wire _17370_;
 wire _17371_;
 wire _17372_;
 wire _17373_;
 wire _17374_;
 wire _17375_;
 wire _17376_;
 wire _17377_;
 wire _17378_;
 wire _17379_;
 wire _17380_;
 wire _17381_;
 wire _17382_;
 wire _17383_;
 wire _17384_;
 wire _17385_;
 wire _17386_;
 wire _17387_;
 wire _17388_;
 wire _17389_;
 wire _17390_;
 wire _17391_;
 wire _17392_;
 wire _17393_;
 wire _17394_;
 wire _17395_;
 wire _17396_;
 wire _17397_;
 wire _17398_;
 wire _17399_;
 wire _17400_;
 wire _17401_;
 wire _17402_;
 wire _17403_;
 wire _17404_;
 wire _17405_;
 wire _17406_;
 wire _17407_;
 wire _17408_;
 wire _17409_;
 wire _17410_;
 wire _17411_;
 wire _17412_;
 wire _17413_;
 wire _17414_;
 wire _17415_;
 wire _17416_;
 wire _17417_;
 wire _17418_;
 wire _17419_;
 wire _17420_;
 wire _17421_;
 wire _17422_;
 wire _17423_;
 wire _17424_;
 wire _17425_;
 wire _17426_;
 wire _17427_;
 wire _17428_;
 wire _17429_;
 wire _17430_;
 wire _17431_;
 wire _17432_;
 wire _17433_;
 wire _17434_;
 wire _17435_;
 wire _17436_;
 wire _17437_;
 wire _17438_;
 wire _17439_;
 wire _17440_;
 wire _17441_;
 wire _17442_;
 wire _17443_;
 wire _17444_;
 wire _17445_;
 wire _17446_;
 wire _17447_;
 wire _17448_;
 wire _17449_;
 wire _17450_;
 wire _17451_;
 wire _17452_;
 wire _17453_;
 wire _17454_;
 wire _17455_;
 wire _17456_;
 wire _17457_;
 wire _17458_;
 wire _17459_;
 wire _17460_;
 wire _17461_;
 wire _17462_;
 wire _17463_;
 wire _17464_;
 wire _17465_;
 wire _17466_;
 wire _17467_;
 wire _17468_;
 wire _17469_;
 wire _17470_;
 wire _17471_;
 wire _17472_;
 wire _17473_;
 wire _17474_;
 wire _17475_;
 wire _17476_;
 wire _17477_;
 wire _17478_;
 wire _17479_;
 wire _17480_;
 wire _17481_;
 wire _17482_;
 wire _17483_;
 wire _17484_;
 wire _17485_;
 wire _17486_;
 wire _17487_;
 wire _17488_;
 wire _17489_;
 wire _17490_;
 wire _17491_;
 wire _17492_;
 wire _17493_;
 wire _17494_;
 wire _17495_;
 wire _17496_;
 wire _17497_;
 wire _17498_;
 wire _17499_;
 wire _17500_;
 wire _17501_;
 wire _17502_;
 wire _17503_;
 wire _17504_;
 wire _17505_;
 wire _17506_;
 wire _17507_;
 wire _17508_;
 wire _17509_;
 wire _17510_;
 wire _17511_;
 wire _17512_;
 wire _17513_;
 wire _17514_;
 wire _17515_;
 wire _17516_;
 wire _17517_;
 wire _17518_;
 wire _17519_;
 wire _17520_;
 wire _17521_;
 wire _17522_;
 wire _17523_;
 wire _17524_;
 wire _17525_;
 wire _17526_;
 wire _17527_;
 wire _17528_;
 wire _17529_;
 wire _17530_;
 wire _17531_;
 wire _17532_;
 wire _17533_;
 wire _17534_;
 wire _17535_;
 wire _17536_;
 wire _17537_;
 wire _17538_;
 wire _17539_;
 wire _17540_;
 wire _17541_;
 wire _17542_;
 wire _17543_;
 wire _17544_;
 wire _17545_;
 wire _17546_;
 wire _17547_;
 wire _17548_;
 wire _17549_;
 wire _17550_;
 wire _17551_;
 wire _17552_;
 wire _17553_;
 wire _17554_;
 wire _17555_;
 wire _17556_;
 wire _17557_;
 wire _17558_;
 wire _17559_;
 wire _17560_;
 wire _17561_;
 wire _17562_;
 wire _17563_;
 wire _17564_;
 wire _17565_;
 wire _17566_;
 wire _17567_;
 wire _17568_;
 wire _17569_;
 wire _17570_;
 wire _17571_;
 wire _17572_;
 wire _17573_;
 wire _17574_;
 wire _17575_;
 wire _17576_;
 wire _17577_;
 wire _17578_;
 wire _17579_;
 wire _17580_;
 wire _17581_;
 wire _17582_;
 wire _17583_;
 wire _17584_;
 wire _17585_;
 wire _17586_;
 wire _17587_;
 wire _17588_;
 wire _17589_;
 wire _17590_;
 wire _17591_;
 wire _17592_;
 wire _17593_;
 wire _17594_;
 wire _17595_;
 wire _17596_;
 wire _17597_;
 wire _17598_;
 wire _17599_;
 wire _17600_;
 wire _17601_;
 wire _17602_;
 wire _17603_;
 wire _17604_;
 wire _17605_;
 wire _17606_;
 wire _17607_;
 wire _17608_;
 wire _17609_;
 wire _17610_;
 wire _17611_;
 wire _17612_;
 wire _17613_;
 wire _17614_;
 wire _17615_;
 wire _17616_;
 wire _17617_;
 wire _17618_;
 wire _17619_;
 wire _17620_;
 wire _17621_;
 wire _17622_;
 wire _17623_;
 wire _17624_;
 wire _17625_;
 wire _17626_;
 wire _17627_;
 wire _17628_;
 wire _17629_;
 wire _17630_;
 wire _17631_;
 wire _17632_;
 wire _17633_;
 wire _17634_;
 wire _17635_;
 wire _17636_;
 wire _17637_;
 wire _17638_;
 wire _17639_;
 wire _17640_;
 wire _17641_;
 wire _17642_;
 wire _17643_;
 wire _17644_;
 wire _17645_;
 wire _17646_;
 wire _17647_;
 wire _17648_;
 wire _17649_;
 wire _17650_;
 wire _17651_;
 wire _17652_;
 wire _17653_;
 wire _17654_;
 wire _17655_;
 wire _17656_;
 wire _17657_;
 wire _17658_;
 wire _17659_;
 wire _17660_;
 wire _17661_;
 wire _17662_;
 wire _17663_;
 wire _17664_;
 wire _17665_;
 wire _17666_;
 wire _17667_;
 wire _17668_;
 wire _17669_;
 wire _17670_;
 wire _17671_;
 wire _17672_;
 wire _17673_;
 wire _17674_;
 wire _17675_;
 wire _17676_;
 wire _17677_;
 wire _17678_;
 wire _17679_;
 wire _17680_;
 wire _17681_;
 wire _17682_;
 wire _17683_;
 wire _17684_;
 wire _17685_;
 wire _17686_;
 wire _17687_;
 wire _17688_;
 wire _17689_;
 wire _17690_;
 wire _17691_;
 wire _17692_;
 wire _17693_;
 wire _17694_;
 wire _17695_;
 wire _17696_;
 wire _17697_;
 wire _17698_;
 wire _17699_;
 wire _17700_;
 wire _17701_;
 wire _17702_;
 wire _17703_;
 wire _17704_;
 wire _17705_;
 wire _17706_;
 wire _17707_;
 wire _17708_;
 wire _17709_;
 wire _17710_;
 wire _17711_;
 wire _17712_;
 wire _17713_;
 wire _17714_;
 wire _17715_;
 wire _17716_;
 wire _17717_;
 wire _17718_;
 wire _17719_;
 wire _17720_;
 wire _17721_;
 wire _17722_;
 wire _17723_;
 wire _17724_;
 wire _17725_;
 wire _17726_;
 wire _17727_;
 wire _17728_;
 wire _17729_;
 wire _17730_;
 wire _17731_;
 wire _17732_;
 wire _17733_;
 wire _17734_;
 wire _17735_;
 wire _17736_;
 wire _17737_;
 wire _17738_;
 wire _17739_;
 wire _17740_;
 wire _17741_;
 wire _17742_;
 wire _17743_;
 wire _17744_;
 wire _17745_;
 wire _17746_;
 wire _17747_;
 wire _17748_;
 wire _17749_;
 wire _17750_;
 wire _17751_;
 wire _17752_;
 wire _17753_;
 wire _17754_;
 wire _17755_;
 wire _17756_;
 wire _17757_;
 wire _17758_;
 wire _17759_;
 wire _17760_;
 wire _17761_;
 wire _17762_;
 wire _17763_;
 wire _17764_;
 wire _17765_;
 wire _17766_;
 wire _17767_;
 wire _17768_;
 wire _17769_;
 wire _17770_;
 wire _17771_;
 wire _17772_;
 wire _17773_;
 wire _17774_;
 wire _17775_;
 wire _17776_;
 wire _17777_;
 wire _17778_;
 wire _17779_;
 wire _17780_;
 wire _17781_;
 wire _17782_;
 wire _17783_;
 wire _17784_;
 wire _17785_;
 wire _17786_;
 wire _17787_;
 wire _17788_;
 wire _17789_;
 wire _17790_;
 wire _17791_;
 wire _17792_;
 wire _17793_;
 wire _17794_;
 wire _17795_;
 wire _17796_;
 wire _17797_;
 wire _17798_;
 wire _17799_;
 wire _17800_;
 wire _17801_;
 wire _17802_;
 wire _17803_;
 wire _17804_;
 wire _17805_;
 wire _17806_;
 wire _17807_;
 wire _17808_;
 wire _17809_;
 wire _17810_;
 wire _17811_;
 wire _17812_;
 wire _17813_;
 wire _17814_;
 wire _17815_;
 wire _17816_;
 wire _17817_;
 wire _17818_;
 wire _17819_;
 wire _17820_;
 wire _17821_;
 wire _17822_;
 wire _17823_;
 wire _17824_;
 wire _17825_;
 wire _17826_;
 wire _17827_;
 wire _17828_;
 wire _17829_;
 wire _17830_;
 wire _17831_;
 wire _17832_;
 wire _17833_;
 wire _17834_;
 wire _17835_;
 wire _17836_;
 wire _17837_;
 wire _17838_;
 wire _17839_;
 wire _17840_;
 wire _17841_;
 wire _17842_;
 wire _17843_;
 wire _17844_;
 wire _17845_;
 wire _17846_;
 wire _17847_;
 wire _17848_;
 wire _17849_;
 wire _17850_;
 wire _17851_;
 wire _17852_;
 wire _17853_;
 wire _17854_;
 wire _17855_;
 wire _17856_;
 wire _17857_;
 wire _17858_;
 wire _17859_;
 wire _17860_;
 wire _17861_;
 wire _17862_;
 wire _17863_;
 wire _17864_;
 wire _17865_;
 wire _17866_;
 wire _17867_;
 wire _17868_;
 wire _17869_;
 wire _17870_;
 wire _17871_;
 wire _17872_;
 wire _17873_;
 wire _17874_;
 wire _17875_;
 wire _17876_;
 wire _17877_;
 wire _17878_;
 wire _17879_;
 wire _17880_;
 wire _17881_;
 wire _17882_;
 wire _17883_;
 wire _17884_;
 wire _17885_;
 wire _17886_;
 wire _17887_;
 wire _17888_;
 wire _17889_;
 wire _17890_;
 wire _17891_;
 wire _17892_;
 wire _17893_;
 wire _17894_;
 wire _17895_;
 wire _17896_;
 wire _17897_;
 wire _17898_;
 wire _17899_;
 wire _17900_;
 wire _17901_;
 wire _17902_;
 wire _17903_;
 wire _17904_;
 wire _17905_;
 wire _17906_;
 wire _17907_;
 wire _17908_;
 wire _17909_;
 wire _17910_;
 wire _17911_;
 wire _17912_;
 wire _17913_;
 wire _17914_;
 wire _17915_;
 wire _17916_;
 wire _17917_;
 wire _17918_;
 wire _17919_;
 wire _17920_;
 wire _17921_;
 wire _17922_;
 wire _17923_;
 wire _17924_;
 wire _17925_;
 wire _17926_;
 wire _17927_;
 wire _17928_;
 wire _17929_;
 wire _17930_;
 wire _17931_;
 wire _17932_;
 wire _17933_;
 wire _17934_;
 wire _17935_;
 wire _17936_;
 wire _17937_;
 wire _17938_;
 wire _17939_;
 wire _17940_;
 wire _17941_;
 wire _17942_;
 wire _17943_;
 wire _17944_;
 wire _17945_;
 wire _17946_;
 wire _17947_;
 wire _17948_;
 wire _17949_;
 wire _17950_;
 wire _17951_;
 wire _17952_;
 wire _17953_;
 wire _17954_;
 wire _17955_;
 wire _17956_;
 wire _17957_;
 wire _17958_;
 wire _17959_;
 wire _17960_;
 wire _17961_;
 wire _17962_;
 wire _17963_;
 wire _17964_;
 wire _17965_;
 wire _17966_;
 wire _17967_;
 wire _17968_;
 wire _17969_;
 wire _17970_;
 wire _17971_;
 wire _17972_;
 wire _17973_;
 wire _17974_;
 wire _17975_;
 wire _17976_;
 wire _17977_;
 wire _17978_;
 wire _17979_;
 wire _17980_;
 wire _17981_;
 wire _17982_;
 wire _17983_;
 wire _17984_;
 wire _17985_;
 wire _17986_;
 wire _17987_;
 wire _17988_;
 wire _17989_;
 wire _17990_;
 wire _17991_;
 wire _17992_;
 wire _17993_;
 wire _17994_;
 wire _17995_;
 wire _17996_;
 wire _17997_;
 wire _17998_;
 wire _17999_;
 wire _18000_;
 wire _18001_;
 wire _18002_;
 wire _18003_;
 wire _18004_;
 wire _18005_;
 wire _18006_;
 wire _18007_;
 wire _18008_;
 wire _18009_;
 wire _18010_;
 wire _18011_;
 wire _18012_;
 wire _18013_;
 wire _18014_;
 wire _18015_;
 wire _18016_;
 wire _18017_;
 wire _18018_;
 wire _18019_;
 wire _18020_;
 wire _18021_;
 wire _18022_;
 wire _18023_;
 wire _18024_;
 wire _18025_;
 wire _18026_;
 wire _18027_;
 wire _18028_;
 wire _18029_;
 wire _18030_;
 wire _18031_;
 wire _18032_;
 wire _18033_;
 wire _18034_;
 wire _18035_;
 wire _18036_;
 wire _18037_;
 wire _18038_;
 wire _18039_;
 wire _18040_;
 wire _18041_;
 wire _18042_;
 wire _18043_;
 wire _18044_;
 wire _18045_;
 wire _18046_;
 wire _18047_;
 wire _18048_;
 wire _18049_;
 wire _18050_;
 wire _18051_;
 wire _18052_;
 wire _18053_;
 wire _18054_;
 wire _18055_;
 wire _18056_;
 wire _18057_;
 wire _18058_;
 wire _18059_;
 wire _18060_;
 wire _18061_;
 wire _18062_;
 wire _18063_;
 wire _18064_;
 wire _18065_;
 wire _18066_;
 wire _18067_;
 wire _18068_;
 wire _18069_;
 wire _18070_;
 wire _18071_;
 wire _18072_;
 wire _18073_;
 wire _18074_;
 wire _18075_;
 wire _18076_;
 wire _18077_;
 wire _18078_;
 wire _18079_;
 wire _18080_;
 wire _18081_;
 wire _18082_;
 wire _18083_;
 wire _18084_;
 wire _18085_;
 wire _18086_;
 wire _18087_;
 wire _18088_;
 wire _18089_;
 wire _18090_;
 wire _18091_;
 wire _18092_;
 wire _18093_;
 wire _18094_;
 wire _18095_;
 wire _18096_;
 wire _18097_;
 wire _18098_;
 wire _18099_;
 wire _18100_;
 wire _18101_;
 wire _18102_;
 wire _18103_;
 wire _18104_;
 wire _18105_;
 wire _18106_;
 wire _18107_;
 wire _18108_;
 wire _18109_;
 wire _18110_;
 wire _18111_;
 wire _18112_;
 wire _18113_;
 wire _18114_;
 wire _18115_;
 wire _18116_;
 wire _18117_;
 wire _18118_;
 wire _18119_;
 wire _18120_;
 wire _18121_;
 wire _18122_;
 wire _18123_;
 wire _18124_;
 wire _18125_;
 wire _18126_;
 wire _18127_;
 wire _18128_;
 wire _18129_;
 wire _18130_;
 wire _18131_;
 wire _18132_;
 wire _18133_;
 wire _18134_;
 wire _18135_;
 wire _18136_;
 wire _18137_;
 wire _18138_;
 wire _18139_;
 wire _18140_;
 wire _18141_;
 wire _18142_;
 wire _18143_;
 wire _18144_;
 wire _18145_;
 wire _18146_;
 wire _18147_;
 wire _18148_;
 wire _18149_;
 wire _18150_;
 wire _18151_;
 wire _18152_;
 wire _18153_;
 wire _18154_;
 wire _18155_;
 wire _18156_;
 wire _18157_;
 wire _18158_;
 wire _18159_;
 wire _18160_;
 wire _18161_;
 wire _18162_;
 wire _18163_;
 wire _18164_;
 wire _18165_;
 wire _18166_;
 wire _18167_;
 wire _18168_;
 wire _18169_;
 wire _18170_;
 wire _18171_;
 wire _18172_;
 wire _18173_;
 wire _18174_;
 wire _18175_;
 wire _18176_;
 wire _18177_;
 wire _18178_;
 wire _18179_;
 wire _18180_;
 wire _18181_;
 wire _18182_;
 wire _18183_;
 wire _18184_;
 wire _18185_;
 wire _18186_;
 wire _18187_;
 wire _18188_;
 wire _18189_;
 wire _18190_;
 wire _18191_;
 wire _18192_;
 wire _18193_;
 wire _18194_;
 wire _18195_;
 wire _18196_;
 wire _18197_;
 wire _18198_;
 wire _18199_;
 wire _18200_;
 wire _18201_;
 wire _18202_;
 wire _18203_;
 wire _18204_;
 wire _18205_;
 wire _18206_;
 wire _18207_;
 wire _18208_;
 wire _18209_;
 wire _18210_;
 wire _18211_;
 wire _18212_;
 wire _18213_;
 wire _18214_;
 wire _18215_;
 wire _18216_;
 wire _18217_;
 wire _18218_;
 wire _18219_;
 wire _18220_;
 wire _18221_;
 wire _18222_;
 wire _18223_;
 wire _18224_;
 wire _18225_;
 wire _18226_;
 wire _18227_;
 wire _18228_;
 wire _18229_;
 wire _18230_;
 wire _18231_;
 wire _18232_;
 wire _18233_;
 wire _18234_;
 wire _18235_;
 wire _18236_;
 wire _18237_;
 wire _18238_;
 wire _18239_;
 wire _18240_;
 wire _18241_;
 wire _18242_;
 wire _18243_;
 wire _18244_;
 wire _18245_;
 wire _18246_;
 wire _18247_;
 wire _18248_;
 wire _18249_;
 wire _18250_;
 wire _18251_;
 wire _18252_;
 wire _18253_;
 wire _18254_;
 wire _18255_;
 wire _18256_;
 wire _18257_;
 wire _18258_;
 wire _18259_;
 wire _18260_;
 wire _18261_;
 wire _18262_;
 wire _18263_;
 wire _18264_;
 wire _18265_;
 wire _18266_;
 wire _18267_;
 wire _18268_;
 wire _18269_;
 wire _18270_;
 wire _18271_;
 wire _18272_;
 wire _18273_;
 wire _18274_;
 wire _18275_;
 wire _18276_;
 wire _18277_;
 wire _18278_;
 wire _18279_;
 wire _18280_;
 wire _18281_;
 wire _18282_;
 wire _18283_;
 wire _18284_;
 wire _18285_;
 wire _18286_;
 wire _18287_;
 wire _18288_;
 wire _18289_;
 wire _18290_;
 wire _18291_;
 wire _18292_;
 wire _18293_;
 wire _18294_;
 wire _18295_;
 wire _18296_;
 wire _18297_;
 wire _18298_;
 wire _18299_;
 wire _18300_;
 wire _18301_;
 wire _18302_;
 wire _18303_;
 wire _18304_;
 wire _18305_;
 wire _18306_;
 wire _18307_;
 wire _18308_;
 wire _18309_;
 wire _18310_;
 wire _18311_;
 wire _18312_;
 wire _18313_;
 wire _18314_;
 wire _18315_;
 wire _18316_;
 wire _18317_;
 wire _18318_;
 wire _18319_;
 wire _18320_;
 wire _18321_;
 wire _18322_;
 wire _18323_;
 wire _18324_;
 wire _18325_;
 wire _18326_;
 wire _18327_;
 wire _18328_;
 wire _18329_;
 wire _18330_;
 wire _18331_;
 wire _18332_;
 wire _18333_;
 wire _18334_;
 wire _18335_;
 wire _18336_;
 wire _18337_;
 wire _18338_;
 wire _18339_;
 wire _18340_;
 wire _18341_;
 wire _18342_;
 wire _18343_;
 wire _18344_;
 wire _18345_;
 wire _18346_;
 wire _18347_;
 wire _18348_;
 wire _18349_;
 wire _18350_;
 wire _18351_;
 wire _18352_;
 wire _18353_;
 wire _18354_;
 wire _18355_;
 wire _18356_;
 wire _18357_;
 wire _18358_;
 wire _18359_;
 wire _18360_;
 wire _18361_;
 wire _18362_;
 wire _18363_;
 wire _18364_;
 wire _18365_;
 wire _18366_;
 wire _18367_;
 wire _18368_;
 wire _18369_;
 wire _18370_;
 wire _18371_;
 wire _18372_;
 wire _18373_;
 wire _18374_;
 wire _18375_;
 wire _18376_;
 wire _18377_;
 wire _18378_;
 wire _18379_;
 wire _18380_;
 wire _18381_;
 wire _18382_;
 wire _18383_;
 wire _18384_;
 wire _18385_;
 wire _18386_;
 wire _18387_;
 wire _18388_;
 wire _18389_;
 wire _18390_;
 wire _18391_;
 wire _18392_;
 wire _18393_;
 wire _18394_;
 wire _18395_;
 wire _18396_;
 wire _18397_;
 wire _18398_;
 wire _18399_;
 wire _18400_;
 wire _18401_;
 wire _18402_;
 wire _18403_;
 wire _18404_;
 wire _18405_;
 wire _18406_;
 wire _18407_;
 wire _18408_;
 wire _18409_;
 wire _18410_;
 wire _18411_;
 wire _18412_;
 wire _18413_;
 wire _18414_;
 wire _18415_;
 wire _18416_;
 wire _18417_;
 wire _18418_;
 wire _18419_;
 wire _18420_;
 wire _18421_;
 wire _18422_;
 wire _18423_;
 wire _18424_;
 wire _18425_;
 wire _18426_;
 wire _18427_;
 wire _18428_;
 wire _18429_;
 wire _18430_;
 wire _18431_;
 wire _18432_;
 wire _18433_;
 wire _18434_;
 wire _18435_;
 wire _18436_;
 wire _18437_;
 wire _18438_;
 wire _18439_;
 wire _18440_;
 wire _18441_;
 wire _18442_;
 wire _18443_;
 wire _18444_;
 wire _18445_;
 wire _18446_;
 wire _18447_;
 wire _18448_;
 wire _18449_;
 wire _18450_;
 wire _18451_;
 wire _18452_;
 wire _18453_;
 wire _18454_;
 wire _18455_;
 wire _18456_;
 wire _18457_;
 wire _18458_;
 wire _18459_;
 wire _18460_;
 wire _18461_;
 wire _18462_;
 wire _18463_;
 wire _18464_;
 wire _18465_;
 wire _18466_;
 wire _18467_;
 wire _18468_;
 wire _18469_;
 wire _18470_;
 wire _18471_;
 wire _18472_;
 wire _18473_;
 wire _18474_;
 wire _18475_;
 wire _18476_;
 wire _18477_;
 wire _18478_;
 wire _18479_;
 wire _18480_;
 wire _18481_;
 wire _18482_;
 wire _18483_;
 wire _18484_;
 wire _18485_;
 wire _18486_;
 wire _18487_;
 wire _18488_;
 wire _18489_;
 wire _18490_;
 wire _18491_;
 wire _18492_;
 wire _18493_;
 wire _18494_;
 wire _18495_;
 wire _18496_;
 wire _18497_;
 wire _18498_;
 wire _18499_;
 wire _18500_;
 wire _18501_;
 wire _18502_;
 wire _18503_;
 wire _18504_;
 wire _18505_;
 wire _18506_;
 wire _18507_;
 wire _18508_;
 wire _18509_;
 wire _18510_;
 wire _18511_;
 wire _18512_;
 wire _18513_;
 wire _18514_;
 wire _18515_;
 wire _18516_;
 wire _18517_;
 wire _18518_;
 wire _18519_;
 wire _18520_;
 wire _18521_;
 wire _18522_;
 wire _18523_;
 wire _18524_;
 wire _18525_;
 wire _18526_;
 wire _18527_;
 wire _18528_;
 wire _18529_;
 wire _18530_;
 wire _18531_;
 wire _18532_;
 wire _18533_;
 wire _18534_;
 wire _18535_;
 wire _18536_;
 wire _18537_;
 wire _18538_;
 wire _18539_;
 wire _18540_;
 wire _18541_;
 wire _18542_;
 wire _18543_;
 wire _18544_;
 wire _18545_;
 wire _18546_;
 wire _18547_;
 wire _18548_;
 wire _18549_;
 wire _18550_;
 wire _18551_;
 wire _18552_;
 wire _18553_;
 wire _18554_;
 wire _18555_;
 wire _18556_;
 wire _18557_;
 wire _18558_;
 wire _18559_;
 wire _18560_;
 wire _18561_;
 wire _18562_;
 wire _18563_;
 wire _18564_;
 wire _18565_;
 wire _18566_;
 wire _18567_;
 wire _18568_;
 wire _18569_;
 wire _18570_;
 wire _18571_;
 wire _18572_;
 wire _18573_;
 wire _18574_;
 wire _18575_;
 wire _18576_;
 wire _18577_;
 wire _18578_;
 wire _18579_;
 wire _18580_;
 wire _18581_;
 wire _18582_;
 wire _18583_;
 wire _18584_;
 wire _18585_;
 wire _18586_;
 wire _18587_;
 wire _18588_;
 wire _18589_;
 wire _18590_;
 wire _18591_;
 wire _18592_;
 wire _18593_;
 wire _18594_;
 wire _18595_;
 wire _18596_;
 wire _18597_;
 wire _18598_;
 wire _18599_;
 wire _18600_;
 wire _18601_;
 wire _18602_;
 wire _18603_;
 wire _18604_;
 wire _18605_;
 wire _18606_;
 wire _18607_;
 wire _18608_;
 wire _18609_;
 wire _18610_;
 wire _18611_;
 wire _18612_;
 wire _18613_;
 wire _18614_;
 wire _18615_;
 wire _18616_;
 wire _18617_;
 wire _18618_;
 wire _18619_;
 wire _18620_;
 wire _18621_;
 wire _18622_;
 wire _18623_;
 wire _18624_;
 wire _18625_;
 wire _18626_;
 wire _18627_;
 wire _18628_;
 wire _18629_;
 wire _18630_;
 wire _18631_;
 wire _18632_;
 wire _18633_;
 wire _18634_;
 wire _18635_;
 wire _18636_;
 wire _18637_;
 wire _18638_;
 wire _18639_;
 wire _18640_;
 wire _18641_;
 wire _18642_;
 wire _18643_;
 wire _18644_;
 wire _18645_;
 wire _18646_;
 wire _18647_;
 wire _18648_;
 wire _18649_;
 wire _18650_;
 wire _18651_;
 wire _18652_;
 wire _18653_;
 wire _18654_;
 wire _18655_;
 wire _18656_;
 wire _18657_;
 wire _18658_;
 wire _18659_;
 wire _18660_;
 wire _18661_;
 wire _18662_;
 wire _18663_;
 wire _18664_;
 wire _18665_;
 wire _18666_;
 wire _18667_;
 wire _18668_;
 wire _18669_;
 wire _18670_;
 wire _18671_;
 wire _18672_;
 wire _18673_;
 wire _18674_;
 wire _18675_;
 wire _18676_;
 wire _18677_;
 wire _18678_;
 wire _18679_;
 wire _18680_;
 wire _18681_;
 wire _18682_;
 wire _18683_;
 wire _18684_;
 wire _18685_;
 wire _18686_;
 wire _18687_;
 wire _18688_;
 wire _18689_;
 wire _18690_;
 wire _18691_;
 wire _18692_;
 wire _18693_;
 wire _18694_;
 wire _18695_;
 wire _18696_;
 wire _18697_;
 wire _18698_;
 wire _18699_;
 wire _18700_;
 wire _18701_;
 wire _18702_;
 wire _18703_;
 wire _18704_;
 wire _18705_;
 wire _18706_;
 wire _18707_;
 wire _18708_;
 wire _18709_;
 wire _18710_;
 wire _18711_;
 wire _18712_;
 wire _18713_;
 wire _18714_;
 wire _18715_;
 wire _18716_;
 wire _18717_;
 wire _18718_;
 wire _18719_;
 wire _18720_;
 wire _18721_;
 wire _18722_;
 wire _18723_;
 wire _18724_;
 wire _18725_;
 wire _18726_;
 wire _18727_;
 wire _18728_;
 wire _18729_;
 wire _18730_;
 wire _18731_;
 wire _18732_;
 wire _18733_;
 wire _18734_;
 wire _18735_;
 wire _18736_;
 wire _18737_;
 wire _18738_;
 wire _18739_;
 wire _18740_;
 wire _18741_;
 wire _18742_;
 wire _18743_;
 wire _18744_;
 wire _18745_;
 wire _18746_;
 wire _18747_;
 wire _18748_;
 wire _18749_;
 wire _18750_;
 wire _18751_;
 wire _18752_;
 wire _18753_;
 wire _18754_;
 wire _18755_;
 wire _18756_;
 wire _18757_;
 wire _18758_;
 wire _18759_;
 wire _18760_;
 wire _18761_;
 wire _18762_;
 wire _18763_;
 wire _18764_;
 wire _18765_;
 wire _18766_;
 wire _18767_;
 wire _18768_;
 wire _18769_;
 wire _18770_;
 wire _18771_;
 wire _18772_;
 wire _18773_;
 wire _18774_;
 wire _18775_;
 wire _18776_;
 wire _18777_;
 wire _18778_;
 wire _18779_;
 wire _18780_;
 wire _18781_;
 wire _18782_;
 wire _18783_;
 wire _18784_;
 wire _18785_;
 wire _18786_;
 wire _18787_;
 wire _18788_;
 wire _18789_;
 wire _18790_;
 wire _18791_;
 wire _18792_;
 wire _18793_;
 wire _18794_;
 wire _18795_;
 wire _18796_;
 wire _18797_;
 wire _18798_;
 wire _18799_;
 wire _18800_;
 wire _18801_;
 wire _18802_;
 wire _18803_;
 wire _18804_;
 wire _18805_;
 wire _18806_;
 wire _18807_;
 wire _18808_;
 wire _18809_;
 wire _18810_;
 wire _18811_;
 wire _18812_;
 wire _18813_;
 wire _18814_;
 wire _18815_;
 wire _18816_;
 wire _18817_;
 wire _18818_;
 wire _18819_;
 wire _18820_;
 wire _18821_;
 wire _18822_;
 wire _18823_;
 wire _18824_;
 wire _18825_;
 wire _18826_;
 wire _18827_;
 wire _18828_;
 wire _18829_;
 wire _18830_;
 wire _18831_;
 wire _18832_;
 wire _18833_;
 wire _18834_;
 wire _18835_;
 wire _18836_;
 wire _18837_;
 wire _18838_;
 wire _18839_;
 wire _18840_;
 wire _18841_;
 wire _18842_;
 wire _18843_;
 wire _18844_;
 wire _18845_;
 wire _18846_;
 wire _18847_;
 wire _18848_;
 wire _18849_;
 wire _18850_;
 wire _18851_;
 wire _18852_;
 wire _18853_;
 wire _18854_;
 wire _18855_;
 wire _18856_;
 wire _18857_;
 wire _18858_;
 wire _18859_;
 wire _18860_;
 wire _18861_;
 wire _18862_;
 wire _18863_;
 wire _18864_;
 wire _18865_;
 wire _18866_;
 wire _18867_;
 wire _18868_;
 wire _18869_;
 wire _18870_;
 wire _18871_;
 wire _18872_;
 wire _18873_;
 wire _18874_;
 wire _18875_;
 wire _18876_;
 wire _18877_;
 wire _18878_;
 wire _18879_;
 wire _18880_;
 wire _18881_;
 wire _18882_;
 wire _18883_;
 wire _18884_;
 wire _18885_;
 wire _18886_;
 wire _18887_;
 wire _18888_;
 wire _18889_;
 wire _18890_;
 wire _18891_;
 wire _18892_;
 wire _18893_;
 wire _18894_;
 wire _18895_;
 wire _18896_;
 wire _18897_;
 wire _18898_;
 wire _18899_;
 wire _18900_;
 wire _18901_;
 wire _18902_;
 wire _18903_;
 wire _18904_;
 wire _18905_;
 wire _18906_;
 wire _18907_;
 wire _18908_;
 wire _18909_;
 wire _18910_;
 wire _18911_;
 wire _18912_;
 wire _18913_;
 wire _18914_;
 wire _18915_;
 wire _18916_;
 wire _18917_;
 wire _18918_;
 wire _18919_;
 wire _18920_;
 wire _18921_;
 wire _18922_;
 wire _18923_;
 wire _18924_;
 wire _18925_;
 wire _18926_;
 wire _18927_;
 wire _18928_;
 wire _18929_;
 wire _18930_;
 wire _18931_;
 wire _18932_;
 wire _18933_;
 wire _18934_;
 wire _18935_;
 wire _18936_;
 wire _18937_;
 wire _18938_;
 wire _18939_;
 wire _18940_;
 wire _18941_;
 wire _18942_;
 wire _18943_;
 wire _18944_;
 wire _18945_;
 wire _18946_;
 wire _18947_;
 wire _18948_;
 wire _18949_;
 wire _18950_;
 wire _18951_;
 wire _18952_;
 wire _18953_;
 wire _18954_;
 wire _18955_;
 wire _18956_;
 wire _18957_;
 wire _18958_;
 wire _18959_;
 wire _18960_;
 wire _18961_;
 wire _18962_;
 wire _18963_;
 wire _18964_;
 wire _18965_;
 wire _18966_;
 wire _18967_;
 wire _18968_;
 wire _18969_;
 wire _18970_;
 wire _18971_;
 wire _18972_;
 wire _18973_;
 wire _18974_;
 wire _18975_;
 wire _18976_;
 wire _18977_;
 wire _18978_;
 wire _18979_;
 wire _18980_;
 wire _18981_;
 wire _18982_;
 wire _18983_;
 wire _18984_;
 wire _18985_;
 wire _18986_;
 wire _18987_;
 wire _18988_;
 wire _18989_;
 wire _18990_;
 wire _18991_;
 wire _18992_;
 wire _18993_;
 wire _18994_;
 wire _18995_;
 wire _18996_;
 wire _18997_;
 wire _18998_;
 wire _18999_;
 wire _19000_;
 wire _19001_;
 wire _19002_;
 wire _19003_;
 wire _19004_;
 wire _19005_;
 wire _19006_;
 wire _19007_;
 wire _19008_;
 wire _19009_;
 wire _19010_;
 wire _19011_;
 wire _19012_;
 wire _19013_;
 wire _19014_;
 wire _19015_;
 wire _19016_;
 wire _19017_;
 wire _19018_;
 wire _19019_;
 wire _19020_;
 wire _19021_;
 wire _19022_;
 wire _19023_;
 wire _19024_;
 wire _19025_;
 wire _19026_;
 wire _19027_;
 wire _19028_;
 wire _19029_;
 wire _19030_;
 wire _19031_;
 wire _19032_;
 wire _19033_;
 wire _19034_;
 wire _19035_;
 wire _19036_;
 wire _19037_;
 wire _19038_;
 wire _19039_;
 wire _19040_;
 wire _19041_;
 wire _19042_;
 wire _19043_;
 wire _19044_;
 wire _19045_;
 wire _19046_;
 wire _19047_;
 wire _19048_;
 wire _19049_;
 wire _19050_;
 wire _19051_;
 wire _19052_;
 wire _19053_;
 wire _19054_;
 wire _19055_;
 wire _19056_;
 wire _19057_;
 wire _19058_;
 wire _19059_;
 wire _19060_;
 wire _19061_;
 wire _19062_;
 wire _19063_;
 wire _19064_;
 wire _19065_;
 wire _19066_;
 wire _19067_;
 wire _19068_;
 wire _19069_;
 wire _19070_;
 wire _19071_;
 wire _19072_;
 wire _19073_;
 wire _19074_;
 wire _19075_;
 wire _19076_;
 wire _19077_;
 wire _19078_;
 wire _19079_;
 wire _19080_;
 wire _19081_;
 wire _19082_;
 wire _19083_;
 wire _19084_;
 wire _19085_;
 wire _19086_;
 wire _19087_;
 wire _19088_;
 wire _19089_;
 wire _19090_;
 wire _19091_;
 wire _19092_;
 wire _19093_;
 wire _19094_;
 wire _19095_;
 wire _19096_;
 wire _19097_;
 wire _19098_;
 wire _19099_;
 wire _19100_;
 wire _19101_;
 wire _19102_;
 wire _19103_;
 wire _19104_;
 wire _19105_;
 wire _19106_;
 wire _19107_;
 wire _19108_;
 wire _19109_;
 wire _19110_;
 wire _19111_;
 wire _19112_;
 wire _19113_;
 wire _19114_;
 wire _19115_;
 wire _19116_;
 wire _19117_;
 wire _19118_;
 wire _19119_;
 wire _19120_;
 wire _19121_;
 wire _19122_;
 wire _19123_;
 wire _19124_;
 wire _19125_;
 wire _19126_;
 wire _19127_;
 wire _19128_;
 wire _19129_;
 wire _19130_;
 wire _19131_;
 wire _19132_;
 wire _19133_;
 wire _19134_;
 wire _19135_;
 wire _19136_;
 wire _19137_;
 wire _19138_;
 wire _19139_;
 wire _19140_;
 wire _19141_;
 wire _19142_;
 wire _19143_;
 wire _19144_;
 wire _19145_;
 wire _19146_;
 wire _19147_;
 wire _19148_;
 wire _19149_;
 wire _19150_;
 wire _19151_;
 wire _19152_;
 wire _19153_;
 wire _19154_;
 wire _19155_;
 wire _19156_;
 wire _19157_;
 wire _19158_;
 wire _19159_;
 wire _19160_;
 wire _19161_;
 wire _19162_;
 wire _19163_;
 wire _19164_;
 wire _19165_;
 wire _19166_;
 wire _19167_;
 wire _19168_;
 wire _19169_;
 wire _19170_;
 wire _19171_;
 wire _19172_;
 wire _19173_;
 wire _19174_;
 wire _19175_;
 wire _19176_;
 wire _19177_;
 wire _19178_;
 wire _19179_;
 wire _19180_;
 wire _19181_;
 wire _19182_;
 wire _19183_;
 wire _19184_;
 wire _19185_;
 wire _19186_;
 wire _19187_;
 wire _19188_;
 wire _19189_;
 wire _19190_;
 wire _19191_;
 wire _19192_;
 wire _19193_;
 wire _19194_;
 wire _19195_;
 wire _19196_;
 wire _19197_;
 wire _19198_;
 wire _19199_;
 wire _19200_;
 wire _19201_;
 wire _19202_;
 wire _19203_;
 wire _19204_;
 wire _19205_;
 wire _19206_;
 wire _19207_;
 wire _19208_;
 wire _19209_;
 wire _19210_;
 wire _19211_;
 wire _19212_;
 wire _19213_;
 wire _19214_;
 wire _19215_;
 wire _19216_;
 wire _19217_;
 wire _19218_;
 wire _19219_;
 wire _19220_;
 wire _19221_;
 wire _19222_;
 wire _19223_;
 wire _19224_;
 wire _19225_;
 wire _19226_;
 wire _19227_;
 wire _19228_;
 wire _19229_;
 wire _19230_;
 wire _19231_;
 wire _19232_;
 wire _19233_;
 wire _19234_;
 wire _19235_;
 wire _19236_;
 wire _19237_;
 wire _19238_;
 wire _19239_;
 wire _19240_;
 wire _19241_;
 wire _19242_;
 wire _19243_;
 wire _19244_;
 wire _19245_;
 wire _19246_;
 wire _19247_;
 wire _19248_;
 wire _19249_;
 wire _19250_;
 wire _19251_;
 wire _19252_;
 wire _19253_;
 wire _19254_;
 wire _19255_;
 wire _19256_;
 wire _19257_;
 wire _19258_;
 wire _19259_;
 wire _19260_;
 wire _19261_;
 wire _19262_;
 wire _19263_;
 wire _19264_;
 wire _19265_;
 wire _19266_;
 wire _19267_;
 wire _19268_;
 wire _19269_;
 wire _19270_;
 wire _19271_;
 wire _19272_;
 wire _19273_;
 wire _19274_;
 wire _19275_;
 wire _19276_;
 wire _19277_;
 wire _19278_;
 wire _19279_;
 wire _19280_;
 wire _19281_;
 wire _19282_;
 wire _19283_;
 wire _19284_;
 wire _19285_;
 wire _19286_;
 wire _19287_;
 wire _19288_;
 wire _19289_;
 wire _19290_;
 wire _19291_;
 wire _19292_;
 wire _19293_;
 wire _19294_;
 wire _19295_;
 wire _19296_;
 wire _19297_;
 wire _19298_;
 wire _19299_;
 wire _19300_;
 wire _19301_;
 wire _19302_;
 wire _19303_;
 wire _19304_;
 wire _19305_;
 wire _19306_;
 wire _19307_;
 wire _19308_;
 wire _19309_;
 wire _19310_;
 wire _19311_;
 wire _19312_;
 wire _19313_;
 wire _19314_;
 wire _19315_;
 wire _19316_;
 wire _19317_;
 wire _19318_;
 wire _19319_;
 wire _19320_;
 wire _19321_;
 wire _19322_;
 wire _19323_;
 wire _19324_;
 wire _19325_;
 wire _19326_;
 wire _19327_;
 wire _19328_;
 wire _19329_;
 wire _19330_;
 wire _19331_;
 wire _19332_;
 wire _19333_;
 wire _19334_;
 wire _19335_;
 wire _19336_;
 wire _19337_;
 wire _19338_;
 wire _19339_;
 wire _19340_;
 wire _19341_;
 wire _19342_;
 wire _19343_;
 wire _19344_;
 wire _19345_;
 wire _19346_;
 wire _19347_;
 wire _19348_;
 wire _19349_;
 wire _19350_;
 wire _19351_;
 wire _19352_;
 wire _19353_;
 wire _19354_;
 wire _19355_;
 wire _19356_;
 wire _19357_;
 wire _19358_;
 wire _19359_;
 wire _19360_;
 wire _19361_;
 wire _19362_;
 wire _19363_;
 wire _19364_;
 wire _19365_;
 wire _19366_;
 wire _19367_;
 wire _19368_;
 wire _19369_;
 wire _19370_;
 wire _19371_;
 wire _19372_;
 wire _19373_;
 wire _19374_;
 wire _19375_;
 wire _19376_;
 wire _19377_;
 wire _19378_;
 wire _19379_;
 wire _19380_;
 wire _19381_;
 wire _19382_;
 wire _19383_;
 wire _19384_;
 wire _19385_;
 wire _19386_;
 wire _19387_;
 wire _19388_;
 wire _19389_;
 wire _19390_;
 wire _19391_;
 wire _19392_;
 wire _19393_;
 wire _19394_;
 wire _19395_;
 wire _19396_;
 wire _19397_;
 wire _19398_;
 wire _19399_;
 wire _19400_;
 wire _19401_;
 wire _19402_;
 wire _19403_;
 wire _19404_;
 wire _19405_;
 wire _19406_;
 wire _19407_;
 wire _19408_;
 wire _19409_;
 wire _19410_;
 wire _19411_;
 wire _19412_;
 wire _19413_;
 wire _19414_;
 wire _19415_;
 wire _19416_;
 wire _19417_;
 wire _19418_;
 wire _19419_;
 wire _19420_;
 wire _19421_;
 wire _19422_;
 wire _19423_;
 wire _19424_;
 wire _19425_;
 wire _19426_;
 wire _19427_;
 wire _19428_;
 wire _19429_;
 wire _19430_;
 wire _19431_;
 wire _19432_;
 wire _19433_;
 wire _19434_;
 wire _19435_;
 wire _19436_;
 wire _19437_;
 wire _19438_;
 wire _19439_;
 wire _19440_;
 wire _19441_;
 wire _19442_;
 wire _19443_;
 wire _19444_;
 wire _19445_;
 wire _19446_;
 wire _19447_;
 wire _19448_;
 wire _19449_;
 wire _19450_;
 wire _19451_;
 wire _19452_;
 wire _19453_;
 wire _19454_;
 wire _19455_;
 wire _19456_;
 wire _19457_;
 wire _19458_;
 wire _19459_;
 wire _19460_;
 wire _19461_;
 wire _19462_;
 wire _19463_;
 wire _19464_;
 wire _19465_;
 wire _19466_;
 wire _19467_;
 wire _19468_;
 wire _19469_;
 wire _19470_;
 wire _19471_;
 wire _19472_;
 wire _19473_;
 wire _19474_;
 wire _19475_;
 wire _19476_;
 wire _19477_;
 wire _19478_;
 wire _19479_;
 wire _19480_;
 wire _19481_;
 wire _19482_;
 wire _19483_;
 wire _19484_;
 wire _19485_;
 wire _19486_;
 wire _19487_;
 wire _19488_;
 wire _19489_;
 wire _19490_;
 wire _19491_;
 wire _19492_;
 wire _19493_;
 wire _19494_;
 wire _19495_;
 wire _19496_;
 wire _19497_;
 wire _19498_;
 wire _19499_;
 wire _19500_;
 wire _19501_;
 wire _19502_;
 wire _19503_;
 wire _19504_;
 wire _19505_;
 wire _19506_;
 wire _19507_;
 wire _19508_;
 wire _19509_;
 wire _19510_;
 wire _19511_;
 wire _19512_;
 wire _19513_;
 wire _19514_;
 wire _19515_;
 wire _19516_;
 wire _19517_;
 wire _19518_;
 wire _19519_;
 wire _19520_;
 wire _19521_;
 wire _19522_;
 wire _19523_;
 wire _19524_;
 wire _19525_;
 wire _19526_;
 wire _19527_;
 wire _19528_;
 wire _19529_;
 wire _19530_;
 wire _19531_;
 wire _19532_;
 wire _19533_;
 wire _19534_;
 wire _19535_;
 wire _19536_;
 wire _19537_;
 wire _19538_;
 wire _19539_;
 wire _19540_;
 wire _19541_;
 wire _19542_;
 wire _19543_;
 wire _19544_;
 wire _19545_;
 wire _19546_;
 wire _19547_;
 wire _19548_;
 wire _19549_;
 wire _19550_;
 wire _19551_;
 wire _19552_;
 wire _19553_;
 wire _19554_;
 wire _19555_;
 wire _19556_;
 wire _19557_;
 wire _19558_;
 wire _19559_;
 wire _19560_;
 wire _19561_;
 wire _19562_;
 wire _19563_;
 wire _19564_;
 wire _19565_;
 wire _19566_;
 wire _19567_;
 wire _19568_;
 wire _19569_;
 wire _19570_;
 wire _19571_;
 wire _19572_;
 wire _19573_;
 wire _19574_;
 wire _19575_;
 wire _19576_;
 wire _19577_;
 wire _19578_;
 wire _19579_;
 wire _19580_;
 wire _19581_;
 wire _19582_;
 wire _19583_;
 wire _19584_;
 wire _19585_;
 wire _19586_;
 wire _19587_;
 wire _19588_;
 wire _19589_;
 wire _19590_;
 wire _19591_;
 wire _19592_;
 wire _19593_;
 wire _19594_;
 wire _19595_;
 wire _19596_;
 wire _19597_;
 wire _19598_;
 wire _19599_;
 wire _19600_;
 wire _19601_;
 wire _19602_;
 wire _19603_;
 wire _19604_;
 wire _19605_;
 wire _19606_;
 wire _19607_;
 wire _19608_;
 wire _19609_;
 wire _19610_;
 wire _19611_;
 wire _19612_;
 wire _19613_;
 wire _19614_;
 wire _19615_;
 wire _19616_;
 wire _19617_;
 wire _19618_;
 wire _19619_;
 wire _19620_;
 wire _19621_;
 wire _19622_;
 wire _19623_;
 wire _19624_;
 wire _19625_;
 wire _19626_;
 wire _19627_;
 wire _19628_;
 wire _19629_;
 wire _19630_;
 wire _19631_;
 wire _19632_;
 wire _19633_;
 wire _19634_;
 wire _19635_;
 wire _19636_;
 wire _19637_;
 wire _19638_;
 wire _19639_;
 wire _19640_;
 wire _19641_;
 wire _19642_;
 wire _19643_;
 wire _19644_;
 wire _19645_;
 wire _19646_;
 wire _19647_;
 wire _19648_;
 wire _19649_;
 wire _19650_;
 wire _19651_;
 wire _19652_;
 wire _19653_;
 wire _19654_;
 wire _19655_;
 wire _19656_;
 wire _19657_;
 wire _19658_;
 wire _19659_;
 wire _19660_;
 wire _19661_;
 wire _19662_;
 wire _19663_;
 wire _19664_;
 wire _19665_;
 wire _19666_;
 wire _19667_;
 wire _19668_;
 wire _19669_;
 wire _19670_;
 wire _19671_;
 wire _19672_;
 wire _19673_;
 wire _19674_;
 wire _19675_;
 wire _19676_;
 wire _19677_;
 wire _19678_;
 wire _19679_;
 wire _19680_;
 wire _19681_;
 wire _19682_;
 wire _19683_;
 wire _19684_;
 wire _19685_;
 wire _19686_;
 wire _19687_;
 wire _19688_;
 wire _19689_;
 wire _19690_;
 wire _19691_;
 wire _19692_;
 wire _19693_;
 wire _19694_;
 wire _19695_;
 wire _19696_;
 wire _19697_;
 wire _19698_;
 wire _19699_;
 wire _19700_;
 wire _19701_;
 wire _19702_;
 wire _19703_;
 wire _19704_;
 wire _19705_;
 wire _19706_;
 wire _19707_;
 wire _19708_;
 wire _19709_;
 wire _19710_;
 wire _19711_;
 wire _19712_;
 wire _19713_;
 wire _19714_;
 wire _19715_;
 wire _19716_;
 wire _19717_;
 wire _19718_;
 wire _19719_;
 wire _19720_;
 wire _19721_;
 wire _19722_;
 wire _19723_;
 wire _19724_;
 wire _19725_;
 wire _19726_;
 wire _19727_;
 wire _19728_;
 wire _19729_;
 wire _19730_;
 wire _19731_;
 wire _19732_;
 wire _19733_;
 wire _19734_;
 wire _19735_;
 wire _19736_;
 wire _19737_;
 wire _19738_;
 wire _19739_;
 wire _19740_;
 wire _19741_;
 wire _19742_;
 wire _19743_;
 wire _19744_;
 wire _19745_;
 wire _19746_;
 wire _19747_;
 wire _19748_;
 wire _19749_;
 wire _19750_;
 wire _19751_;
 wire _19752_;
 wire _19753_;
 wire _19754_;
 wire _19755_;
 wire _19756_;
 wire _19757_;
 wire _19758_;
 wire _19759_;
 wire _19760_;
 wire _19761_;
 wire _19762_;
 wire _19763_;
 wire _19764_;
 wire _19765_;
 wire _19766_;
 wire _19767_;
 wire _19768_;
 wire _19769_;
 wire _19770_;
 wire _19771_;
 wire _19772_;
 wire _19773_;
 wire _19774_;
 wire _19775_;
 wire _19776_;
 wire _19777_;
 wire _19778_;
 wire _19779_;
 wire _19780_;
 wire _19781_;
 wire _19782_;
 wire _19783_;
 wire _19784_;
 wire _19785_;
 wire _19786_;
 wire _19787_;
 wire _19788_;
 wire _19789_;
 wire _19790_;
 wire _19791_;
 wire _19792_;
 wire _19793_;
 wire _19794_;
 wire _19795_;
 wire _19796_;
 wire _19797_;
 wire _19798_;
 wire _19799_;
 wire _19800_;
 wire _19801_;
 wire _19802_;
 wire _19803_;
 wire _19804_;
 wire _19805_;
 wire _19806_;
 wire _19807_;
 wire _19808_;
 wire _19809_;
 wire _19810_;
 wire _19811_;
 wire _19812_;
 wire _19813_;
 wire _19814_;
 wire _19815_;
 wire _19816_;
 wire _19817_;
 wire _19818_;
 wire _19819_;
 wire _19820_;
 wire _19821_;
 wire _19822_;
 wire _19823_;
 wire _19824_;
 wire _19825_;
 wire _19826_;
 wire _19827_;
 wire _19828_;
 wire _19829_;
 wire _19830_;
 wire _19831_;
 wire _19832_;
 wire _19833_;
 wire _19834_;
 wire _19835_;
 wire _19836_;
 wire _19837_;
 wire _19838_;
 wire _19839_;
 wire _19840_;
 wire _19841_;
 wire _19842_;
 wire _19843_;
 wire _19844_;
 wire _19845_;
 wire _19846_;
 wire _19847_;
 wire _19848_;
 wire _19849_;
 wire _19850_;
 wire _19851_;
 wire _19852_;
 wire _19853_;
 wire _19854_;
 wire _19855_;
 wire _19856_;
 wire _19857_;
 wire _19858_;
 wire _19859_;
 wire _19860_;
 wire _19861_;
 wire _19862_;
 wire _19863_;
 wire _19864_;
 wire _19865_;
 wire _19866_;
 wire \alu_add_sub[0] ;
 wire \alu_add_sub[10] ;
 wire \alu_add_sub[11] ;
 wire \alu_add_sub[12] ;
 wire \alu_add_sub[13] ;
 wire \alu_add_sub[14] ;
 wire \alu_add_sub[15] ;
 wire \alu_add_sub[16] ;
 wire \alu_add_sub[17] ;
 wire \alu_add_sub[18] ;
 wire \alu_add_sub[19] ;
 wire \alu_add_sub[1] ;
 wire \alu_add_sub[20] ;
 wire \alu_add_sub[21] ;
 wire \alu_add_sub[22] ;
 wire \alu_add_sub[23] ;
 wire \alu_add_sub[24] ;
 wire \alu_add_sub[25] ;
 wire \alu_add_sub[26] ;
 wire \alu_add_sub[27] ;
 wire \alu_add_sub[28] ;
 wire \alu_add_sub[29] ;
 wire \alu_add_sub[2] ;
 wire \alu_add_sub[30] ;
 wire \alu_add_sub[31] ;
 wire \alu_add_sub[3] ;
 wire \alu_add_sub[4] ;
 wire \alu_add_sub[5] ;
 wire \alu_add_sub[6] ;
 wire \alu_add_sub[7] ;
 wire \alu_add_sub[8] ;
 wire \alu_add_sub[9] ;
 wire alu_eq;
 wire alu_lts;
 wire alu_ltu;
 wire \alu_out[0] ;
 wire \alu_out[10] ;
 wire \alu_out[11] ;
 wire \alu_out[12] ;
 wire \alu_out[13] ;
 wire \alu_out[14] ;
 wire \alu_out[15] ;
 wire \alu_out[16] ;
 wire \alu_out[17] ;
 wire \alu_out[18] ;
 wire \alu_out[19] ;
 wire \alu_out[1] ;
 wire \alu_out[20] ;
 wire \alu_out[21] ;
 wire \alu_out[22] ;
 wire \alu_out[23] ;
 wire \alu_out[24] ;
 wire \alu_out[25] ;
 wire \alu_out[26] ;
 wire \alu_out[27] ;
 wire \alu_out[28] ;
 wire \alu_out[29] ;
 wire \alu_out[2] ;
 wire \alu_out[30] ;
 wire \alu_out[31] ;
 wire \alu_out[3] ;
 wire \alu_out[4] ;
 wire \alu_out[5] ;
 wire \alu_out[6] ;
 wire \alu_out[7] ;
 wire \alu_out[8] ;
 wire \alu_out[9] ;
 wire \alu_out_q[0] ;
 wire \alu_out_q[10] ;
 wire \alu_out_q[11] ;
 wire \alu_out_q[12] ;
 wire \alu_out_q[13] ;
 wire \alu_out_q[14] ;
 wire \alu_out_q[15] ;
 wire \alu_out_q[16] ;
 wire \alu_out_q[17] ;
 wire \alu_out_q[18] ;
 wire \alu_out_q[19] ;
 wire \alu_out_q[1] ;
 wire \alu_out_q[20] ;
 wire \alu_out_q[21] ;
 wire \alu_out_q[22] ;
 wire \alu_out_q[23] ;
 wire \alu_out_q[24] ;
 wire \alu_out_q[25] ;
 wire \alu_out_q[26] ;
 wire \alu_out_q[27] ;
 wire \alu_out_q[28] ;
 wire \alu_out_q[29] ;
 wire \alu_out_q[2] ;
 wire \alu_out_q[30] ;
 wire \alu_out_q[31] ;
 wire \alu_out_q[3] ;
 wire \alu_out_q[4] ;
 wire \alu_out_q[5] ;
 wire \alu_out_q[6] ;
 wire \alu_out_q[7] ;
 wire \alu_out_q[8] ;
 wire \alu_out_q[9] ;
 wire \alu_shl[0] ;
 wire \alu_shl[10] ;
 wire \alu_shl[11] ;
 wire \alu_shl[12] ;
 wire \alu_shl[13] ;
 wire \alu_shl[14] ;
 wire \alu_shl[15] ;
 wire \alu_shl[16] ;
 wire \alu_shl[17] ;
 wire \alu_shl[18] ;
 wire \alu_shl[19] ;
 wire \alu_shl[1] ;
 wire \alu_shl[20] ;
 wire \alu_shl[21] ;
 wire \alu_shl[22] ;
 wire \alu_shl[23] ;
 wire \alu_shl[24] ;
 wire \alu_shl[25] ;
 wire \alu_shl[26] ;
 wire \alu_shl[27] ;
 wire \alu_shl[28] ;
 wire \alu_shl[29] ;
 wire \alu_shl[2] ;
 wire \alu_shl[30] ;
 wire \alu_shl[31] ;
 wire \alu_shl[3] ;
 wire \alu_shl[4] ;
 wire \alu_shl[5] ;
 wire \alu_shl[6] ;
 wire \alu_shl[7] ;
 wire \alu_shl[8] ;
 wire \alu_shl[9] ;
 wire \alu_shr[0] ;
 wire \alu_shr[10] ;
 wire \alu_shr[11] ;
 wire \alu_shr[12] ;
 wire \alu_shr[13] ;
 wire \alu_shr[14] ;
 wire \alu_shr[15] ;
 wire \alu_shr[16] ;
 wire \alu_shr[17] ;
 wire \alu_shr[18] ;
 wire \alu_shr[19] ;
 wire \alu_shr[1] ;
 wire \alu_shr[20] ;
 wire \alu_shr[21] ;
 wire \alu_shr[22] ;
 wire \alu_shr[23] ;
 wire \alu_shr[24] ;
 wire \alu_shr[25] ;
 wire \alu_shr[26] ;
 wire \alu_shr[27] ;
 wire \alu_shr[28] ;
 wire \alu_shr[29] ;
 wire \alu_shr[2] ;
 wire \alu_shr[30] ;
 wire \alu_shr[31] ;
 wire \alu_shr[3] ;
 wire \alu_shr[4] ;
 wire \alu_shr[5] ;
 wire \alu_shr[6] ;
 wire \alu_shr[7] ;
 wire \alu_shr[8] ;
 wire \alu_shr[9] ;
 wire alu_wait;
 wire \count_cycle[0] ;
 wire \count_cycle[10] ;
 wire \count_cycle[11] ;
 wire \count_cycle[12] ;
 wire \count_cycle[13] ;
 wire \count_cycle[14] ;
 wire \count_cycle[15] ;
 wire \count_cycle[16] ;
 wire \count_cycle[17] ;
 wire \count_cycle[18] ;
 wire \count_cycle[19] ;
 wire \count_cycle[1] ;
 wire \count_cycle[20] ;
 wire \count_cycle[21] ;
 wire \count_cycle[22] ;
 wire \count_cycle[23] ;
 wire \count_cycle[24] ;
 wire \count_cycle[25] ;
 wire \count_cycle[26] ;
 wire \count_cycle[27] ;
 wire \count_cycle[28] ;
 wire \count_cycle[29] ;
 wire \count_cycle[2] ;
 wire \count_cycle[30] ;
 wire \count_cycle[31] ;
 wire \count_cycle[32] ;
 wire \count_cycle[33] ;
 wire \count_cycle[34] ;
 wire \count_cycle[35] ;
 wire \count_cycle[36] ;
 wire \count_cycle[37] ;
 wire \count_cycle[38] ;
 wire \count_cycle[39] ;
 wire \count_cycle[3] ;
 wire \count_cycle[40] ;
 wire \count_cycle[41] ;
 wire \count_cycle[42] ;
 wire \count_cycle[43] ;
 wire \count_cycle[44] ;
 wire \count_cycle[45] ;
 wire \count_cycle[46] ;
 wire \count_cycle[47] ;
 wire \count_cycle[48] ;
 wire \count_cycle[49] ;
 wire \count_cycle[4] ;
 wire \count_cycle[50] ;
 wire \count_cycle[51] ;
 wire \count_cycle[52] ;
 wire \count_cycle[53] ;
 wire \count_cycle[54] ;
 wire \count_cycle[55] ;
 wire \count_cycle[56] ;
 wire \count_cycle[57] ;
 wire \count_cycle[58] ;
 wire \count_cycle[59] ;
 wire \count_cycle[5] ;
 wire \count_cycle[60] ;
 wire \count_cycle[61] ;
 wire \count_cycle[62] ;
 wire \count_cycle[63] ;
 wire \count_cycle[6] ;
 wire \count_cycle[7] ;
 wire \count_cycle[8] ;
 wire \count_cycle[9] ;
 wire \count_instr[0] ;
 wire \count_instr[10] ;
 wire \count_instr[11] ;
 wire \count_instr[12] ;
 wire \count_instr[13] ;
 wire \count_instr[14] ;
 wire \count_instr[15] ;
 wire \count_instr[16] ;
 wire \count_instr[17] ;
 wire \count_instr[18] ;
 wire \count_instr[19] ;
 wire \count_instr[1] ;
 wire \count_instr[20] ;
 wire \count_instr[21] ;
 wire \count_instr[22] ;
 wire \count_instr[23] ;
 wire \count_instr[24] ;
 wire \count_instr[25] ;
 wire \count_instr[26] ;
 wire \count_instr[27] ;
 wire \count_instr[28] ;
 wire \count_instr[29] ;
 wire \count_instr[2] ;
 wire \count_instr[30] ;
 wire \count_instr[31] ;
 wire \count_instr[32] ;
 wire \count_instr[33] ;
 wire \count_instr[34] ;
 wire \count_instr[35] ;
 wire \count_instr[36] ;
 wire \count_instr[37] ;
 wire \count_instr[38] ;
 wire \count_instr[39] ;
 wire \count_instr[3] ;
 wire \count_instr[40] ;
 wire \count_instr[41] ;
 wire \count_instr[42] ;
 wire \count_instr[43] ;
 wire \count_instr[44] ;
 wire \count_instr[45] ;
 wire \count_instr[46] ;
 wire \count_instr[47] ;
 wire \count_instr[48] ;
 wire \count_instr[49] ;
 wire \count_instr[4] ;
 wire \count_instr[50] ;
 wire \count_instr[51] ;
 wire \count_instr[52] ;
 wire \count_instr[53] ;
 wire \count_instr[54] ;
 wire \count_instr[55] ;
 wire \count_instr[56] ;
 wire \count_instr[57] ;
 wire \count_instr[58] ;
 wire \count_instr[59] ;
 wire \count_instr[5] ;
 wire \count_instr[60] ;
 wire \count_instr[61] ;
 wire \count_instr[62] ;
 wire \count_instr[63] ;
 wire \count_instr[6] ;
 wire \count_instr[7] ;
 wire \count_instr[8] ;
 wire \count_instr[9] ;
 wire \cpu_state[0] ;
 wire \cpu_state[1] ;
 wire \cpu_state[2] ;
 wire \cpu_state[3] ;
 wire \cpu_state[4] ;
 wire \cpu_state[5] ;
 wire \cpu_state[6] ;
 wire \cpuregs[0][0] ;
 wire \cpuregs[0][10] ;
 wire \cpuregs[0][11] ;
 wire \cpuregs[0][12] ;
 wire \cpuregs[0][13] ;
 wire \cpuregs[0][14] ;
 wire \cpuregs[0][15] ;
 wire \cpuregs[0][16] ;
 wire \cpuregs[0][17] ;
 wire \cpuregs[0][18] ;
 wire \cpuregs[0][19] ;
 wire \cpuregs[0][1] ;
 wire \cpuregs[0][20] ;
 wire \cpuregs[0][21] ;
 wire \cpuregs[0][22] ;
 wire \cpuregs[0][23] ;
 wire \cpuregs[0][24] ;
 wire \cpuregs[0][25] ;
 wire \cpuregs[0][26] ;
 wire \cpuregs[0][27] ;
 wire \cpuregs[0][28] ;
 wire \cpuregs[0][29] ;
 wire \cpuregs[0][2] ;
 wire \cpuregs[0][30] ;
 wire \cpuregs[0][31] ;
 wire \cpuregs[0][3] ;
 wire \cpuregs[0][4] ;
 wire \cpuregs[0][5] ;
 wire \cpuregs[0][6] ;
 wire \cpuregs[0][7] ;
 wire \cpuregs[0][8] ;
 wire \cpuregs[0][9] ;
 wire \cpuregs[10][0] ;
 wire \cpuregs[10][10] ;
 wire \cpuregs[10][11] ;
 wire \cpuregs[10][12] ;
 wire \cpuregs[10][13] ;
 wire \cpuregs[10][14] ;
 wire \cpuregs[10][15] ;
 wire \cpuregs[10][16] ;
 wire \cpuregs[10][17] ;
 wire \cpuregs[10][18] ;
 wire \cpuregs[10][19] ;
 wire \cpuregs[10][1] ;
 wire \cpuregs[10][20] ;
 wire \cpuregs[10][21] ;
 wire \cpuregs[10][22] ;
 wire \cpuregs[10][23] ;
 wire \cpuregs[10][24] ;
 wire \cpuregs[10][25] ;
 wire \cpuregs[10][26] ;
 wire \cpuregs[10][27] ;
 wire \cpuregs[10][28] ;
 wire \cpuregs[10][29] ;
 wire \cpuregs[10][2] ;
 wire \cpuregs[10][30] ;
 wire \cpuregs[10][31] ;
 wire \cpuregs[10][3] ;
 wire \cpuregs[10][4] ;
 wire \cpuregs[10][5] ;
 wire \cpuregs[10][6] ;
 wire \cpuregs[10][7] ;
 wire \cpuregs[10][8] ;
 wire \cpuregs[10][9] ;
 wire \cpuregs[11][0] ;
 wire \cpuregs[11][10] ;
 wire \cpuregs[11][11] ;
 wire \cpuregs[11][12] ;
 wire \cpuregs[11][13] ;
 wire \cpuregs[11][14] ;
 wire \cpuregs[11][15] ;
 wire \cpuregs[11][16] ;
 wire \cpuregs[11][17] ;
 wire \cpuregs[11][18] ;
 wire \cpuregs[11][19] ;
 wire \cpuregs[11][1] ;
 wire \cpuregs[11][20] ;
 wire \cpuregs[11][21] ;
 wire \cpuregs[11][22] ;
 wire \cpuregs[11][23] ;
 wire \cpuregs[11][24] ;
 wire \cpuregs[11][25] ;
 wire \cpuregs[11][26] ;
 wire \cpuregs[11][27] ;
 wire \cpuregs[11][28] ;
 wire \cpuregs[11][29] ;
 wire \cpuregs[11][2] ;
 wire \cpuregs[11][30] ;
 wire \cpuregs[11][31] ;
 wire \cpuregs[11][3] ;
 wire \cpuregs[11][4] ;
 wire \cpuregs[11][5] ;
 wire \cpuregs[11][6] ;
 wire \cpuregs[11][7] ;
 wire \cpuregs[11][8] ;
 wire \cpuregs[11][9] ;
 wire \cpuregs[12][0] ;
 wire \cpuregs[12][10] ;
 wire \cpuregs[12][11] ;
 wire \cpuregs[12][12] ;
 wire \cpuregs[12][13] ;
 wire \cpuregs[12][14] ;
 wire \cpuregs[12][15] ;
 wire \cpuregs[12][16] ;
 wire \cpuregs[12][17] ;
 wire \cpuregs[12][18] ;
 wire \cpuregs[12][19] ;
 wire \cpuregs[12][1] ;
 wire \cpuregs[12][20] ;
 wire \cpuregs[12][21] ;
 wire \cpuregs[12][22] ;
 wire \cpuregs[12][23] ;
 wire \cpuregs[12][24] ;
 wire \cpuregs[12][25] ;
 wire \cpuregs[12][26] ;
 wire \cpuregs[12][27] ;
 wire \cpuregs[12][28] ;
 wire \cpuregs[12][29] ;
 wire \cpuregs[12][2] ;
 wire \cpuregs[12][30] ;
 wire \cpuregs[12][31] ;
 wire \cpuregs[12][3] ;
 wire \cpuregs[12][4] ;
 wire \cpuregs[12][5] ;
 wire \cpuregs[12][6] ;
 wire \cpuregs[12][7] ;
 wire \cpuregs[12][8] ;
 wire \cpuregs[12][9] ;
 wire \cpuregs[13][0] ;
 wire \cpuregs[13][10] ;
 wire \cpuregs[13][11] ;
 wire \cpuregs[13][12] ;
 wire \cpuregs[13][13] ;
 wire \cpuregs[13][14] ;
 wire \cpuregs[13][15] ;
 wire \cpuregs[13][16] ;
 wire \cpuregs[13][17] ;
 wire \cpuregs[13][18] ;
 wire \cpuregs[13][19] ;
 wire \cpuregs[13][1] ;
 wire \cpuregs[13][20] ;
 wire \cpuregs[13][21] ;
 wire \cpuregs[13][22] ;
 wire \cpuregs[13][23] ;
 wire \cpuregs[13][24] ;
 wire \cpuregs[13][25] ;
 wire \cpuregs[13][26] ;
 wire \cpuregs[13][27] ;
 wire \cpuregs[13][28] ;
 wire \cpuregs[13][29] ;
 wire \cpuregs[13][2] ;
 wire \cpuregs[13][30] ;
 wire \cpuregs[13][31] ;
 wire \cpuregs[13][3] ;
 wire \cpuregs[13][4] ;
 wire \cpuregs[13][5] ;
 wire \cpuregs[13][6] ;
 wire \cpuregs[13][7] ;
 wire \cpuregs[13][8] ;
 wire \cpuregs[13][9] ;
 wire \cpuregs[14][0] ;
 wire \cpuregs[14][10] ;
 wire \cpuregs[14][11] ;
 wire \cpuregs[14][12] ;
 wire \cpuregs[14][13] ;
 wire \cpuregs[14][14] ;
 wire \cpuregs[14][15] ;
 wire \cpuregs[14][16] ;
 wire \cpuregs[14][17] ;
 wire \cpuregs[14][18] ;
 wire \cpuregs[14][19] ;
 wire \cpuregs[14][1] ;
 wire \cpuregs[14][20] ;
 wire \cpuregs[14][21] ;
 wire \cpuregs[14][22] ;
 wire \cpuregs[14][23] ;
 wire \cpuregs[14][24] ;
 wire \cpuregs[14][25] ;
 wire \cpuregs[14][26] ;
 wire \cpuregs[14][27] ;
 wire \cpuregs[14][28] ;
 wire \cpuregs[14][29] ;
 wire \cpuregs[14][2] ;
 wire \cpuregs[14][30] ;
 wire \cpuregs[14][31] ;
 wire \cpuregs[14][3] ;
 wire \cpuregs[14][4] ;
 wire \cpuregs[14][5] ;
 wire \cpuregs[14][6] ;
 wire \cpuregs[14][7] ;
 wire \cpuregs[14][8] ;
 wire \cpuregs[14][9] ;
 wire \cpuregs[15][0] ;
 wire \cpuregs[15][10] ;
 wire \cpuregs[15][11] ;
 wire \cpuregs[15][12] ;
 wire \cpuregs[15][13] ;
 wire \cpuregs[15][14] ;
 wire \cpuregs[15][15] ;
 wire \cpuregs[15][16] ;
 wire \cpuregs[15][17] ;
 wire \cpuregs[15][18] ;
 wire \cpuregs[15][19] ;
 wire \cpuregs[15][1] ;
 wire \cpuregs[15][20] ;
 wire \cpuregs[15][21] ;
 wire \cpuregs[15][22] ;
 wire \cpuregs[15][23] ;
 wire \cpuregs[15][24] ;
 wire \cpuregs[15][25] ;
 wire \cpuregs[15][26] ;
 wire \cpuregs[15][27] ;
 wire \cpuregs[15][28] ;
 wire \cpuregs[15][29] ;
 wire \cpuregs[15][2] ;
 wire \cpuregs[15][30] ;
 wire \cpuregs[15][31] ;
 wire \cpuregs[15][3] ;
 wire \cpuregs[15][4] ;
 wire \cpuregs[15][5] ;
 wire \cpuregs[15][6] ;
 wire \cpuregs[15][7] ;
 wire \cpuregs[15][8] ;
 wire \cpuregs[15][9] ;
 wire \cpuregs[16][0] ;
 wire \cpuregs[16][10] ;
 wire \cpuregs[16][11] ;
 wire \cpuregs[16][12] ;
 wire \cpuregs[16][13] ;
 wire \cpuregs[16][14] ;
 wire \cpuregs[16][15] ;
 wire \cpuregs[16][16] ;
 wire \cpuregs[16][17] ;
 wire \cpuregs[16][18] ;
 wire \cpuregs[16][19] ;
 wire \cpuregs[16][1] ;
 wire \cpuregs[16][20] ;
 wire \cpuregs[16][21] ;
 wire \cpuregs[16][22] ;
 wire \cpuregs[16][23] ;
 wire \cpuregs[16][24] ;
 wire \cpuregs[16][25] ;
 wire \cpuregs[16][26] ;
 wire \cpuregs[16][27] ;
 wire \cpuregs[16][28] ;
 wire \cpuregs[16][29] ;
 wire \cpuregs[16][2] ;
 wire \cpuregs[16][30] ;
 wire \cpuregs[16][31] ;
 wire \cpuregs[16][3] ;
 wire \cpuregs[16][4] ;
 wire \cpuregs[16][5] ;
 wire \cpuregs[16][6] ;
 wire \cpuregs[16][7] ;
 wire \cpuregs[16][8] ;
 wire \cpuregs[16][9] ;
 wire \cpuregs[17][0] ;
 wire \cpuregs[17][10] ;
 wire \cpuregs[17][11] ;
 wire \cpuregs[17][12] ;
 wire \cpuregs[17][13] ;
 wire \cpuregs[17][14] ;
 wire \cpuregs[17][15] ;
 wire \cpuregs[17][16] ;
 wire \cpuregs[17][17] ;
 wire \cpuregs[17][18] ;
 wire \cpuregs[17][19] ;
 wire \cpuregs[17][1] ;
 wire \cpuregs[17][20] ;
 wire \cpuregs[17][21] ;
 wire \cpuregs[17][22] ;
 wire \cpuregs[17][23] ;
 wire \cpuregs[17][24] ;
 wire \cpuregs[17][25] ;
 wire \cpuregs[17][26] ;
 wire \cpuregs[17][27] ;
 wire \cpuregs[17][28] ;
 wire \cpuregs[17][29] ;
 wire \cpuregs[17][2] ;
 wire \cpuregs[17][30] ;
 wire \cpuregs[17][31] ;
 wire \cpuregs[17][3] ;
 wire \cpuregs[17][4] ;
 wire \cpuregs[17][5] ;
 wire \cpuregs[17][6] ;
 wire \cpuregs[17][7] ;
 wire \cpuregs[17][8] ;
 wire \cpuregs[17][9] ;
 wire \cpuregs[18][0] ;
 wire \cpuregs[18][10] ;
 wire \cpuregs[18][11] ;
 wire \cpuregs[18][12] ;
 wire \cpuregs[18][13] ;
 wire \cpuregs[18][14] ;
 wire \cpuregs[18][15] ;
 wire \cpuregs[18][16] ;
 wire \cpuregs[18][17] ;
 wire \cpuregs[18][18] ;
 wire \cpuregs[18][19] ;
 wire \cpuregs[18][1] ;
 wire \cpuregs[18][20] ;
 wire \cpuregs[18][21] ;
 wire \cpuregs[18][22] ;
 wire \cpuregs[18][23] ;
 wire \cpuregs[18][24] ;
 wire \cpuregs[18][25] ;
 wire \cpuregs[18][26] ;
 wire \cpuregs[18][27] ;
 wire \cpuregs[18][28] ;
 wire \cpuregs[18][29] ;
 wire \cpuregs[18][2] ;
 wire \cpuregs[18][30] ;
 wire \cpuregs[18][31] ;
 wire \cpuregs[18][3] ;
 wire \cpuregs[18][4] ;
 wire \cpuregs[18][5] ;
 wire \cpuregs[18][6] ;
 wire \cpuregs[18][7] ;
 wire \cpuregs[18][8] ;
 wire \cpuregs[18][9] ;
 wire \cpuregs[19][0] ;
 wire \cpuregs[19][10] ;
 wire \cpuregs[19][11] ;
 wire \cpuregs[19][12] ;
 wire \cpuregs[19][13] ;
 wire \cpuregs[19][14] ;
 wire \cpuregs[19][15] ;
 wire \cpuregs[19][16] ;
 wire \cpuregs[19][17] ;
 wire \cpuregs[19][18] ;
 wire \cpuregs[19][19] ;
 wire \cpuregs[19][1] ;
 wire \cpuregs[19][20] ;
 wire \cpuregs[19][21] ;
 wire \cpuregs[19][22] ;
 wire \cpuregs[19][23] ;
 wire \cpuregs[19][24] ;
 wire \cpuregs[19][25] ;
 wire \cpuregs[19][26] ;
 wire \cpuregs[19][27] ;
 wire \cpuregs[19][28] ;
 wire \cpuregs[19][29] ;
 wire \cpuregs[19][2] ;
 wire \cpuregs[19][30] ;
 wire \cpuregs[19][31] ;
 wire \cpuregs[19][3] ;
 wire \cpuregs[19][4] ;
 wire \cpuregs[19][5] ;
 wire \cpuregs[19][6] ;
 wire \cpuregs[19][7] ;
 wire \cpuregs[19][8] ;
 wire \cpuregs[19][9] ;
 wire \cpuregs[1][0] ;
 wire \cpuregs[1][10] ;
 wire \cpuregs[1][11] ;
 wire \cpuregs[1][12] ;
 wire \cpuregs[1][13] ;
 wire \cpuregs[1][14] ;
 wire \cpuregs[1][15] ;
 wire \cpuregs[1][16] ;
 wire \cpuregs[1][17] ;
 wire \cpuregs[1][18] ;
 wire \cpuregs[1][19] ;
 wire \cpuregs[1][1] ;
 wire \cpuregs[1][20] ;
 wire \cpuregs[1][21] ;
 wire \cpuregs[1][22] ;
 wire \cpuregs[1][23] ;
 wire \cpuregs[1][24] ;
 wire \cpuregs[1][25] ;
 wire \cpuregs[1][26] ;
 wire \cpuregs[1][27] ;
 wire \cpuregs[1][28] ;
 wire \cpuregs[1][29] ;
 wire \cpuregs[1][2] ;
 wire \cpuregs[1][30] ;
 wire \cpuregs[1][31] ;
 wire \cpuregs[1][3] ;
 wire \cpuregs[1][4] ;
 wire \cpuregs[1][5] ;
 wire \cpuregs[1][6] ;
 wire \cpuregs[1][7] ;
 wire \cpuregs[1][8] ;
 wire \cpuregs[1][9] ;
 wire \cpuregs[2][0] ;
 wire \cpuregs[2][10] ;
 wire \cpuregs[2][11] ;
 wire \cpuregs[2][12] ;
 wire \cpuregs[2][13] ;
 wire \cpuregs[2][14] ;
 wire \cpuregs[2][15] ;
 wire \cpuregs[2][16] ;
 wire \cpuregs[2][17] ;
 wire \cpuregs[2][18] ;
 wire \cpuregs[2][19] ;
 wire \cpuregs[2][1] ;
 wire \cpuregs[2][20] ;
 wire \cpuregs[2][21] ;
 wire \cpuregs[2][22] ;
 wire \cpuregs[2][23] ;
 wire \cpuregs[2][24] ;
 wire \cpuregs[2][25] ;
 wire \cpuregs[2][26] ;
 wire \cpuregs[2][27] ;
 wire \cpuregs[2][28] ;
 wire \cpuregs[2][29] ;
 wire \cpuregs[2][2] ;
 wire \cpuregs[2][30] ;
 wire \cpuregs[2][31] ;
 wire \cpuregs[2][3] ;
 wire \cpuregs[2][4] ;
 wire \cpuregs[2][5] ;
 wire \cpuregs[2][6] ;
 wire \cpuregs[2][7] ;
 wire \cpuregs[2][8] ;
 wire \cpuregs[2][9] ;
 wire \cpuregs[3][0] ;
 wire \cpuregs[3][10] ;
 wire \cpuregs[3][11] ;
 wire \cpuregs[3][12] ;
 wire \cpuregs[3][13] ;
 wire \cpuregs[3][14] ;
 wire \cpuregs[3][15] ;
 wire \cpuregs[3][16] ;
 wire \cpuregs[3][17] ;
 wire \cpuregs[3][18] ;
 wire \cpuregs[3][19] ;
 wire \cpuregs[3][1] ;
 wire \cpuregs[3][20] ;
 wire \cpuregs[3][21] ;
 wire \cpuregs[3][22] ;
 wire \cpuregs[3][23] ;
 wire \cpuregs[3][24] ;
 wire \cpuregs[3][25] ;
 wire \cpuregs[3][26] ;
 wire \cpuregs[3][27] ;
 wire \cpuregs[3][28] ;
 wire \cpuregs[3][29] ;
 wire \cpuregs[3][2] ;
 wire \cpuregs[3][30] ;
 wire \cpuregs[3][31] ;
 wire \cpuregs[3][3] ;
 wire \cpuregs[3][4] ;
 wire \cpuregs[3][5] ;
 wire \cpuregs[3][6] ;
 wire \cpuregs[3][7] ;
 wire \cpuregs[3][8] ;
 wire \cpuregs[3][9] ;
 wire \cpuregs[4][0] ;
 wire \cpuregs[4][10] ;
 wire \cpuregs[4][11] ;
 wire \cpuregs[4][12] ;
 wire \cpuregs[4][13] ;
 wire \cpuregs[4][14] ;
 wire \cpuregs[4][15] ;
 wire \cpuregs[4][16] ;
 wire \cpuregs[4][17] ;
 wire \cpuregs[4][18] ;
 wire \cpuregs[4][19] ;
 wire \cpuregs[4][1] ;
 wire \cpuregs[4][20] ;
 wire \cpuregs[4][21] ;
 wire \cpuregs[4][22] ;
 wire \cpuregs[4][23] ;
 wire \cpuregs[4][24] ;
 wire \cpuregs[4][25] ;
 wire \cpuregs[4][26] ;
 wire \cpuregs[4][27] ;
 wire \cpuregs[4][28] ;
 wire \cpuregs[4][29] ;
 wire \cpuregs[4][2] ;
 wire \cpuregs[4][30] ;
 wire \cpuregs[4][31] ;
 wire \cpuregs[4][3] ;
 wire \cpuregs[4][4] ;
 wire \cpuregs[4][5] ;
 wire \cpuregs[4][6] ;
 wire \cpuregs[4][7] ;
 wire \cpuregs[4][8] ;
 wire \cpuregs[4][9] ;
 wire \cpuregs[5][0] ;
 wire \cpuregs[5][10] ;
 wire \cpuregs[5][11] ;
 wire \cpuregs[5][12] ;
 wire \cpuregs[5][13] ;
 wire \cpuregs[5][14] ;
 wire \cpuregs[5][15] ;
 wire \cpuregs[5][16] ;
 wire \cpuregs[5][17] ;
 wire \cpuregs[5][18] ;
 wire \cpuregs[5][19] ;
 wire \cpuregs[5][1] ;
 wire \cpuregs[5][20] ;
 wire \cpuregs[5][21] ;
 wire \cpuregs[5][22] ;
 wire \cpuregs[5][23] ;
 wire \cpuregs[5][24] ;
 wire \cpuregs[5][25] ;
 wire \cpuregs[5][26] ;
 wire \cpuregs[5][27] ;
 wire \cpuregs[5][28] ;
 wire \cpuregs[5][29] ;
 wire \cpuregs[5][2] ;
 wire \cpuregs[5][30] ;
 wire \cpuregs[5][31] ;
 wire \cpuregs[5][3] ;
 wire \cpuregs[5][4] ;
 wire \cpuregs[5][5] ;
 wire \cpuregs[5][6] ;
 wire \cpuregs[5][7] ;
 wire \cpuregs[5][8] ;
 wire \cpuregs[5][9] ;
 wire \cpuregs[6][0] ;
 wire \cpuregs[6][10] ;
 wire \cpuregs[6][11] ;
 wire \cpuregs[6][12] ;
 wire \cpuregs[6][13] ;
 wire \cpuregs[6][14] ;
 wire \cpuregs[6][15] ;
 wire \cpuregs[6][16] ;
 wire \cpuregs[6][17] ;
 wire \cpuregs[6][18] ;
 wire \cpuregs[6][19] ;
 wire \cpuregs[6][1] ;
 wire \cpuregs[6][20] ;
 wire \cpuregs[6][21] ;
 wire \cpuregs[6][22] ;
 wire \cpuregs[6][23] ;
 wire \cpuregs[6][24] ;
 wire \cpuregs[6][25] ;
 wire \cpuregs[6][26] ;
 wire \cpuregs[6][27] ;
 wire \cpuregs[6][28] ;
 wire \cpuregs[6][29] ;
 wire \cpuregs[6][2] ;
 wire \cpuregs[6][30] ;
 wire \cpuregs[6][31] ;
 wire \cpuregs[6][3] ;
 wire \cpuregs[6][4] ;
 wire \cpuregs[6][5] ;
 wire \cpuregs[6][6] ;
 wire \cpuregs[6][7] ;
 wire \cpuregs[6][8] ;
 wire \cpuregs[6][9] ;
 wire \cpuregs[7][0] ;
 wire \cpuregs[7][10] ;
 wire \cpuregs[7][11] ;
 wire \cpuregs[7][12] ;
 wire \cpuregs[7][13] ;
 wire \cpuregs[7][14] ;
 wire \cpuregs[7][15] ;
 wire \cpuregs[7][16] ;
 wire \cpuregs[7][17] ;
 wire \cpuregs[7][18] ;
 wire \cpuregs[7][19] ;
 wire \cpuregs[7][1] ;
 wire \cpuregs[7][20] ;
 wire \cpuregs[7][21] ;
 wire \cpuregs[7][22] ;
 wire \cpuregs[7][23] ;
 wire \cpuregs[7][24] ;
 wire \cpuregs[7][25] ;
 wire \cpuregs[7][26] ;
 wire \cpuregs[7][27] ;
 wire \cpuregs[7][28] ;
 wire \cpuregs[7][29] ;
 wire \cpuregs[7][2] ;
 wire \cpuregs[7][30] ;
 wire \cpuregs[7][31] ;
 wire \cpuregs[7][3] ;
 wire \cpuregs[7][4] ;
 wire \cpuregs[7][5] ;
 wire \cpuregs[7][6] ;
 wire \cpuregs[7][7] ;
 wire \cpuregs[7][8] ;
 wire \cpuregs[7][9] ;
 wire \cpuregs[8][0] ;
 wire \cpuregs[8][10] ;
 wire \cpuregs[8][11] ;
 wire \cpuregs[8][12] ;
 wire \cpuregs[8][13] ;
 wire \cpuregs[8][14] ;
 wire \cpuregs[8][15] ;
 wire \cpuregs[8][16] ;
 wire \cpuregs[8][17] ;
 wire \cpuregs[8][18] ;
 wire \cpuregs[8][19] ;
 wire \cpuregs[8][1] ;
 wire \cpuregs[8][20] ;
 wire \cpuregs[8][21] ;
 wire \cpuregs[8][22] ;
 wire \cpuregs[8][23] ;
 wire \cpuregs[8][24] ;
 wire \cpuregs[8][25] ;
 wire \cpuregs[8][26] ;
 wire \cpuregs[8][27] ;
 wire \cpuregs[8][28] ;
 wire \cpuregs[8][29] ;
 wire \cpuregs[8][2] ;
 wire \cpuregs[8][30] ;
 wire \cpuregs[8][31] ;
 wire \cpuregs[8][3] ;
 wire \cpuregs[8][4] ;
 wire \cpuregs[8][5] ;
 wire \cpuregs[8][6] ;
 wire \cpuregs[8][7] ;
 wire \cpuregs[8][8] ;
 wire \cpuregs[8][9] ;
 wire \cpuregs[9][0] ;
 wire \cpuregs[9][10] ;
 wire \cpuregs[9][11] ;
 wire \cpuregs[9][12] ;
 wire \cpuregs[9][13] ;
 wire \cpuregs[9][14] ;
 wire \cpuregs[9][15] ;
 wire \cpuregs[9][16] ;
 wire \cpuregs[9][17] ;
 wire \cpuregs[9][18] ;
 wire \cpuregs[9][19] ;
 wire \cpuregs[9][1] ;
 wire \cpuregs[9][20] ;
 wire \cpuregs[9][21] ;
 wire \cpuregs[9][22] ;
 wire \cpuregs[9][23] ;
 wire \cpuregs[9][24] ;
 wire \cpuregs[9][25] ;
 wire \cpuregs[9][26] ;
 wire \cpuregs[9][27] ;
 wire \cpuregs[9][28] ;
 wire \cpuregs[9][29] ;
 wire \cpuregs[9][2] ;
 wire \cpuregs[9][30] ;
 wire \cpuregs[9][31] ;
 wire \cpuregs[9][3] ;
 wire \cpuregs[9][4] ;
 wire \cpuregs[9][5] ;
 wire \cpuregs[9][6] ;
 wire \cpuregs[9][7] ;
 wire \cpuregs[9][8] ;
 wire \cpuregs[9][9] ;
 wire \cpuregs_rs1[0] ;
 wire \cpuregs_rs1[10] ;
 wire \cpuregs_rs1[11] ;
 wire \cpuregs_rs1[12] ;
 wire \cpuregs_rs1[13] ;
 wire \cpuregs_rs1[14] ;
 wire \cpuregs_rs1[15] ;
 wire \cpuregs_rs1[16] ;
 wire \cpuregs_rs1[17] ;
 wire \cpuregs_rs1[18] ;
 wire \cpuregs_rs1[19] ;
 wire \cpuregs_rs1[1] ;
 wire \cpuregs_rs1[20] ;
 wire \cpuregs_rs1[21] ;
 wire \cpuregs_rs1[22] ;
 wire \cpuregs_rs1[23] ;
 wire \cpuregs_rs1[24] ;
 wire \cpuregs_rs1[25] ;
 wire \cpuregs_rs1[26] ;
 wire \cpuregs_rs1[27] ;
 wire \cpuregs_rs1[28] ;
 wire \cpuregs_rs1[29] ;
 wire \cpuregs_rs1[2] ;
 wire \cpuregs_rs1[30] ;
 wire \cpuregs_rs1[31] ;
 wire \cpuregs_rs1[3] ;
 wire \cpuregs_rs1[4] ;
 wire \cpuregs_rs1[5] ;
 wire \cpuregs_rs1[6] ;
 wire \cpuregs_rs1[7] ;
 wire \cpuregs_rs1[8] ;
 wire \cpuregs_rs1[9] ;
 wire \cpuregs_wrdata[0] ;
 wire \cpuregs_wrdata[10] ;
 wire \cpuregs_wrdata[11] ;
 wire \cpuregs_wrdata[12] ;
 wire \cpuregs_wrdata[13] ;
 wire \cpuregs_wrdata[14] ;
 wire \cpuregs_wrdata[15] ;
 wire \cpuregs_wrdata[16] ;
 wire \cpuregs_wrdata[17] ;
 wire \cpuregs_wrdata[18] ;
 wire \cpuregs_wrdata[19] ;
 wire \cpuregs_wrdata[1] ;
 wire \cpuregs_wrdata[20] ;
 wire \cpuregs_wrdata[21] ;
 wire \cpuregs_wrdata[22] ;
 wire \cpuregs_wrdata[23] ;
 wire \cpuregs_wrdata[24] ;
 wire \cpuregs_wrdata[25] ;
 wire \cpuregs_wrdata[26] ;
 wire \cpuregs_wrdata[27] ;
 wire \cpuregs_wrdata[28] ;
 wire \cpuregs_wrdata[29] ;
 wire \cpuregs_wrdata[2] ;
 wire \cpuregs_wrdata[30] ;
 wire \cpuregs_wrdata[31] ;
 wire \cpuregs_wrdata[3] ;
 wire \cpuregs_wrdata[4] ;
 wire \cpuregs_wrdata[5] ;
 wire \cpuregs_wrdata[6] ;
 wire \cpuregs_wrdata[7] ;
 wire \cpuregs_wrdata[8] ;
 wire \cpuregs_wrdata[9] ;
 wire \decoded_imm[0] ;
 wire \decoded_imm[10] ;
 wire \decoded_imm[11] ;
 wire \decoded_imm[12] ;
 wire \decoded_imm[13] ;
 wire \decoded_imm[14] ;
 wire \decoded_imm[15] ;
 wire \decoded_imm[16] ;
 wire \decoded_imm[17] ;
 wire \decoded_imm[18] ;
 wire \decoded_imm[19] ;
 wire \decoded_imm[1] ;
 wire \decoded_imm[20] ;
 wire \decoded_imm[21] ;
 wire \decoded_imm[22] ;
 wire \decoded_imm[23] ;
 wire \decoded_imm[24] ;
 wire \decoded_imm[25] ;
 wire \decoded_imm[26] ;
 wire \decoded_imm[27] ;
 wire \decoded_imm[28] ;
 wire \decoded_imm[29] ;
 wire \decoded_imm[2] ;
 wire \decoded_imm[30] ;
 wire \decoded_imm[31] ;
 wire \decoded_imm[3] ;
 wire \decoded_imm[4] ;
 wire \decoded_imm[5] ;
 wire \decoded_imm[6] ;
 wire \decoded_imm[7] ;
 wire \decoded_imm[8] ;
 wire \decoded_imm[9] ;
 wire \decoded_imm_uj[10] ;
 wire \decoded_imm_uj[11] ;
 wire \decoded_imm_uj[12] ;
 wire \decoded_imm_uj[13] ;
 wire \decoded_imm_uj[14] ;
 wire \decoded_imm_uj[15] ;
 wire \decoded_imm_uj[16] ;
 wire \decoded_imm_uj[17] ;
 wire \decoded_imm_uj[18] ;
 wire \decoded_imm_uj[19] ;
 wire \decoded_imm_uj[1] ;
 wire \decoded_imm_uj[20] ;
 wire \decoded_imm_uj[2] ;
 wire \decoded_imm_uj[3] ;
 wire \decoded_imm_uj[4] ;
 wire \decoded_imm_uj[5] ;
 wire \decoded_imm_uj[6] ;
 wire \decoded_imm_uj[7] ;
 wire \decoded_imm_uj[8] ;
 wire \decoded_imm_uj[9] ;
 wire \decoded_rd[0] ;
 wire \decoded_rd[1] ;
 wire \decoded_rd[2] ;
 wire \decoded_rd[3] ;
 wire \decoded_rd[4] ;
 wire \decoded_rs1[0] ;
 wire \decoded_rs1[1] ;
 wire \decoded_rs1[2] ;
 wire \decoded_rs1[3] ;
 wire \decoded_rs1[4] ;
 wire decoder_pseudo_trigger;
 wire decoder_trigger;
 wire do_waitirq;
 wire instr_add;
 wire instr_addi;
 wire instr_and;
 wire instr_andi;
 wire instr_auipc;
 wire instr_beq;
 wire instr_bge;
 wire instr_bgeu;
 wire instr_blt;
 wire instr_bltu;
 wire instr_bne;
 wire instr_ecall_ebreak;
 wire instr_getq;
 wire instr_jal;
 wire instr_jalr;
 wire instr_lb;
 wire instr_lbu;
 wire instr_lh;
 wire instr_lhu;
 wire instr_lui;
 wire instr_lw;
 wire instr_maskirq;
 wire instr_or;
 wire instr_ori;
 wire instr_rdcycle;
 wire instr_rdcycleh;
 wire instr_rdinstr;
 wire instr_rdinstrh;
 wire instr_retirq;
 wire instr_sb;
 wire instr_setq;
 wire instr_sh;
 wire instr_sll;
 wire instr_slli;
 wire instr_slt;
 wire instr_slti;
 wire instr_sltiu;
 wire instr_sltu;
 wire instr_sra;
 wire instr_srai;
 wire instr_srl;
 wire instr_srli;
 wire instr_sub;
 wire instr_sw;
 wire instr_timer;
 wire instr_waitirq;
 wire instr_xor;
 wire instr_xori;
 wire irq_active;
 wire irq_delay;
 wire \irq_mask[0] ;
 wire \irq_mask[10] ;
 wire \irq_mask[11] ;
 wire \irq_mask[12] ;
 wire \irq_mask[13] ;
 wire \irq_mask[14] ;
 wire \irq_mask[15] ;
 wire \irq_mask[16] ;
 wire \irq_mask[17] ;
 wire \irq_mask[18] ;
 wire \irq_mask[19] ;
 wire \irq_mask[1] ;
 wire \irq_mask[20] ;
 wire \irq_mask[21] ;
 wire \irq_mask[22] ;
 wire \irq_mask[23] ;
 wire \irq_mask[24] ;
 wire \irq_mask[25] ;
 wire \irq_mask[26] ;
 wire \irq_mask[27] ;
 wire \irq_mask[28] ;
 wire \irq_mask[29] ;
 wire \irq_mask[2] ;
 wire \irq_mask[30] ;
 wire \irq_mask[31] ;
 wire \irq_mask[3] ;
 wire \irq_mask[4] ;
 wire \irq_mask[5] ;
 wire \irq_mask[6] ;
 wire \irq_mask[7] ;
 wire \irq_mask[8] ;
 wire \irq_mask[9] ;
 wire \irq_pending[0] ;
 wire \irq_pending[10] ;
 wire \irq_pending[11] ;
 wire \irq_pending[12] ;
 wire \irq_pending[13] ;
 wire \irq_pending[14] ;
 wire \irq_pending[15] ;
 wire \irq_pending[16] ;
 wire \irq_pending[17] ;
 wire \irq_pending[18] ;
 wire \irq_pending[19] ;
 wire \irq_pending[1] ;
 wire \irq_pending[20] ;
 wire \irq_pending[21] ;
 wire \irq_pending[22] ;
 wire \irq_pending[23] ;
 wire \irq_pending[24] ;
 wire \irq_pending[25] ;
 wire \irq_pending[26] ;
 wire \irq_pending[27] ;
 wire \irq_pending[28] ;
 wire \irq_pending[29] ;
 wire \irq_pending[2] ;
 wire \irq_pending[30] ;
 wire \irq_pending[31] ;
 wire \irq_pending[3] ;
 wire \irq_pending[4] ;
 wire \irq_pending[5] ;
 wire \irq_pending[6] ;
 wire \irq_pending[7] ;
 wire \irq_pending[8] ;
 wire \irq_pending[9] ;
 wire \irq_state[0] ;
 wire \irq_state[1] ;
 wire is_alu_reg_imm;
 wire is_alu_reg_reg;
 wire is_beq_bne_blt_bge_bltu_bgeu;
 wire is_compare;
 wire is_jalr_addi_slti_sltiu_xori_ori_andi;
 wire is_lb_lh_lw_lbu_lhu;
 wire is_lui_auipc_jal;
 wire is_sb_sh_sw;
 wire is_slli_srli_srai;
 wire is_slti_blt_slt;
 wire is_sltiu_bltu_sltu;
 wire latched_branch;
 wire latched_is_lb;
 wire latched_is_lh;
 wire \latched_rd[0] ;
 wire \latched_rd[1] ;
 wire \latched_rd[2] ;
 wire \latched_rd[3] ;
 wire \latched_rd[4] ;
 wire latched_stalu;
 wire latched_store;
 wire mem_do_prefetch;
 wire mem_do_rdata;
 wire mem_do_rinst;
 wire mem_do_wdata;
 wire \mem_rdata_latched[10] ;
 wire \mem_rdata_latched[11] ;
 wire \mem_rdata_latched[12] ;
 wire \mem_rdata_latched[13] ;
 wire \mem_rdata_latched[14] ;
 wire \mem_rdata_latched[15] ;
 wire \mem_rdata_latched[16] ;
 wire \mem_rdata_latched[17] ;
 wire \mem_rdata_latched[18] ;
 wire \mem_rdata_latched[19] ;
 wire \mem_rdata_latched[20] ;
 wire \mem_rdata_latched[21] ;
 wire \mem_rdata_latched[22] ;
 wire \mem_rdata_latched[23] ;
 wire \mem_rdata_latched[24] ;
 wire \mem_rdata_latched[25] ;
 wire \mem_rdata_latched[26] ;
 wire \mem_rdata_latched[27] ;
 wire \mem_rdata_latched[28] ;
 wire \mem_rdata_latched[29] ;
 wire \mem_rdata_latched[30] ;
 wire \mem_rdata_latched[31] ;
 wire \mem_rdata_latched[7] ;
 wire \mem_rdata_latched[8] ;
 wire \mem_rdata_latched[9] ;
 wire \mem_rdata_q[0] ;
 wire \mem_rdata_q[10] ;
 wire \mem_rdata_q[11] ;
 wire \mem_rdata_q[12] ;
 wire \mem_rdata_q[13] ;
 wire \mem_rdata_q[14] ;
 wire \mem_rdata_q[15] ;
 wire \mem_rdata_q[16] ;
 wire \mem_rdata_q[17] ;
 wire \mem_rdata_q[18] ;
 wire \mem_rdata_q[19] ;
 wire \mem_rdata_q[1] ;
 wire \mem_rdata_q[20] ;
 wire \mem_rdata_q[21] ;
 wire \mem_rdata_q[22] ;
 wire \mem_rdata_q[23] ;
 wire \mem_rdata_q[24] ;
 wire \mem_rdata_q[25] ;
 wire \mem_rdata_q[26] ;
 wire \mem_rdata_q[27] ;
 wire \mem_rdata_q[28] ;
 wire \mem_rdata_q[29] ;
 wire \mem_rdata_q[2] ;
 wire \mem_rdata_q[30] ;
 wire \mem_rdata_q[31] ;
 wire \mem_rdata_q[3] ;
 wire \mem_rdata_q[4] ;
 wire \mem_rdata_q[5] ;
 wire \mem_rdata_q[6] ;
 wire \mem_rdata_q[7] ;
 wire \mem_rdata_q[8] ;
 wire \mem_rdata_q[9] ;
 wire \mem_state[0] ;
 wire \mem_state[1] ;
 wire \mem_wordsize[0] ;
 wire \mem_wordsize[1] ;
 wire \mem_wordsize[2] ;
 wire mem_xfer;
 wire \pcpi_mul.active[0] ;
 wire \pcpi_mul.active[1] ;
 wire \pcpi_mul.instr_any_mulh ;
 wire \pcpi_mul.rd[0] ;
 wire \pcpi_mul.rd[10] ;
 wire \pcpi_mul.rd[11] ;
 wire \pcpi_mul.rd[12] ;
 wire \pcpi_mul.rd[13] ;
 wire \pcpi_mul.rd[14] ;
 wire \pcpi_mul.rd[15] ;
 wire \pcpi_mul.rd[16] ;
 wire \pcpi_mul.rd[17] ;
 wire \pcpi_mul.rd[18] ;
 wire \pcpi_mul.rd[19] ;
 wire \pcpi_mul.rd[1] ;
 wire \pcpi_mul.rd[20] ;
 wire \pcpi_mul.rd[21] ;
 wire \pcpi_mul.rd[22] ;
 wire \pcpi_mul.rd[23] ;
 wire \pcpi_mul.rd[24] ;
 wire \pcpi_mul.rd[25] ;
 wire \pcpi_mul.rd[26] ;
 wire \pcpi_mul.rd[27] ;
 wire \pcpi_mul.rd[28] ;
 wire \pcpi_mul.rd[29] ;
 wire \pcpi_mul.rd[2] ;
 wire \pcpi_mul.rd[30] ;
 wire \pcpi_mul.rd[31] ;
 wire \pcpi_mul.rd[32] ;
 wire \pcpi_mul.rd[33] ;
 wire \pcpi_mul.rd[34] ;
 wire \pcpi_mul.rd[35] ;
 wire \pcpi_mul.rd[36] ;
 wire \pcpi_mul.rd[37] ;
 wire \pcpi_mul.rd[38] ;
 wire \pcpi_mul.rd[39] ;
 wire \pcpi_mul.rd[3] ;
 wire \pcpi_mul.rd[40] ;
 wire \pcpi_mul.rd[41] ;
 wire \pcpi_mul.rd[42] ;
 wire \pcpi_mul.rd[43] ;
 wire \pcpi_mul.rd[44] ;
 wire \pcpi_mul.rd[45] ;
 wire \pcpi_mul.rd[46] ;
 wire \pcpi_mul.rd[47] ;
 wire \pcpi_mul.rd[48] ;
 wire \pcpi_mul.rd[49] ;
 wire \pcpi_mul.rd[4] ;
 wire \pcpi_mul.rd[50] ;
 wire \pcpi_mul.rd[51] ;
 wire \pcpi_mul.rd[52] ;
 wire \pcpi_mul.rd[53] ;
 wire \pcpi_mul.rd[54] ;
 wire \pcpi_mul.rd[55] ;
 wire \pcpi_mul.rd[56] ;
 wire \pcpi_mul.rd[57] ;
 wire \pcpi_mul.rd[58] ;
 wire \pcpi_mul.rd[59] ;
 wire \pcpi_mul.rd[5] ;
 wire \pcpi_mul.rd[60] ;
 wire \pcpi_mul.rd[61] ;
 wire \pcpi_mul.rd[62] ;
 wire \pcpi_mul.rd[63] ;
 wire \pcpi_mul.rd[6] ;
 wire \pcpi_mul.rd[7] ;
 wire \pcpi_mul.rd[8] ;
 wire \pcpi_mul.rd[9] ;
 wire \pcpi_mul.rs1[0] ;
 wire \pcpi_mul.rs1[10] ;
 wire \pcpi_mul.rs1[11] ;
 wire \pcpi_mul.rs1[12] ;
 wire \pcpi_mul.rs1[13] ;
 wire \pcpi_mul.rs1[14] ;
 wire \pcpi_mul.rs1[15] ;
 wire \pcpi_mul.rs1[16] ;
 wire \pcpi_mul.rs1[17] ;
 wire \pcpi_mul.rs1[18] ;
 wire \pcpi_mul.rs1[19] ;
 wire \pcpi_mul.rs1[1] ;
 wire \pcpi_mul.rs1[20] ;
 wire \pcpi_mul.rs1[21] ;
 wire \pcpi_mul.rs1[22] ;
 wire \pcpi_mul.rs1[23] ;
 wire \pcpi_mul.rs1[24] ;
 wire \pcpi_mul.rs1[25] ;
 wire \pcpi_mul.rs1[26] ;
 wire \pcpi_mul.rs1[27] ;
 wire \pcpi_mul.rs1[28] ;
 wire \pcpi_mul.rs1[29] ;
 wire \pcpi_mul.rs1[2] ;
 wire \pcpi_mul.rs1[30] ;
 wire \pcpi_mul.rs1[31] ;
 wire \pcpi_mul.rs1[32] ;
 wire \pcpi_mul.rs1[3] ;
 wire \pcpi_mul.rs1[4] ;
 wire \pcpi_mul.rs1[5] ;
 wire \pcpi_mul.rs1[6] ;
 wire \pcpi_mul.rs1[7] ;
 wire \pcpi_mul.rs1[8] ;
 wire \pcpi_mul.rs1[9] ;
 wire \pcpi_mul.rs2[0] ;
 wire \pcpi_mul.rs2[10] ;
 wire \pcpi_mul.rs2[11] ;
 wire \pcpi_mul.rs2[12] ;
 wire \pcpi_mul.rs2[13] ;
 wire \pcpi_mul.rs2[14] ;
 wire \pcpi_mul.rs2[15] ;
 wire \pcpi_mul.rs2[16] ;
 wire \pcpi_mul.rs2[17] ;
 wire \pcpi_mul.rs2[18] ;
 wire \pcpi_mul.rs2[19] ;
 wire \pcpi_mul.rs2[1] ;
 wire \pcpi_mul.rs2[20] ;
 wire \pcpi_mul.rs2[21] ;
 wire \pcpi_mul.rs2[22] ;
 wire \pcpi_mul.rs2[23] ;
 wire \pcpi_mul.rs2[24] ;
 wire \pcpi_mul.rs2[25] ;
 wire \pcpi_mul.rs2[26] ;
 wire \pcpi_mul.rs2[27] ;
 wire \pcpi_mul.rs2[28] ;
 wire \pcpi_mul.rs2[29] ;
 wire \pcpi_mul.rs2[2] ;
 wire \pcpi_mul.rs2[30] ;
 wire \pcpi_mul.rs2[31] ;
 wire \pcpi_mul.rs2[32] ;
 wire \pcpi_mul.rs2[3] ;
 wire \pcpi_mul.rs2[4] ;
 wire \pcpi_mul.rs2[5] ;
 wire \pcpi_mul.rs2[6] ;
 wire \pcpi_mul.rs2[7] ;
 wire \pcpi_mul.rs2[8] ;
 wire \pcpi_mul.rs2[9] ;
 wire \pcpi_mul.shift_out ;
 wire pcpi_timeout;
 wire \pcpi_timeout_counter[0] ;
 wire \pcpi_timeout_counter[1] ;
 wire \pcpi_timeout_counter[2] ;
 wire \pcpi_timeout_counter[3] ;
 wire \reg_next_pc[0] ;
 wire \reg_next_pc[10] ;
 wire \reg_next_pc[11] ;
 wire \reg_next_pc[12] ;
 wire \reg_next_pc[13] ;
 wire \reg_next_pc[14] ;
 wire \reg_next_pc[15] ;
 wire \reg_next_pc[16] ;
 wire \reg_next_pc[17] ;
 wire \reg_next_pc[18] ;
 wire \reg_next_pc[19] ;
 wire \reg_next_pc[1] ;
 wire \reg_next_pc[20] ;
 wire \reg_next_pc[21] ;
 wire \reg_next_pc[22] ;
 wire \reg_next_pc[23] ;
 wire \reg_next_pc[24] ;
 wire \reg_next_pc[25] ;
 wire \reg_next_pc[26] ;
 wire \reg_next_pc[27] ;
 wire \reg_next_pc[28] ;
 wire \reg_next_pc[29] ;
 wire \reg_next_pc[2] ;
 wire \reg_next_pc[30] ;
 wire \reg_next_pc[31] ;
 wire \reg_next_pc[3] ;
 wire \reg_next_pc[4] ;
 wire \reg_next_pc[5] ;
 wire \reg_next_pc[6] ;
 wire \reg_next_pc[7] ;
 wire \reg_next_pc[8] ;
 wire \reg_next_pc[9] ;
 wire \reg_out[0] ;
 wire \reg_out[10] ;
 wire \reg_out[11] ;
 wire \reg_out[12] ;
 wire \reg_out[13] ;
 wire \reg_out[14] ;
 wire \reg_out[15] ;
 wire \reg_out[16] ;
 wire \reg_out[17] ;
 wire \reg_out[18] ;
 wire \reg_out[19] ;
 wire \reg_out[1] ;
 wire \reg_out[20] ;
 wire \reg_out[21] ;
 wire \reg_out[22] ;
 wire \reg_out[23] ;
 wire \reg_out[24] ;
 wire \reg_out[25] ;
 wire \reg_out[26] ;
 wire \reg_out[27] ;
 wire \reg_out[28] ;
 wire \reg_out[29] ;
 wire \reg_out[2] ;
 wire \reg_out[30] ;
 wire \reg_out[31] ;
 wire \reg_out[3] ;
 wire \reg_out[4] ;
 wire \reg_out[5] ;
 wire \reg_out[6] ;
 wire \reg_out[7] ;
 wire \reg_out[8] ;
 wire \reg_out[9] ;
 wire \reg_pc[10] ;
 wire \reg_pc[11] ;
 wire \reg_pc[12] ;
 wire \reg_pc[13] ;
 wire \reg_pc[14] ;
 wire \reg_pc[15] ;
 wire \reg_pc[16] ;
 wire \reg_pc[17] ;
 wire \reg_pc[18] ;
 wire \reg_pc[19] ;
 wire \reg_pc[1] ;
 wire \reg_pc[20] ;
 wire \reg_pc[21] ;
 wire \reg_pc[22] ;
 wire \reg_pc[23] ;
 wire \reg_pc[24] ;
 wire \reg_pc[25] ;
 wire \reg_pc[26] ;
 wire \reg_pc[27] ;
 wire \reg_pc[28] ;
 wire \reg_pc[29] ;
 wire \reg_pc[2] ;
 wire \reg_pc[30] ;
 wire \reg_pc[31] ;
 wire \reg_pc[3] ;
 wire \reg_pc[4] ;
 wire \reg_pc[5] ;
 wire \reg_pc[6] ;
 wire \reg_pc[7] ;
 wire \reg_pc[8] ;
 wire \reg_pc[9] ;
 wire \timer[0] ;
 wire \timer[10] ;
 wire \timer[11] ;
 wire \timer[12] ;
 wire \timer[13] ;
 wire \timer[14] ;
 wire \timer[15] ;
 wire \timer[16] ;
 wire \timer[17] ;
 wire \timer[18] ;
 wire \timer[19] ;
 wire \timer[1] ;
 wire \timer[20] ;
 wire \timer[21] ;
 wire \timer[22] ;
 wire \timer[23] ;
 wire \timer[24] ;
 wire \timer[25] ;
 wire \timer[26] ;
 wire \timer[27] ;
 wire \timer[28] ;
 wire \timer[29] ;
 wire \timer[2] ;
 wire \timer[30] ;
 wire \timer[31] ;
 wire \timer[3] ;
 wire \timer[4] ;
 wire \timer[5] ;
 wire \timer[6] ;
 wire \timer[7] ;
 wire \timer[8] ;
 wire \timer[9] ;

 sky130_fd_sc_hd__and2_2 _19867_ (.A(mem_valid),
    .B(mem_ready),
    .X(_16796_));
 sky130_fd_sc_hd__buf_1 _19868_ (.A(\mem_state[0] ),
    .X(_16797_));
 sky130_fd_sc_hd__and2_2 _19869_ (.A(\mem_state[1] ),
    .B(_16797_),
    .X(_16798_));
 sky130_fd_sc_hd__buf_1 _19870_ (.A(mem_do_rinst),
    .X(_16799_));
 sky130_fd_sc_hd__buf_1 _19871_ (.A(mem_ready),
    .X(_16800_));
 sky130_fd_sc_hd__o211a_2 _19872_ (.A1(mem_do_wdata),
    .A2(mem_do_rdata),
    .B1(mem_valid),
    .C1(_16800_),
    .X(_16801_));
 sky130_fd_sc_hd__nor2_2 _19873_ (.A(\mem_state[1] ),
    .B(\mem_state[0] ),
    .Y(_00290_));
 sky130_vsdinv _19874_ (.A(_00290_),
    .Y(_16802_));
 sky130_fd_sc_hd__o221ai_2 _19875_ (.A1(_16796_),
    .A2(_16798_),
    .B1(_16799_),
    .B2(_16801_),
    .C1(_16802_),
    .Y(_16803_));
 sky130_fd_sc_hd__buf_1 _19876_ (.A(_16803_),
    .X(_16804_));
 sky130_fd_sc_hd__buf_1 _19877_ (.A(mem_do_prefetch),
    .X(_16805_));
 sky130_fd_sc_hd__buf_1 _19878_ (.A(resetn),
    .X(_16806_));
 sky130_vsdinv _19879_ (.A(_16806_),
    .Y(_16807_));
 sky130_fd_sc_hd__buf_1 _19880_ (.A(_16807_),
    .X(_16808_));
 sky130_fd_sc_hd__buf_1 _19881_ (.A(_16808_),
    .X(_16809_));
 sky130_fd_sc_hd__a21oi_2 _19882_ (.A1(_16804_),
    .A2(_16805_),
    .B1(_16809_),
    .Y(_16810_));
 sky130_fd_sc_hd__buf_1 _19883_ (.A(mem_do_rdata),
    .X(_16811_));
 sky130_fd_sc_hd__and2_2 _19884_ (.A(_16811_),
    .B(\cpu_state[6] ),
    .X(_16812_));
 sky130_fd_sc_hd__buf_1 _19885_ (.A(_16812_),
    .X(_00319_));
 sky130_fd_sc_hd__a21oi_2 _19886_ (.A1(_16810_),
    .A2(_00319_),
    .B1(_00332_),
    .Y(_16813_));
 sky130_fd_sc_hd__buf_1 _19887_ (.A(_16806_),
    .X(_16814_));
 sky130_fd_sc_hd__buf_1 _19888_ (.A(_16814_),
    .X(_16815_));
 sky130_fd_sc_hd__buf_1 _19889_ (.A(_16815_),
    .X(_16816_));
 sky130_fd_sc_hd__buf_1 _19890_ (.A(_16816_),
    .X(_16817_));
 sky130_fd_sc_hd__buf_1 _19891_ (.A(_16817_),
    .X(_16818_));
 sky130_fd_sc_hd__buf_1 _19892_ (.A(_16818_),
    .X(_16819_));
 sky130_vsdinv _19893_ (.A(instr_lb),
    .Y(_16820_));
 sky130_fd_sc_hd__buf_1 _19894_ (.A(\cpu_state[6] ),
    .X(_16821_));
 sky130_vsdinv _19895_ (.A(_16821_),
    .Y(_16822_));
 sky130_fd_sc_hd__buf_1 _19896_ (.A(_16822_),
    .X(_16823_));
 sky130_fd_sc_hd__buf_1 _19897_ (.A(_16823_),
    .X(_16824_));
 sky130_fd_sc_hd__o21ai_2 _19898_ (.A1(_16820_),
    .A2(_16824_),
    .B1(_16813_),
    .Y(_16825_));
 sky130_fd_sc_hd__o211a_2 _19899_ (.A1(latched_is_lb),
    .A2(_16813_),
    .B1(_16819_),
    .C1(_16825_),
    .X(_04071_));
 sky130_vsdinv _19900_ (.A(instr_lh),
    .Y(_16826_));
 sky130_fd_sc_hd__o21ai_2 _19901_ (.A1(_16826_),
    .A2(_16824_),
    .B1(_16813_),
    .Y(_16827_));
 sky130_fd_sc_hd__o211a_2 _19902_ (.A1(latched_is_lh),
    .A2(_16813_),
    .B1(_16819_),
    .C1(_16827_),
    .X(_04070_));
 sky130_fd_sc_hd__buf_1 _19903_ (.A(\cpu_state[2] ),
    .X(_16828_));
 sky130_fd_sc_hd__buf_1 _19904_ (.A(_16828_),
    .X(_16829_));
 sky130_fd_sc_hd__and2b_2 _19905_ (.A_N(instr_retirq),
    .B(_16829_),
    .X(_16830_));
 sky130_fd_sc_hd__buf_1 _19906_ (.A(_16817_),
    .X(_16831_));
 sky130_fd_sc_hd__buf_1 _19907_ (.A(_16831_),
    .X(_16832_));
 sky130_fd_sc_hd__buf_1 _19908_ (.A(latched_branch),
    .X(_16833_));
 sky130_fd_sc_hd__o21bai_2 _19909_ (.A1(_00331_),
    .A2(_16830_),
    .B1_N(_16833_),
    .Y(_16834_));
 sky130_fd_sc_hd__o311a_2 _19910_ (.A1(_19816_),
    .A2(_00331_),
    .A3(_16830_),
    .B1(_16832_),
    .C1(_16834_),
    .X(_04069_));
 sky130_fd_sc_hd__buf_1 _19911_ (.A(\mem_state[1] ),
    .X(_16835_));
 sky130_fd_sc_hd__buf_1 _19912_ (.A(trap),
    .X(_16836_));
 sky130_fd_sc_hd__buf_1 _19913_ (.A(_16815_),
    .X(_16837_));
 sky130_fd_sc_hd__buf_1 _19914_ (.A(_16837_),
    .X(_16838_));
 sky130_fd_sc_hd__nand3b_2 _19915_ (.A_N(_16836_),
    .B(_16838_),
    .C(_19781_),
    .Y(_16839_));
 sky130_vsdinv _19916_ (.A(_16839_),
    .Y(_16840_));
 sky130_fd_sc_hd__buf_1 _19917_ (.A(_16808_),
    .X(_16841_));
 sky130_fd_sc_hd__buf_1 _19918_ (.A(_16841_),
    .X(_16842_));
 sky130_fd_sc_hd__nand3b_2 _19919_ (.A_N(_16797_),
    .B(mem_valid),
    .C(_16800_),
    .Y(_16843_));
 sky130_fd_sc_hd__buf_1 _19920_ (.A(_16797_),
    .X(_16844_));
 sky130_fd_sc_hd__buf_1 _19921_ (.A(_16799_),
    .X(_16845_));
 sky130_fd_sc_hd__nand2_2 _19922_ (.A(_16844_),
    .B(_16845_),
    .Y(_16846_));
 sky130_fd_sc_hd__nor2_2 _19923_ (.A(_16799_),
    .B(mem_do_prefetch),
    .Y(_16847_));
 sky130_fd_sc_hd__buf_1 _19924_ (.A(mem_do_wdata),
    .X(_16848_));
 sky130_fd_sc_hd__inv_2 _19925_ (.A(_16848_),
    .Y(_00291_));
 sky130_vsdinv _19926_ (.A(_16811_),
    .Y(_16849_));
 sky130_fd_sc_hd__nand3_2 _19927_ (.A(_16847_),
    .B(_00291_),
    .C(_16849_),
    .Y(_16850_));
 sky130_fd_sc_hd__nor2_2 _19928_ (.A(_16802_),
    .B(_16850_),
    .Y(_16851_));
 sky130_fd_sc_hd__a311oi_2 _19929_ (.A1(_16835_),
    .A2(_16843_),
    .A3(_16846_),
    .B1(trap),
    .C1(_16851_),
    .Y(_16852_));
 sky130_fd_sc_hd__o21a_2 _19930_ (.A1(_16842_),
    .A2(_16852_),
    .B1(_00300_),
    .X(_16853_));
 sky130_fd_sc_hd__mux2_2 _19931_ (.A0(_16835_),
    .A1(_16840_),
    .S(_16853_),
    .X(_04068_));
 sky130_fd_sc_hd__buf_1 _19932_ (.A(_16815_),
    .X(_16854_));
 sky130_fd_sc_hd__and2b_2 _19933_ (.A_N(_16836_),
    .B(_16854_),
    .X(_16855_));
 sky130_fd_sc_hd__buf_1 _19934_ (.A(_16855_),
    .X(_16856_));
 sky130_fd_sc_hd__and2b_2 _19935_ (.A_N(_16853_),
    .B(_16844_),
    .X(_16857_));
 sky130_fd_sc_hd__a31o_2 _19936_ (.A1(_19780_),
    .A2(_16853_),
    .A3(_16856_),
    .B1(_16857_),
    .X(_04067_));
 sky130_vsdinv _19937_ (.A(_16845_),
    .Y(_16858_));
 sky130_fd_sc_hd__nor3_2 _19938_ (.A(_16808_),
    .B(_16858_),
    .C(_16804_),
    .Y(_16859_));
 sky130_fd_sc_hd__buf_1 _19939_ (.A(_16859_),
    .X(_16860_));
 sky130_fd_sc_hd__buf_1 _19940_ (.A(_16860_),
    .X(_16861_));
 sky130_fd_sc_hd__buf_1 _19941_ (.A(_16861_),
    .X(_19783_));
 sky130_fd_sc_hd__inv_2 _19942_ (.A(\decoded_rs1[4] ),
    .Y(_00366_));
 sky130_fd_sc_hd__buf_1 _19943_ (.A(_16860_),
    .X(_16862_));
 sky130_fd_sc_hd__buf_1 _19944_ (.A(_16862_),
    .X(_16863_));
 sky130_fd_sc_hd__or3_2 _19945_ (.A(\mem_rdata_latched[31] ),
    .B(\mem_rdata_latched[30] ),
    .C(\mem_rdata_latched[29] ),
    .X(_16864_));
 sky130_fd_sc_hd__or2b_2 _19946_ (.A(\mem_rdata_latched[25] ),
    .B_N(\mem_rdata_latched[26] ),
    .X(_16865_));
 sky130_fd_sc_hd__nand3b_2 _19947_ (.A_N(_00326_),
    .B(_00325_),
    .C(_00324_),
    .Y(_16866_));
 sky130_fd_sc_hd__nor2_2 _19948_ (.A(_00329_),
    .B(_00328_),
    .Y(_16867_));
 sky130_fd_sc_hd__nor3b_2 _19949_ (.A(\mem_rdata_latched[28] ),
    .B(_00330_),
    .C_N(_00327_),
    .Y(_16868_));
 sky130_fd_sc_hd__nand3b_2 _19950_ (.A_N(_16866_),
    .B(_16867_),
    .C(_16868_),
    .Y(_16869_));
 sky130_fd_sc_hd__or2_2 _19951_ (.A(\mem_rdata_latched[27] ),
    .B(_16869_),
    .X(_16870_));
 sky130_fd_sc_hd__nor3_2 _19952_ (.A(_16864_),
    .B(_16865_),
    .C(_16870_),
    .Y(_16871_));
 sky130_fd_sc_hd__buf_1 _19953_ (.A(_16860_),
    .X(_16872_));
 sky130_fd_sc_hd__nand2_2 _19954_ (.A(_16871_),
    .B(_16872_),
    .Y(_16873_));
 sky130_fd_sc_hd__or3_2 _19955_ (.A(\mem_rdata_latched[26] ),
    .B(\mem_rdata_latched[25] ),
    .C(_16864_),
    .X(_16874_));
 sky130_fd_sc_hd__nor2_2 _19956_ (.A(_16870_),
    .B(_16874_),
    .Y(_16875_));
 sky130_fd_sc_hd__buf_1 _19957_ (.A(_16861_),
    .X(_16876_));
 sky130_fd_sc_hd__o21ai_2 _19958_ (.A1(\mem_rdata_latched[19] ),
    .A2(_16875_),
    .B1(_16876_),
    .Y(_16877_));
 sky130_fd_sc_hd__o211ai_2 _19959_ (.A1(_00366_),
    .A2(_16863_),
    .B1(_16873_),
    .C1(_16877_),
    .Y(_04066_));
 sky130_vsdinv _19960_ (.A(irq_delay),
    .Y(_16878_));
 sky130_vsdinv _19961_ (.A(instr_waitirq),
    .Y(_16879_));
 sky130_fd_sc_hd__nor2_2 _19962_ (.A(decoder_trigger),
    .B(do_waitirq),
    .Y(_16880_));
 sky130_fd_sc_hd__nor2_2 _19963_ (.A(\irq_state[1] ),
    .B(\irq_state[0] ),
    .Y(_16881_));
 sky130_vsdinv _19964_ (.A(\irq_mask[11] ),
    .Y(_16882_));
 sky130_fd_sc_hd__and2b_2 _19965_ (.A_N(\irq_mask[8] ),
    .B(\irq_pending[8] ),
    .X(_16883_));
 sky130_fd_sc_hd__and2b_2 _19966_ (.A_N(\irq_mask[10] ),
    .B(\irq_pending[10] ),
    .X(_16884_));
 sky130_fd_sc_hd__and2b_2 _19967_ (.A_N(\irq_mask[9] ),
    .B(\irq_pending[9] ),
    .X(_16885_));
 sky130_fd_sc_hd__a2111oi_2 _19968_ (.A1(_16882_),
    .A2(\irq_pending[11] ),
    .B1(_16883_),
    .C1(_16884_),
    .D1(_16885_),
    .Y(_16886_));
 sky130_vsdinv _19969_ (.A(\irq_mask[2] ),
    .Y(_16887_));
 sky130_fd_sc_hd__and2b_2 _19970_ (.A_N(\irq_mask[0] ),
    .B(\irq_pending[0] ),
    .X(_16888_));
 sky130_fd_sc_hd__and2b_2 _19971_ (.A_N(\irq_mask[3] ),
    .B(\irq_pending[3] ),
    .X(_16889_));
 sky130_fd_sc_hd__and2b_2 _19972_ (.A_N(\irq_mask[1] ),
    .B(\irq_pending[1] ),
    .X(_16890_));
 sky130_fd_sc_hd__a2111oi_2 _19973_ (.A1(_16887_),
    .A2(\irq_pending[2] ),
    .B1(_16888_),
    .C1(_16889_),
    .D1(_16890_),
    .Y(_16891_));
 sky130_vsdinv _19974_ (.A(\irq_mask[23] ),
    .Y(_16892_));
 sky130_fd_sc_hd__and2b_2 _19975_ (.A_N(\irq_mask[20] ),
    .B(\irq_pending[20] ),
    .X(_16893_));
 sky130_fd_sc_hd__and2b_2 _19976_ (.A_N(\irq_mask[22] ),
    .B(\irq_pending[22] ),
    .X(_16894_));
 sky130_fd_sc_hd__and2b_2 _19977_ (.A_N(\irq_mask[21] ),
    .B(\irq_pending[21] ),
    .X(_16895_));
 sky130_fd_sc_hd__a2111oi_2 _19978_ (.A1(_16892_),
    .A2(\irq_pending[23] ),
    .B1(_16893_),
    .C1(_16894_),
    .D1(_16895_),
    .Y(_16896_));
 sky130_vsdinv _19979_ (.A(\irq_mask[7] ),
    .Y(_16897_));
 sky130_fd_sc_hd__and2b_2 _19980_ (.A_N(\irq_mask[4] ),
    .B(\irq_pending[4] ),
    .X(_16898_));
 sky130_fd_sc_hd__and2b_2 _19981_ (.A_N(\irq_mask[6] ),
    .B(\irq_pending[6] ),
    .X(_16899_));
 sky130_fd_sc_hd__and2b_2 _19982_ (.A_N(\irq_mask[5] ),
    .B(\irq_pending[5] ),
    .X(_16900_));
 sky130_fd_sc_hd__a2111oi_2 _19983_ (.A1(_16897_),
    .A2(\irq_pending[7] ),
    .B1(_16898_),
    .C1(_16899_),
    .D1(_16900_),
    .Y(_16901_));
 sky130_fd_sc_hd__and4_2 _19984_ (.A(_16886_),
    .B(_16891_),
    .C(_16896_),
    .D(_16901_),
    .X(_16902_));
 sky130_fd_sc_hd__and2b_2 _19985_ (.A_N(\irq_mask[16] ),
    .B(\irq_pending[16] ),
    .X(_16903_));
 sky130_fd_sc_hd__and2b_2 _19986_ (.A_N(\irq_mask[18] ),
    .B(\irq_pending[18] ),
    .X(_16904_));
 sky130_fd_sc_hd__and2b_2 _19987_ (.A_N(\irq_mask[19] ),
    .B(\irq_pending[19] ),
    .X(_16905_));
 sky130_fd_sc_hd__and2b_2 _19988_ (.A_N(\irq_mask[17] ),
    .B(\irq_pending[17] ),
    .X(_16906_));
 sky130_fd_sc_hd__or4_2 _19989_ (.A(_16903_),
    .B(_16904_),
    .C(_16905_),
    .D(_16906_),
    .X(_16907_));
 sky130_fd_sc_hd__and2b_2 _19990_ (.A_N(\irq_mask[28] ),
    .B(\irq_pending[28] ),
    .X(_16908_));
 sky130_fd_sc_hd__and2b_2 _19991_ (.A_N(\irq_mask[30] ),
    .B(\irq_pending[30] ),
    .X(_16909_));
 sky130_fd_sc_hd__and2b_2 _19992_ (.A_N(\irq_mask[31] ),
    .B(\irq_pending[31] ),
    .X(_16910_));
 sky130_fd_sc_hd__and2b_2 _19993_ (.A_N(\irq_mask[29] ),
    .B(\irq_pending[29] ),
    .X(_16911_));
 sky130_fd_sc_hd__or4_2 _19994_ (.A(_16908_),
    .B(_16909_),
    .C(_16910_),
    .D(_16911_),
    .X(_16912_));
 sky130_fd_sc_hd__nor2_2 _19995_ (.A(_16907_),
    .B(_16912_),
    .Y(_16913_));
 sky130_vsdinv _19996_ (.A(\irq_mask[27] ),
    .Y(_16914_));
 sky130_fd_sc_hd__and2b_2 _19997_ (.A_N(\irq_mask[24] ),
    .B(\irq_pending[24] ),
    .X(_16915_));
 sky130_fd_sc_hd__and2b_2 _19998_ (.A_N(\irq_mask[26] ),
    .B(\irq_pending[26] ),
    .X(_16916_));
 sky130_fd_sc_hd__and2b_2 _19999_ (.A_N(\irq_mask[25] ),
    .B(\irq_pending[25] ),
    .X(_16917_));
 sky130_fd_sc_hd__a2111oi_2 _20000_ (.A1(_16914_),
    .A2(\irq_pending[27] ),
    .B1(_16915_),
    .C1(_16916_),
    .D1(_16917_),
    .Y(_16918_));
 sky130_vsdinv _20001_ (.A(\irq_mask[15] ),
    .Y(_16919_));
 sky130_fd_sc_hd__and2b_2 _20002_ (.A_N(\irq_mask[12] ),
    .B(\irq_pending[12] ),
    .X(_16920_));
 sky130_fd_sc_hd__and2b_2 _20003_ (.A_N(\irq_mask[14] ),
    .B(\irq_pending[14] ),
    .X(_16921_));
 sky130_fd_sc_hd__and2b_2 _20004_ (.A_N(\irq_mask[13] ),
    .B(\irq_pending[13] ),
    .X(_16922_));
 sky130_fd_sc_hd__a2111oi_2 _20005_ (.A1(_16919_),
    .A2(\irq_pending[15] ),
    .B1(_16920_),
    .C1(_16921_),
    .D1(_16922_),
    .Y(_16923_));
 sky130_fd_sc_hd__nand3b_2 _20006_ (.A_N(irq_active),
    .B(_16878_),
    .C(decoder_trigger),
    .Y(_16924_));
 sky130_fd_sc_hd__a41o_2 _20007_ (.A1(_16902_),
    .A2(_16913_),
    .A3(_16918_),
    .A4(_16923_),
    .B1(_16924_),
    .X(_16925_));
 sky130_fd_sc_hd__o211a_2 _20008_ (.A1(_16879_),
    .A2(_16880_),
    .B1(_16881_),
    .C1(_16925_),
    .X(_16926_));
 sky130_fd_sc_hd__buf_1 _20009_ (.A(decoder_trigger),
    .X(_16927_));
 sky130_fd_sc_hd__nand3_2 _20010_ (.A(_16926_),
    .B(\cpu_state[1] ),
    .C(_16927_),
    .Y(_16928_));
 sky130_fd_sc_hd__buf_1 _20011_ (.A(_16928_),
    .X(_16929_));
 sky130_fd_sc_hd__buf_1 _20012_ (.A(_16807_),
    .X(_16930_));
 sky130_fd_sc_hd__buf_1 _20013_ (.A(_16930_),
    .X(_16931_));
 sky130_fd_sc_hd__buf_1 _20014_ (.A(_16931_),
    .X(_16932_));
 sky130_fd_sc_hd__buf_1 _20015_ (.A(_16932_),
    .X(_16933_));
 sky130_fd_sc_hd__buf_1 _20016_ (.A(_16933_),
    .X(_16934_));
 sky130_fd_sc_hd__buf_1 _20017_ (.A(irq_active),
    .X(_16935_));
 sky130_fd_sc_hd__buf_1 _20018_ (.A(_16935_),
    .X(_16936_));
 sky130_fd_sc_hd__nor2_2 _20019_ (.A(_16936_),
    .B(_16929_),
    .Y(_16937_));
 sky130_fd_sc_hd__a211oi_2 _20020_ (.A1(_16878_),
    .A2(_16929_),
    .B1(_16934_),
    .C1(_16937_),
    .Y(_04065_));
 sky130_fd_sc_hd__buf_1 _20021_ (.A(pcpi_insn[13]),
    .X(_16938_));
 sky130_fd_sc_hd__nand3b_2 _20022_ (.A_N(pcpi_insn[2]),
    .B(pcpi_insn[1]),
    .C(pcpi_insn[0]),
    .Y(_16939_));
 sky130_fd_sc_hd__nor2_2 _20023_ (.A(pcpi_insn[27]),
    .B(pcpi_insn[26]),
    .Y(_16940_));
 sky130_fd_sc_hd__nand3b_2 _20024_ (.A_N(pcpi_insn[14]),
    .B(_16940_),
    .C(pcpi_insn[25]),
    .Y(_16941_));
 sky130_fd_sc_hd__and2b_2 _20025_ (.A_N(pcpi_insn[3]),
    .B(pcpi_insn[4]),
    .X(_16942_));
 sky130_fd_sc_hd__nand3b_2 _20026_ (.A_N(pcpi_insn[6]),
    .B(_16942_),
    .C(pcpi_insn[5]),
    .Y(_16943_));
 sky130_fd_sc_hd__nor3_2 _20027_ (.A(_16939_),
    .B(_16941_),
    .C(_16943_),
    .Y(_16944_));
 sky130_fd_sc_hd__and2_2 _20028_ (.A(_16806_),
    .B(pcpi_valid),
    .X(_16945_));
 sky130_fd_sc_hd__nor2_2 _20029_ (.A(pcpi_insn[31]),
    .B(pcpi_insn[30]),
    .Y(_16946_));
 sky130_fd_sc_hd__nor2_2 _20030_ (.A(pcpi_insn[29]),
    .B(pcpi_insn[28]),
    .Y(_16947_));
 sky130_fd_sc_hd__and3_2 _20031_ (.A(_16945_),
    .B(_16946_),
    .C(_16947_),
    .X(_16948_));
 sky130_fd_sc_hd__nand3_2 _20032_ (.A(_16944_),
    .B(pcpi_insn[12]),
    .C(_16948_),
    .Y(_16949_));
 sky130_fd_sc_hd__and2_2 _20033_ (.A(_16944_),
    .B(_16948_),
    .X(_16950_));
 sky130_fd_sc_hd__nand3b_2 _20034_ (.A_N(pcpi_insn[12]),
    .B(_16950_),
    .C(pcpi_insn[13]),
    .Y(_16951_));
 sky130_fd_sc_hd__o21ai_2 _20035_ (.A1(_16938_),
    .A2(_16949_),
    .B1(_16951_),
    .Y(_16952_));
 sky130_vsdinv _20036_ (.A(\pcpi_mul.active[0] ),
    .Y(_16953_));
 sky130_vsdinv _20037_ (.A(\pcpi_mul.active[1] ),
    .Y(_16954_));
 sky130_fd_sc_hd__and4_2 _20038_ (.A(_16944_),
    .B(_16953_),
    .C(_16954_),
    .D(_16948_),
    .X(_16955_));
 sky130_fd_sc_hd__buf_1 _20039_ (.A(_16955_),
    .X(_16956_));
 sky130_fd_sc_hd__buf_1 _20040_ (.A(pcpi_rs1[31]),
    .X(_16957_));
 sky130_fd_sc_hd__buf_1 _20041_ (.A(_16957_),
    .X(_16958_));
 sky130_fd_sc_hd__and2_2 _20042_ (.A(_16956_),
    .B(_16958_),
    .X(_16959_));
 sky130_fd_sc_hd__buf_1 _20043_ (.A(\pcpi_mul.rs1[32] ),
    .X(_16960_));
 sky130_fd_sc_hd__buf_1 _20044_ (.A(_16960_),
    .X(_16961_));
 sky130_vsdinv _20045_ (.A(_16961_),
    .Y(_16962_));
 sky130_fd_sc_hd__buf_1 _20046_ (.A(_16962_),
    .X(_16963_));
 sky130_fd_sc_hd__buf_1 _20047_ (.A(_16955_),
    .X(_16964_));
 sky130_fd_sc_hd__buf_1 _20048_ (.A(_16964_),
    .X(_16965_));
 sky130_fd_sc_hd__buf_1 _20049_ (.A(_16965_),
    .X(_16966_));
 sky130_fd_sc_hd__o2bb2ai_2 _20050_ (.A1_N(_16952_),
    .A2_N(_16959_),
    .B1(_16963_),
    .B2(_16966_),
    .Y(_04064_));
 sky130_vsdinv _20051_ (.A(\pcpi_mul.rs2[32] ),
    .Y(_16967_));
 sky130_fd_sc_hd__buf_1 _20052_ (.A(_16967_),
    .X(_16968_));
 sky130_fd_sc_hd__buf_1 _20053_ (.A(_16968_),
    .X(_16969_));
 sky130_fd_sc_hd__buf_1 _20054_ (.A(_16969_),
    .X(_16970_));
 sky130_fd_sc_hd__buf_1 _20055_ (.A(_16970_),
    .X(_16971_));
 sky130_fd_sc_hd__buf_1 _20056_ (.A(_16971_),
    .X(_16972_));
 sky130_fd_sc_hd__buf_1 _20057_ (.A(_16972_),
    .X(_16973_));
 sky130_fd_sc_hd__buf_1 _20058_ (.A(_16964_),
    .X(_16974_));
 sky130_fd_sc_hd__buf_1 _20059_ (.A(_16974_),
    .X(_03728_));
 sky130_fd_sc_hd__buf_1 _20060_ (.A(_16956_),
    .X(_16975_));
 sky130_fd_sc_hd__nor2_2 _20061_ (.A(_16938_),
    .B(_16949_),
    .Y(_16976_));
 sky130_fd_sc_hd__buf_1 _20062_ (.A(pcpi_rs2[31]),
    .X(_16977_));
 sky130_fd_sc_hd__buf_1 _20063_ (.A(_16977_),
    .X(_16978_));
 sky130_fd_sc_hd__nand3_2 _20064_ (.A(_16975_),
    .B(_16976_),
    .C(_16978_),
    .Y(_16979_));
 sky130_fd_sc_hd__o21ai_2 _20065_ (.A1(_16973_),
    .A2(_03728_),
    .B1(_16979_),
    .Y(_04063_));
 sky130_fd_sc_hd__inv_2 _20066_ (.A(alu_wait),
    .Y(_00302_));
 sky130_fd_sc_hd__buf_1 _20067_ (.A(is_beq_bne_blt_bge_bltu_bgeu),
    .X(_16980_));
 sky130_fd_sc_hd__buf_1 _20068_ (.A(_16980_),
    .X(_16981_));
 sky130_fd_sc_hd__a21boi_2 _20069_ (.A1(_00302_),
    .A2(_16981_),
    .B1_N(_00333_),
    .Y(_16982_));
 sky130_vsdinv _20070_ (.A(\cpu_state[4] ),
    .Y(_16983_));
 sky130_fd_sc_hd__buf_1 _20071_ (.A(_16983_),
    .X(_16984_));
 sky130_fd_sc_hd__buf_1 _20072_ (.A(_16984_),
    .X(_16985_));
 sky130_fd_sc_hd__nand2_2 _20073_ (.A(_16985_),
    .B(_00333_),
    .Y(_16986_));
 sky130_fd_sc_hd__o211a_2 _20074_ (.A1(latched_stalu),
    .A2(_16982_),
    .B1(_16819_),
    .C1(_16986_),
    .X(_04062_));
 sky130_fd_sc_hd__buf_1 _20075_ (.A(latched_store),
    .X(_16987_));
 sky130_fd_sc_hd__nor2_2 _20076_ (.A(instr_auipc),
    .B(instr_lui),
    .Y(_16988_));
 sky130_vsdinv _20077_ (.A(instr_jal),
    .Y(_16989_));
 sky130_fd_sc_hd__nand2_2 _20078_ (.A(_16988_),
    .B(_16989_),
    .Y(_00005_));
 sky130_fd_sc_hd__nor2_2 _20079_ (.A(instr_sra),
    .B(instr_srai),
    .Y(_16990_));
 sky130_vsdinv _20080_ (.A(instr_srl),
    .Y(_16991_));
 sky130_vsdinv _20081_ (.A(instr_srli),
    .Y(_16992_));
 sky130_fd_sc_hd__and3_2 _20082_ (.A(_16990_),
    .B(_16991_),
    .C(_16992_),
    .X(_16993_));
 sky130_vsdinv _20083_ (.A(_16993_),
    .Y(_16994_));
 sky130_fd_sc_hd__or4_2 _20084_ (.A(instr_lw),
    .B(instr_lh),
    .C(instr_lb),
    .D(instr_jalr),
    .X(_16995_));
 sky130_fd_sc_hd__or4_2 _20085_ (.A(instr_sh),
    .B(instr_sb),
    .C(instr_lhu),
    .D(instr_lbu),
    .X(_16996_));
 sky130_fd_sc_hd__or4_2 _20086_ (.A(_00005_),
    .B(_16994_),
    .C(_16995_),
    .D(_16996_),
    .X(_16997_));
 sky130_fd_sc_hd__or4_2 _20087_ (.A(instr_andi),
    .B(instr_ori),
    .C(instr_xori),
    .D(instr_addi),
    .X(_16998_));
 sky130_fd_sc_hd__or4_2 _20088_ (.A(instr_slt),
    .B(instr_sll),
    .C(instr_sub),
    .D(instr_add),
    .X(_16999_));
 sky130_fd_sc_hd__or4_2 _20089_ (.A(instr_timer),
    .B(instr_waitirq),
    .C(instr_slli),
    .D(instr_sw),
    .X(_17000_));
 sky130_fd_sc_hd__or4_2 _20090_ (.A(instr_bltu),
    .B(instr_blt),
    .C(instr_bne),
    .D(instr_beq),
    .X(_17001_));
 sky130_fd_sc_hd__or4_2 _20091_ (.A(_16998_),
    .B(_16999_),
    .C(_17000_),
    .D(_17001_),
    .X(_17002_));
 sky130_fd_sc_hd__nor2_2 _20092_ (.A(_16997_),
    .B(_17002_),
    .Y(_17003_));
 sky130_fd_sc_hd__buf_1 _20093_ (.A(_17003_),
    .X(_17004_));
 sky130_fd_sc_hd__nor2_2 _20094_ (.A(instr_setq),
    .B(instr_getq),
    .Y(_17005_));
 sky130_vsdinv _20095_ (.A(instr_maskirq),
    .Y(_17006_));
 sky130_vsdinv _20096_ (.A(instr_retirq),
    .Y(_17007_));
 sky130_fd_sc_hd__nand3_2 _20097_ (.A(_17005_),
    .B(_17006_),
    .C(_17007_),
    .Y(_17008_));
 sky130_fd_sc_hd__nor3_2 _20098_ (.A(instr_rdinstrh),
    .B(instr_rdinstr),
    .C(instr_rdcycleh),
    .Y(_01714_));
 sky130_fd_sc_hd__or2b_2 _20099_ (.A(instr_rdcycle),
    .B_N(_01714_),
    .X(_17009_));
 sky130_fd_sc_hd__or4_2 _20100_ (.A(instr_and),
    .B(instr_or),
    .C(instr_xor),
    .D(instr_sltu),
    .X(_17010_));
 sky130_fd_sc_hd__nor2_2 _20101_ (.A(instr_sltiu),
    .B(instr_slti),
    .Y(_17011_));
 sky130_fd_sc_hd__nor2_2 _20102_ (.A(instr_bgeu),
    .B(instr_bge),
    .Y(_17012_));
 sky130_fd_sc_hd__nand3b_2 _20103_ (.A_N(_17010_),
    .B(_17011_),
    .C(_17012_),
    .Y(_17013_));
 sky130_fd_sc_hd__nor3_2 _20104_ (.A(_17008_),
    .B(_17009_),
    .C(_17013_),
    .Y(_17014_));
 sky130_fd_sc_hd__buf_1 _20105_ (.A(_17014_),
    .X(_17015_));
 sky130_fd_sc_hd__nand3_2 _20106_ (.A(_17004_),
    .B(\pcpi_mul.active[1] ),
    .C(_17015_),
    .Y(_17016_));
 sky130_fd_sc_hd__buf_1 _20107_ (.A(\cpu_state[3] ),
    .X(_17017_));
 sky130_fd_sc_hd__buf_1 _20108_ (.A(_17017_),
    .X(_17018_));
 sky130_fd_sc_hd__buf_1 _20109_ (.A(\cpu_state[2] ),
    .X(_17019_));
 sky130_vsdinv _20110_ (.A(_17019_),
    .Y(_17020_));
 sky130_fd_sc_hd__buf_1 _20111_ (.A(_17020_),
    .X(_17021_));
 sky130_fd_sc_hd__buf_1 _20112_ (.A(instr_timer),
    .X(_17022_));
 sky130_fd_sc_hd__nor2_2 _20113_ (.A(_17022_),
    .B(_17008_),
    .Y(_01717_));
 sky130_fd_sc_hd__nor3b_2 _20114_ (.A(_17021_),
    .B(_17009_),
    .C_N(_01717_),
    .Y(_17023_));
 sky130_fd_sc_hd__and2_2 _20115_ (.A(\cpu_state[4] ),
    .B(alu_wait),
    .X(_17024_));
 sky130_fd_sc_hd__buf_1 _20116_ (.A(\cpu_state[1] ),
    .X(_17025_));
 sky130_fd_sc_hd__buf_1 _20117_ (.A(_17025_),
    .X(_17026_));
 sky130_fd_sc_hd__buf_1 _20118_ (.A(_17026_),
    .X(_17027_));
 sky130_fd_sc_hd__nor2_2 _20119_ (.A(_17019_),
    .B(\cpu_state[3] ),
    .Y(_17028_));
 sky130_fd_sc_hd__nand3_2 _20120_ (.A(_17028_),
    .B(_16983_),
    .C(_16822_),
    .Y(_17029_));
 sky130_fd_sc_hd__nor2_2 _20121_ (.A(_17027_),
    .B(_17029_),
    .Y(_17030_));
 sky130_fd_sc_hd__a2111oi_2 _20122_ (.A1(_17016_),
    .A2(_17018_),
    .B1(_17023_),
    .C1(_17024_),
    .D1(_17030_),
    .Y(_17031_));
 sky130_fd_sc_hd__or2b_2 _20123_ (.A(_19817_),
    .B_N(_17031_),
    .X(_17032_));
 sky130_fd_sc_hd__o211a_2 _20124_ (.A1(_16987_),
    .A2(_17031_),
    .B1(_16819_),
    .C1(_17032_),
    .X(_04061_));
 sky130_fd_sc_hd__buf_1 _20125_ (.A(\irq_state[1] ),
    .X(_17033_));
 sky130_fd_sc_hd__buf_1 _20126_ (.A(_17033_),
    .X(_17034_));
 sky130_fd_sc_hd__buf_1 _20127_ (.A(_17034_),
    .X(_17035_));
 sky130_fd_sc_hd__buf_1 _20128_ (.A(\irq_state[0] ),
    .X(_17036_));
 sky130_fd_sc_hd__buf_1 _20129_ (.A(_17036_),
    .X(_17037_));
 sky130_fd_sc_hd__buf_1 _20130_ (.A(_17037_),
    .X(_17038_));
 sky130_fd_sc_hd__buf_1 _20131_ (.A(_17027_),
    .X(_17039_));
 sky130_fd_sc_hd__buf_1 _20132_ (.A(_17039_),
    .X(_17040_));
 sky130_fd_sc_hd__nand3b_2 _20133_ (.A_N(_17035_),
    .B(_17038_),
    .C(_17040_),
    .Y(_17041_));
 sky130_vsdinv _20134_ (.A(_17025_),
    .Y(_17042_));
 sky130_fd_sc_hd__buf_1 _20135_ (.A(_17042_),
    .X(_17043_));
 sky130_fd_sc_hd__buf_1 _20136_ (.A(_17043_),
    .X(_17044_));
 sky130_fd_sc_hd__buf_1 _20137_ (.A(_17044_),
    .X(_17045_));
 sky130_fd_sc_hd__buf_1 _20138_ (.A(_17034_),
    .X(_17046_));
 sky130_fd_sc_hd__nand2_2 _20139_ (.A(_17045_),
    .B(_17046_),
    .Y(_17047_));
 sky130_fd_sc_hd__buf_1 _20140_ (.A(_16931_),
    .X(_17048_));
 sky130_fd_sc_hd__buf_1 _20141_ (.A(_17048_),
    .X(_17049_));
 sky130_fd_sc_hd__buf_1 _20142_ (.A(_17049_),
    .X(_17050_));
 sky130_fd_sc_hd__a21oi_2 _20143_ (.A1(_17041_),
    .A2(_17047_),
    .B1(_17050_),
    .Y(_04060_));
 sky130_fd_sc_hd__buf_1 _20144_ (.A(_16925_),
    .X(_17051_));
 sky130_fd_sc_hd__or4_2 _20145_ (.A(_17034_),
    .B(_17037_),
    .C(_17044_),
    .D(_17051_),
    .X(_17052_));
 sky130_fd_sc_hd__nand2_2 _20146_ (.A(_17045_),
    .B(_17038_),
    .Y(_17053_));
 sky130_fd_sc_hd__buf_1 _20147_ (.A(_17049_),
    .X(_17054_));
 sky130_fd_sc_hd__a21oi_2 _20148_ (.A1(_17052_),
    .A2(_17053_),
    .B1(_17054_),
    .Y(_04059_));
 sky130_fd_sc_hd__and2_2 _20149_ (.A(_16803_),
    .B(_16814_),
    .X(_17055_));
 sky130_vsdinv _20150_ (.A(_17055_),
    .Y(_17056_));
 sky130_fd_sc_hd__buf_1 _20151_ (.A(\cpu_state[4] ),
    .X(_17057_));
 sky130_fd_sc_hd__a21oi_2 _20152_ (.A1(_17028_),
    .A2(_17042_),
    .B1(_17057_),
    .Y(_17058_));
 sky130_vsdinv _20153_ (.A(is_lb_lh_lw_lbu_lhu),
    .Y(_17059_));
 sky130_fd_sc_hd__a21oi_2 _20154_ (.A1(_17004_),
    .A2(_17015_),
    .B1(_17059_),
    .Y(_17060_));
 sky130_vsdinv _20155_ (.A(is_sb_sh_sw),
    .Y(_17061_));
 sky130_fd_sc_hd__buf_1 _20156_ (.A(_17061_),
    .X(_17062_));
 sky130_vsdinv _20157_ (.A(_17014_),
    .Y(_17063_));
 sky130_fd_sc_hd__nor3_2 _20158_ (.A(_16997_),
    .B(_17063_),
    .C(_17002_),
    .Y(_17064_));
 sky130_fd_sc_hd__buf_1 _20159_ (.A(\cpu_state[3] ),
    .X(_17065_));
 sky130_fd_sc_hd__o211ai_2 _20160_ (.A1(_17062_),
    .A2(_17064_),
    .B1(_17065_),
    .C1(_17016_),
    .Y(_17066_));
 sky130_fd_sc_hd__o221a_2 _20161_ (.A1(_17024_),
    .A2(_17058_),
    .B1(_17021_),
    .B2(_17060_),
    .C1(_17066_),
    .X(_17067_));
 sky130_fd_sc_hd__buf_1 _20162_ (.A(_17055_),
    .X(_17068_));
 sky130_fd_sc_hd__buf_1 _20163_ (.A(_17068_),
    .X(_17069_));
 sky130_fd_sc_hd__nand3b_2 _20164_ (.A_N(_00356_),
    .B(_17067_),
    .C(_17069_),
    .Y(_17070_));
 sky130_fd_sc_hd__and2b_2 _20165_ (.A_N(alu_wait),
    .B(is_beq_bne_blt_bge_bltu_bgeu),
    .X(_17071_));
 sky130_vsdinv _20166_ (.A(_00343_),
    .Y(_17072_));
 sky130_fd_sc_hd__nor2_2 _20167_ (.A(_16821_),
    .B(\cpu_state[5] ),
    .Y(_17073_));
 sky130_fd_sc_hd__and4_2 _20168_ (.A(_17071_),
    .B(_16817_),
    .C(_17072_),
    .D(_17073_),
    .X(_17074_));
 sky130_vsdinv _20169_ (.A(\cpu_state[0] ),
    .Y(_17075_));
 sky130_fd_sc_hd__nand3_2 _20170_ (.A(_17028_),
    .B(_17043_),
    .C(_17075_),
    .Y(_17076_));
 sky130_vsdinv _20171_ (.A(_17076_),
    .Y(_17077_));
 sky130_fd_sc_hd__nand2_2 _20172_ (.A(_17074_),
    .B(_17077_),
    .Y(_17078_));
 sky130_fd_sc_hd__o311ai_2 _20173_ (.A1(_16858_),
    .A2(_17056_),
    .A3(_17067_),
    .B1(_17070_),
    .C1(_17078_),
    .Y(_04058_));
 sky130_fd_sc_hd__buf_1 _20174_ (.A(_16805_),
    .X(_17079_));
 sky130_fd_sc_hd__buf_1 _20175_ (.A(_17079_),
    .X(_17080_));
 sky130_fd_sc_hd__buf_1 _20176_ (.A(_17080_),
    .X(_17081_));
 sky130_fd_sc_hd__buf_1 _20177_ (.A(instr_jal),
    .X(_17082_));
 sky130_fd_sc_hd__buf_1 _20178_ (.A(_17082_),
    .X(_17083_));
 sky130_fd_sc_hd__buf_1 _20179_ (.A(_17083_),
    .X(_17084_));
 sky130_fd_sc_hd__nor2_2 _20180_ (.A(_17084_),
    .B(_16929_),
    .Y(_17085_));
 sky130_fd_sc_hd__buf_1 _20181_ (.A(instr_jalr),
    .X(_17086_));
 sky130_fd_sc_hd__o21ai_2 _20182_ (.A1(instr_retirq),
    .A2(_17086_),
    .B1(_17085_),
    .Y(_17087_));
 sky130_fd_sc_hd__o211a_2 _20183_ (.A1(_17081_),
    .A2(_17085_),
    .B1(_17069_),
    .C1(_17087_),
    .X(_04057_));
 sky130_fd_sc_hd__buf_1 _20184_ (.A(\irq_mask[31] ),
    .X(_17088_));
 sky130_fd_sc_hd__and2_2 _20185_ (.A(instr_maskirq),
    .B(_17019_),
    .X(_17089_));
 sky130_vsdinv _20186_ (.A(_17089_),
    .Y(_17090_));
 sky130_fd_sc_hd__buf_1 _20187_ (.A(_17090_),
    .X(_17091_));
 sky130_fd_sc_hd__buf_1 _20188_ (.A(_17091_),
    .X(_17092_));
 sky130_fd_sc_hd__buf_1 _20189_ (.A(_16842_),
    .X(_17093_));
 sky130_fd_sc_hd__buf_1 _20190_ (.A(_17093_),
    .X(_17094_));
 sky130_fd_sc_hd__nor3b_2 _20191_ (.A(_00362_),
    .B(_00360_),
    .C_N(_00368_),
    .Y(_17095_));
 sky130_fd_sc_hd__nor3b_2 _20192_ (.A(_00358_),
    .B(_00357_),
    .C_N(_17095_),
    .Y(_17096_));
 sky130_fd_sc_hd__buf_1 _20193_ (.A(_17096_),
    .X(_17097_));
 sky130_fd_sc_hd__buf_1 _20194_ (.A(_17097_),
    .X(_17098_));
 sky130_fd_sc_hd__nor2_2 _20195_ (.A(_01207_),
    .B(_17098_),
    .Y(\cpuregs_rs1[31] ));
 sky130_fd_sc_hd__buf_1 _20196_ (.A(_17089_),
    .X(_17099_));
 sky130_fd_sc_hd__nand2_2 _20197_ (.A(\cpuregs_rs1[31] ),
    .B(_17099_),
    .Y(_17100_));
 sky130_vsdinv _20198_ (.A(_17100_),
    .Y(_17101_));
 sky130_fd_sc_hd__a211o_2 _20199_ (.A1(_17088_),
    .A2(_17092_),
    .B1(_17094_),
    .C1(_17101_),
    .X(_04056_));
 sky130_fd_sc_hd__buf_1 _20200_ (.A(_17090_),
    .X(_17102_));
 sky130_fd_sc_hd__buf_1 _20201_ (.A(_17102_),
    .X(_17103_));
 sky130_fd_sc_hd__buf_1 _20202_ (.A(_17096_),
    .X(_17104_));
 sky130_fd_sc_hd__buf_1 _20203_ (.A(_17104_),
    .X(_17105_));
 sky130_fd_sc_hd__buf_1 _20204_ (.A(_17105_),
    .X(_17106_));
 sky130_fd_sc_hd__buf_1 _20205_ (.A(_17090_),
    .X(_17107_));
 sky130_fd_sc_hd__buf_1 _20206_ (.A(\irq_mask[30] ),
    .X(_17108_));
 sky130_fd_sc_hd__buf_1 _20207_ (.A(_17048_),
    .X(_17109_));
 sky130_fd_sc_hd__a21oi_2 _20208_ (.A1(_17107_),
    .A2(_17108_),
    .B1(_17109_),
    .Y(_17110_));
 sky130_fd_sc_hd__o31ai_2 _20209_ (.A1(_01180_),
    .A2(_17103_),
    .A3(_17106_),
    .B1(_17110_),
    .Y(_04055_));
 sky130_fd_sc_hd__buf_1 _20210_ (.A(_17096_),
    .X(_17111_));
 sky130_fd_sc_hd__buf_1 _20211_ (.A(_17111_),
    .X(_17112_));
 sky130_fd_sc_hd__nor2_2 _20212_ (.A(_01180_),
    .B(_17112_),
    .Y(\cpuregs_rs1[30] ));
 sky130_fd_sc_hd__buf_1 _20213_ (.A(\irq_mask[29] ),
    .X(_17113_));
 sky130_fd_sc_hd__nor2_2 _20214_ (.A(_01153_),
    .B(_17098_),
    .Y(\cpuregs_rs1[29] ));
 sky130_fd_sc_hd__nand2_2 _20215_ (.A(\cpuregs_rs1[29] ),
    .B(_17099_),
    .Y(_17114_));
 sky130_vsdinv _20216_ (.A(_17114_),
    .Y(_17115_));
 sky130_fd_sc_hd__a211o_2 _20217_ (.A1(_17113_),
    .A2(_17092_),
    .B1(_17094_),
    .C1(_17115_),
    .X(_04054_));
 sky130_fd_sc_hd__buf_1 _20218_ (.A(\irq_mask[28] ),
    .X(_17116_));
 sky130_fd_sc_hd__a21oi_2 _20219_ (.A1(_17107_),
    .A2(_17116_),
    .B1(_17109_),
    .Y(_17117_));
 sky130_fd_sc_hd__o31ai_2 _20220_ (.A1(_01126_),
    .A2(_17103_),
    .A3(_17106_),
    .B1(_17117_),
    .Y(_04053_));
 sky130_fd_sc_hd__nor2_2 _20221_ (.A(_01126_),
    .B(_17112_),
    .Y(\cpuregs_rs1[28] ));
 sky130_fd_sc_hd__buf_1 _20222_ (.A(_17099_),
    .X(_17118_));
 sky130_fd_sc_hd__buf_1 _20223_ (.A(_16816_),
    .X(_17119_));
 sky130_fd_sc_hd__buf_1 _20224_ (.A(_17119_),
    .X(_17120_));
 sky130_fd_sc_hd__buf_1 _20225_ (.A(_17120_),
    .X(_17121_));
 sky130_fd_sc_hd__buf_1 _20226_ (.A(_17111_),
    .X(_17122_));
 sky130_fd_sc_hd__nor2_2 _20227_ (.A(_01099_),
    .B(_17122_),
    .Y(\cpuregs_rs1[27] ));
 sky130_fd_sc_hd__buf_1 _20228_ (.A(_17089_),
    .X(_17123_));
 sky130_fd_sc_hd__buf_1 _20229_ (.A(_17123_),
    .X(_17124_));
 sky130_fd_sc_hd__nand2_2 _20230_ (.A(\cpuregs_rs1[27] ),
    .B(_17124_),
    .Y(_17125_));
 sky130_fd_sc_hd__o211ai_2 _20231_ (.A1(_16914_),
    .A2(_17118_),
    .B1(_17121_),
    .C1(_17125_),
    .Y(_04052_));
 sky130_fd_sc_hd__buf_1 _20232_ (.A(\irq_mask[26] ),
    .X(_17126_));
 sky130_fd_sc_hd__nor2_2 _20233_ (.A(_01072_),
    .B(_17098_),
    .Y(\cpuregs_rs1[26] ));
 sky130_fd_sc_hd__nand2_2 _20234_ (.A(\cpuregs_rs1[26] ),
    .B(_17099_),
    .Y(_17127_));
 sky130_vsdinv _20235_ (.A(_17127_),
    .Y(_17128_));
 sky130_fd_sc_hd__a211o_2 _20236_ (.A1(_17126_),
    .A2(_17092_),
    .B1(_17094_),
    .C1(_17128_),
    .X(_04051_));
 sky130_fd_sc_hd__buf_1 _20237_ (.A(\irq_mask[25] ),
    .X(_17129_));
 sky130_fd_sc_hd__nor2_2 _20238_ (.A(_01045_),
    .B(_17098_),
    .Y(\cpuregs_rs1[25] ));
 sky130_fd_sc_hd__buf_1 _20239_ (.A(_17089_),
    .X(_17130_));
 sky130_fd_sc_hd__buf_1 _20240_ (.A(_17130_),
    .X(_17131_));
 sky130_fd_sc_hd__nand2_2 _20241_ (.A(\cpuregs_rs1[25] ),
    .B(_17131_),
    .Y(_17132_));
 sky130_vsdinv _20242_ (.A(_17132_),
    .Y(_17133_));
 sky130_fd_sc_hd__a211o_2 _20243_ (.A1(_17129_),
    .A2(_17092_),
    .B1(_17094_),
    .C1(_17133_),
    .X(_04050_));
 sky130_fd_sc_hd__buf_1 _20244_ (.A(\irq_mask[24] ),
    .X(_17134_));
 sky130_fd_sc_hd__buf_1 _20245_ (.A(_17102_),
    .X(_17135_));
 sky130_fd_sc_hd__buf_1 _20246_ (.A(_17093_),
    .X(_17136_));
 sky130_fd_sc_hd__buf_1 _20247_ (.A(_17097_),
    .X(_17137_));
 sky130_fd_sc_hd__nor2_2 _20248_ (.A(_01018_),
    .B(_17137_),
    .Y(\cpuregs_rs1[24] ));
 sky130_fd_sc_hd__nand2_2 _20249_ (.A(\cpuregs_rs1[24] ),
    .B(_17131_),
    .Y(_17138_));
 sky130_vsdinv _20250_ (.A(_17138_),
    .Y(_17139_));
 sky130_fd_sc_hd__a211o_2 _20251_ (.A1(_17134_),
    .A2(_17135_),
    .B1(_17136_),
    .C1(_17139_),
    .X(_04049_));
 sky130_fd_sc_hd__nor2_2 _20252_ (.A(_00991_),
    .B(_17122_),
    .Y(\cpuregs_rs1[23] ));
 sky130_fd_sc_hd__nand2_2 _20253_ (.A(\cpuregs_rs1[23] ),
    .B(_17124_),
    .Y(_17140_));
 sky130_fd_sc_hd__o211ai_2 _20254_ (.A1(_16892_),
    .A2(_17118_),
    .B1(_17121_),
    .C1(_17140_),
    .Y(_04048_));
 sky130_fd_sc_hd__buf_1 _20255_ (.A(_17091_),
    .X(_17141_));
 sky130_fd_sc_hd__buf_1 _20256_ (.A(_17090_),
    .X(_17142_));
 sky130_fd_sc_hd__buf_1 _20257_ (.A(\irq_mask[22] ),
    .X(_17143_));
 sky130_fd_sc_hd__a21oi_2 _20258_ (.A1(_17142_),
    .A2(_17143_),
    .B1(_17109_),
    .Y(_17144_));
 sky130_fd_sc_hd__o31ai_2 _20259_ (.A1(_00964_),
    .A2(_17141_),
    .A3(_17106_),
    .B1(_17144_),
    .Y(_04047_));
 sky130_fd_sc_hd__nor2_2 _20260_ (.A(_00964_),
    .B(_17112_),
    .Y(\cpuregs_rs1[22] ));
 sky130_fd_sc_hd__buf_1 _20261_ (.A(_17105_),
    .X(_17145_));
 sky130_fd_sc_hd__buf_1 _20262_ (.A(\irq_mask[21] ),
    .X(_17146_));
 sky130_fd_sc_hd__buf_1 _20263_ (.A(_16841_),
    .X(_17147_));
 sky130_fd_sc_hd__buf_1 _20264_ (.A(_17147_),
    .X(_17148_));
 sky130_fd_sc_hd__buf_1 _20265_ (.A(_17148_),
    .X(_17149_));
 sky130_fd_sc_hd__a21oi_2 _20266_ (.A1(_17142_),
    .A2(_17146_),
    .B1(_17149_),
    .Y(_17150_));
 sky130_fd_sc_hd__o31ai_2 _20267_ (.A1(_00937_),
    .A2(_17141_),
    .A3(_17145_),
    .B1(_17150_),
    .Y(_04046_));
 sky130_fd_sc_hd__nor2_2 _20268_ (.A(_00937_),
    .B(_17112_),
    .Y(\cpuregs_rs1[21] ));
 sky130_fd_sc_hd__buf_1 _20269_ (.A(\irq_mask[20] ),
    .X(_17151_));
 sky130_fd_sc_hd__nor2_2 _20270_ (.A(_00910_),
    .B(_17137_),
    .Y(\cpuregs_rs1[20] ));
 sky130_fd_sc_hd__nand2_2 _20271_ (.A(\cpuregs_rs1[20] ),
    .B(_17131_),
    .Y(_17152_));
 sky130_vsdinv _20272_ (.A(_17152_),
    .Y(_17153_));
 sky130_fd_sc_hd__a211o_2 _20273_ (.A1(_17151_),
    .A2(_17135_),
    .B1(_17136_),
    .C1(_17153_),
    .X(_04045_));
 sky130_fd_sc_hd__buf_1 _20274_ (.A(\irq_mask[19] ),
    .X(_17154_));
 sky130_fd_sc_hd__a21oi_2 _20275_ (.A1(_17142_),
    .A2(_17154_),
    .B1(_17149_),
    .Y(_17155_));
 sky130_fd_sc_hd__o31ai_2 _20276_ (.A1(_00883_),
    .A2(_17141_),
    .A3(_17145_),
    .B1(_17155_),
    .Y(_04044_));
 sky130_fd_sc_hd__buf_1 _20277_ (.A(_17111_),
    .X(_17156_));
 sky130_fd_sc_hd__nor2_2 _20278_ (.A(_00883_),
    .B(_17156_),
    .Y(\cpuregs_rs1[19] ));
 sky130_fd_sc_hd__buf_1 _20279_ (.A(\irq_mask[18] ),
    .X(_17157_));
 sky130_fd_sc_hd__a21oi_2 _20280_ (.A1(_17142_),
    .A2(_17157_),
    .B1(_17149_),
    .Y(_17158_));
 sky130_fd_sc_hd__o31ai_2 _20281_ (.A1(_00856_),
    .A2(_17141_),
    .A3(_17145_),
    .B1(_17158_),
    .Y(_04043_));
 sky130_fd_sc_hd__nor2_2 _20282_ (.A(_00856_),
    .B(_17156_),
    .Y(\cpuregs_rs1[18] ));
 sky130_fd_sc_hd__buf_1 _20283_ (.A(\irq_mask[17] ),
    .X(_17159_));
 sky130_fd_sc_hd__nor2_2 _20284_ (.A(_00829_),
    .B(_17137_),
    .Y(\cpuregs_rs1[17] ));
 sky130_fd_sc_hd__nand2_2 _20285_ (.A(\cpuregs_rs1[17] ),
    .B(_17131_),
    .Y(_17160_));
 sky130_vsdinv _20286_ (.A(_17160_),
    .Y(_17161_));
 sky130_fd_sc_hd__a211o_2 _20287_ (.A1(_17159_),
    .A2(_17135_),
    .B1(_17136_),
    .C1(_17161_),
    .X(_04042_));
 sky130_fd_sc_hd__buf_1 _20288_ (.A(\irq_mask[16] ),
    .X(_17162_));
 sky130_fd_sc_hd__a21oi_2 _20289_ (.A1(_17091_),
    .A2(_17162_),
    .B1(_17149_),
    .Y(_17163_));
 sky130_fd_sc_hd__o31ai_2 _20290_ (.A1(_00802_),
    .A2(_17107_),
    .A3(_17145_),
    .B1(_17163_),
    .Y(_04041_));
 sky130_fd_sc_hd__nor2_2 _20291_ (.A(_00802_),
    .B(_17156_),
    .Y(\cpuregs_rs1[16] ));
 sky130_fd_sc_hd__nor2_2 _20292_ (.A(_00775_),
    .B(_17122_),
    .Y(\cpuregs_rs1[15] ));
 sky130_fd_sc_hd__buf_1 _20293_ (.A(_17130_),
    .X(_17164_));
 sky130_fd_sc_hd__nand2_2 _20294_ (.A(\cpuregs_rs1[15] ),
    .B(_17164_),
    .Y(_17165_));
 sky130_fd_sc_hd__o211ai_2 _20295_ (.A1(_16919_),
    .A2(_17118_),
    .B1(_17121_),
    .C1(_17165_),
    .Y(_04040_));
 sky130_fd_sc_hd__buf_1 _20296_ (.A(\irq_mask[14] ),
    .X(_17166_));
 sky130_fd_sc_hd__nor2_2 _20297_ (.A(_00748_),
    .B(_17137_),
    .Y(\cpuregs_rs1[14] ));
 sky130_fd_sc_hd__buf_1 _20298_ (.A(_17130_),
    .X(_17167_));
 sky130_fd_sc_hd__nand2_2 _20299_ (.A(\cpuregs_rs1[14] ),
    .B(_17167_),
    .Y(_17168_));
 sky130_vsdinv _20300_ (.A(_17168_),
    .Y(_17169_));
 sky130_fd_sc_hd__a211o_2 _20301_ (.A1(_17166_),
    .A2(_17135_),
    .B1(_17136_),
    .C1(_17169_),
    .X(_04039_));
 sky130_fd_sc_hd__buf_1 _20302_ (.A(\irq_mask[13] ),
    .X(_17170_));
 sky130_fd_sc_hd__buf_1 _20303_ (.A(_17102_),
    .X(_17171_));
 sky130_fd_sc_hd__buf_1 _20304_ (.A(_17093_),
    .X(_17172_));
 sky130_fd_sc_hd__buf_1 _20305_ (.A(_17097_),
    .X(_17173_));
 sky130_fd_sc_hd__nor2_2 _20306_ (.A(_00721_),
    .B(_17173_),
    .Y(\cpuregs_rs1[13] ));
 sky130_fd_sc_hd__nand2_2 _20307_ (.A(\cpuregs_rs1[13] ),
    .B(_17167_),
    .Y(_17174_));
 sky130_vsdinv _20308_ (.A(_17174_),
    .Y(_17175_));
 sky130_fd_sc_hd__a211o_2 _20309_ (.A1(_17170_),
    .A2(_17171_),
    .B1(_17172_),
    .C1(_17175_),
    .X(_04038_));
 sky130_fd_sc_hd__buf_1 _20310_ (.A(\irq_mask[12] ),
    .X(_17176_));
 sky130_fd_sc_hd__nor2_2 _20311_ (.A(_00694_),
    .B(_17173_),
    .Y(\cpuregs_rs1[12] ));
 sky130_fd_sc_hd__nand2_2 _20312_ (.A(\cpuregs_rs1[12] ),
    .B(_17167_),
    .Y(_17177_));
 sky130_vsdinv _20313_ (.A(_17177_),
    .Y(_17178_));
 sky130_fd_sc_hd__a211o_2 _20314_ (.A1(_17176_),
    .A2(_17171_),
    .B1(_17172_),
    .C1(_17178_),
    .X(_04037_));
 sky130_fd_sc_hd__nor2_2 _20315_ (.A(_00667_),
    .B(_17122_),
    .Y(\cpuregs_rs1[11] ));
 sky130_fd_sc_hd__nand2_2 _20316_ (.A(\cpuregs_rs1[11] ),
    .B(_17164_),
    .Y(_17179_));
 sky130_fd_sc_hd__o211ai_2 _20317_ (.A1(_16882_),
    .A2(_17118_),
    .B1(_17121_),
    .C1(_17179_),
    .Y(_04036_));
 sky130_fd_sc_hd__buf_1 _20318_ (.A(\irq_mask[10] ),
    .X(_17180_));
 sky130_fd_sc_hd__nor2_2 _20319_ (.A(_00640_),
    .B(_17173_),
    .Y(\cpuregs_rs1[10] ));
 sky130_fd_sc_hd__nand2_2 _20320_ (.A(\cpuregs_rs1[10] ),
    .B(_17167_),
    .Y(_17181_));
 sky130_vsdinv _20321_ (.A(_17181_),
    .Y(_17182_));
 sky130_fd_sc_hd__a211o_2 _20322_ (.A1(_17180_),
    .A2(_17171_),
    .B1(_17172_),
    .C1(_17182_),
    .X(_04035_));
 sky130_fd_sc_hd__buf_1 _20323_ (.A(\irq_mask[9] ),
    .X(_17183_));
 sky130_fd_sc_hd__nor2_2 _20324_ (.A(_00613_),
    .B(_17173_),
    .Y(\cpuregs_rs1[9] ));
 sky130_fd_sc_hd__buf_1 _20325_ (.A(_17130_),
    .X(_17184_));
 sky130_fd_sc_hd__nand2_2 _20326_ (.A(\cpuregs_rs1[9] ),
    .B(_17184_),
    .Y(_17185_));
 sky130_vsdinv _20327_ (.A(_17185_),
    .Y(_17186_));
 sky130_fd_sc_hd__a211o_2 _20328_ (.A1(_17183_),
    .A2(_17171_),
    .B1(_17172_),
    .C1(_17186_),
    .X(_04034_));
 sky130_fd_sc_hd__buf_1 _20329_ (.A(\irq_mask[8] ),
    .X(_17187_));
 sky130_fd_sc_hd__buf_1 _20330_ (.A(_17102_),
    .X(_17188_));
 sky130_fd_sc_hd__buf_1 _20331_ (.A(_16842_),
    .X(_17189_));
 sky130_fd_sc_hd__buf_1 _20332_ (.A(_17189_),
    .X(_17190_));
 sky130_fd_sc_hd__buf_1 _20333_ (.A(_17097_),
    .X(_17191_));
 sky130_fd_sc_hd__nor2_2 _20334_ (.A(_00586_),
    .B(_17191_),
    .Y(\cpuregs_rs1[8] ));
 sky130_fd_sc_hd__nand2_2 _20335_ (.A(\cpuregs_rs1[8] ),
    .B(_17184_),
    .Y(_17192_));
 sky130_vsdinv _20336_ (.A(_17192_),
    .Y(_17193_));
 sky130_fd_sc_hd__a211o_2 _20337_ (.A1(_17187_),
    .A2(_17188_),
    .B1(_17190_),
    .C1(_17193_),
    .X(_04033_));
 sky130_fd_sc_hd__buf_1 _20338_ (.A(_16831_),
    .X(_17194_));
 sky130_fd_sc_hd__nor2_2 _20339_ (.A(_00559_),
    .B(_17104_),
    .Y(\cpuregs_rs1[7] ));
 sky130_fd_sc_hd__nand2_2 _20340_ (.A(\cpuregs_rs1[7] ),
    .B(_17164_),
    .Y(_17195_));
 sky130_fd_sc_hd__o211ai_2 _20341_ (.A1(_16897_),
    .A2(_17124_),
    .B1(_17194_),
    .C1(_17195_),
    .Y(_04032_));
 sky130_fd_sc_hd__buf_1 _20342_ (.A(\irq_mask[6] ),
    .X(_17196_));
 sky130_fd_sc_hd__buf_1 _20343_ (.A(_17148_),
    .X(_17197_));
 sky130_fd_sc_hd__a21oi_2 _20344_ (.A1(_17091_),
    .A2(_17196_),
    .B1(_17197_),
    .Y(_17198_));
 sky130_fd_sc_hd__o31ai_2 _20345_ (.A1(_00532_),
    .A2(_17107_),
    .A3(_17105_),
    .B1(_17198_),
    .Y(_04031_));
 sky130_fd_sc_hd__nor2_2 _20346_ (.A(_00532_),
    .B(_17156_),
    .Y(\cpuregs_rs1[6] ));
 sky130_fd_sc_hd__buf_1 _20347_ (.A(\irq_mask[5] ),
    .X(_17199_));
 sky130_fd_sc_hd__nor2_2 _20348_ (.A(_00505_),
    .B(_17191_),
    .Y(\cpuregs_rs1[5] ));
 sky130_fd_sc_hd__nand2_2 _20349_ (.A(\cpuregs_rs1[5] ),
    .B(_17184_),
    .Y(_17200_));
 sky130_vsdinv _20350_ (.A(_17200_),
    .Y(_17201_));
 sky130_fd_sc_hd__a211o_2 _20351_ (.A1(_17199_),
    .A2(_17188_),
    .B1(_17190_),
    .C1(_17201_),
    .X(_04030_));
 sky130_fd_sc_hd__buf_1 _20352_ (.A(\irq_mask[4] ),
    .X(_17202_));
 sky130_fd_sc_hd__nor2_2 _20353_ (.A(_00478_),
    .B(_17191_),
    .Y(\cpuregs_rs1[4] ));
 sky130_fd_sc_hd__nand2_2 _20354_ (.A(\cpuregs_rs1[4] ),
    .B(_17184_),
    .Y(_17203_));
 sky130_vsdinv _20355_ (.A(_17203_),
    .Y(_17204_));
 sky130_fd_sc_hd__a211o_2 _20356_ (.A1(_17202_),
    .A2(_17188_),
    .B1(_17190_),
    .C1(_17204_),
    .X(_04029_));
 sky130_fd_sc_hd__buf_1 _20357_ (.A(\irq_mask[3] ),
    .X(_17205_));
 sky130_fd_sc_hd__nor2_2 _20358_ (.A(_00451_),
    .B(_17191_),
    .Y(\cpuregs_rs1[3] ));
 sky130_fd_sc_hd__nand2_2 _20359_ (.A(\cpuregs_rs1[3] ),
    .B(_17123_),
    .Y(_17206_));
 sky130_vsdinv _20360_ (.A(_17206_),
    .Y(_17207_));
 sky130_fd_sc_hd__a211o_2 _20361_ (.A1(_17205_),
    .A2(_17188_),
    .B1(_17190_),
    .C1(_17207_),
    .X(_04028_));
 sky130_fd_sc_hd__nor2_2 _20362_ (.A(_00424_),
    .B(_17104_),
    .Y(\cpuregs_rs1[2] ));
 sky130_fd_sc_hd__nand2_2 _20363_ (.A(\cpuregs_rs1[2] ),
    .B(_17164_),
    .Y(_17208_));
 sky130_fd_sc_hd__o211ai_2 _20364_ (.A1(_16887_),
    .A2(_17124_),
    .B1(_17194_),
    .C1(_17208_),
    .Y(_04027_));
 sky130_fd_sc_hd__buf_1 _20365_ (.A(\irq_mask[1] ),
    .X(_17209_));
 sky130_fd_sc_hd__buf_1 _20366_ (.A(_17209_),
    .X(_17210_));
 sky130_fd_sc_hd__buf_1 _20367_ (.A(_17189_),
    .X(_17211_));
 sky130_fd_sc_hd__nor2_2 _20368_ (.A(_00397_),
    .B(_17111_),
    .Y(\cpuregs_rs1[1] ));
 sky130_fd_sc_hd__nand2_2 _20369_ (.A(\cpuregs_rs1[1] ),
    .B(_17123_),
    .Y(_17212_));
 sky130_vsdinv _20370_ (.A(_17212_),
    .Y(_17213_));
 sky130_fd_sc_hd__a211o_2 _20371_ (.A1(_17210_),
    .A2(_17103_),
    .B1(_17211_),
    .C1(_17213_),
    .X(_04026_));
 sky130_fd_sc_hd__buf_1 _20372_ (.A(\irq_mask[0] ),
    .X(_17214_));
 sky130_fd_sc_hd__nand3b_2 _20373_ (.A_N(_17104_),
    .B(_00370_),
    .C(_17123_),
    .Y(_17215_));
 sky130_vsdinv _20374_ (.A(_17215_),
    .Y(_17216_));
 sky130_fd_sc_hd__a211o_2 _20375_ (.A1(_17214_),
    .A2(_17103_),
    .B1(_17211_),
    .C1(_17216_),
    .X(_04025_));
 sky130_fd_sc_hd__nor2b_2 _20376_ (.A(_17106_),
    .B_N(_00370_),
    .Y(\cpuregs_rs1[0] ));
 sky130_fd_sc_hd__buf_1 _20377_ (.A(_16848_),
    .X(_17217_));
 sky130_fd_sc_hd__buf_1 _20378_ (.A(_17217_),
    .X(_17218_));
 sky130_fd_sc_hd__o21ba_2 _20379_ (.A1(_16845_),
    .A2(_17080_),
    .B1_N(_17218_),
    .X(_17219_));
 sky130_vsdinv _20380_ (.A(trap),
    .Y(_17220_));
 sky130_fd_sc_hd__buf_1 _20381_ (.A(_16814_),
    .X(_17221_));
 sky130_fd_sc_hd__nor3b_2 _20382_ (.A(\mem_state[1] ),
    .B(_16797_),
    .C_N(_17221_),
    .Y(_17222_));
 sky130_fd_sc_hd__nand3_2 _20383_ (.A(_16850_),
    .B(_17220_),
    .C(_17222_),
    .Y(_17223_));
 sky130_fd_sc_hd__buf_1 _20384_ (.A(_17223_),
    .X(_17224_));
 sky130_fd_sc_hd__buf_1 _20385_ (.A(_17224_),
    .X(_17225_));
 sky130_fd_sc_hd__mux2_2 _20386_ (.A0(_17219_),
    .A1(mem_instr),
    .S(_17225_),
    .X(_04024_));
 sky130_fd_sc_hd__buf_1 _20387_ (.A(_16981_),
    .X(_17226_));
 sky130_fd_sc_hd__buf_1 _20388_ (.A(_16818_),
    .X(_17227_));
 sky130_fd_sc_hd__buf_1 _20389_ (.A(_00327_),
    .X(_17228_));
 sky130_fd_sc_hd__buf_1 _20390_ (.A(_00328_),
    .X(_17229_));
 sky130_fd_sc_hd__buf_1 _20391_ (.A(_00329_),
    .X(_17230_));
 sky130_fd_sc_hd__nand3b_2 _20392_ (.A_N(_17229_),
    .B(_17230_),
    .C(_00330_),
    .Y(_17231_));
 sky130_fd_sc_hd__o31ai_2 _20393_ (.A1(_17228_),
    .A2(_16866_),
    .A3(_17231_),
    .B1(_16872_),
    .Y(_17232_));
 sky130_fd_sc_hd__o211a_2 _20394_ (.A1(_17226_),
    .A2(_16863_),
    .B1(_17227_),
    .C1(_17232_),
    .X(_04023_));
 sky130_vsdinv _20395_ (.A(_16860_),
    .Y(_17233_));
 sky130_fd_sc_hd__buf_1 _20396_ (.A(_17233_),
    .X(_17234_));
 sky130_fd_sc_hd__and2_2 _20397_ (.A(_16861_),
    .B(\mem_rdata_latched[18] ),
    .X(_17235_));
 sky130_vsdinv _20398_ (.A(_16871_),
    .Y(_17236_));
 sky130_fd_sc_hd__a22o_2 _20399_ (.A1(\decoded_rs1[3] ),
    .A2(_17234_),
    .B1(_17235_),
    .B2(_17236_),
    .X(_04022_));
 sky130_fd_sc_hd__buf_1 _20400_ (.A(_17233_),
    .X(_17237_));
 sky130_fd_sc_hd__and2_2 _20401_ (.A(_16861_),
    .B(\mem_rdata_latched[17] ),
    .X(_17238_));
 sky130_fd_sc_hd__a22o_2 _20402_ (.A1(\decoded_rs1[2] ),
    .A2(_17237_),
    .B1(_17238_),
    .B2(_17236_),
    .X(_04021_));
 sky130_fd_sc_hd__and2_2 _20403_ (.A(_16862_),
    .B(\mem_rdata_latched[16] ),
    .X(_17239_));
 sky130_fd_sc_hd__a22o_2 _20404_ (.A1(\decoded_rs1[1] ),
    .A2(_17237_),
    .B1(_17239_),
    .B2(_17236_),
    .X(_04020_));
 sky130_fd_sc_hd__and2_2 _20405_ (.A(_16862_),
    .B(\mem_rdata_latched[15] ),
    .X(_17240_));
 sky130_fd_sc_hd__a22o_2 _20406_ (.A1(\decoded_rs1[0] ),
    .A2(_17237_),
    .B1(_17240_),
    .B2(_17236_),
    .X(_04019_));
 sky130_fd_sc_hd__buf_1 _20407_ (.A(\mem_rdata_q[14] ),
    .X(_17241_));
 sky130_fd_sc_hd__buf_1 _20408_ (.A(_17241_),
    .X(_17242_));
 sky130_fd_sc_hd__buf_1 _20409_ (.A(\mem_rdata_q[13] ),
    .X(_17243_));
 sky130_fd_sc_hd__buf_1 _20410_ (.A(_17243_),
    .X(_17244_));
 sky130_fd_sc_hd__buf_1 _20411_ (.A(\mem_rdata_q[12] ),
    .X(_17245_));
 sky130_fd_sc_hd__nand3_2 _20412_ (.A(_17242_),
    .B(_17244_),
    .C(_17245_),
    .Y(_17246_));
 sky130_vsdinv _20413_ (.A(\mem_rdata_q[31] ),
    .Y(_17247_));
 sky130_fd_sc_hd__buf_1 _20414_ (.A(_17247_),
    .X(_17248_));
 sky130_vsdinv _20415_ (.A(\mem_rdata_q[30] ),
    .Y(_17249_));
 sky130_vsdinv _20416_ (.A(\mem_rdata_q[29] ),
    .Y(_17250_));
 sky130_fd_sc_hd__nand3_2 _20417_ (.A(_17248_),
    .B(_17249_),
    .C(_17250_),
    .Y(_17251_));
 sky130_fd_sc_hd__nor2_2 _20418_ (.A(\mem_rdata_q[28] ),
    .B(\mem_rdata_q[26] ),
    .Y(_17252_));
 sky130_fd_sc_hd__nor2_2 _20419_ (.A(\mem_rdata_q[27] ),
    .B(\mem_rdata_q[25] ),
    .Y(_17253_));
 sky130_fd_sc_hd__nand2_2 _20420_ (.A(_17252_),
    .B(_17253_),
    .Y(_17254_));
 sky130_fd_sc_hd__buf_1 _20421_ (.A(_16927_),
    .X(_17255_));
 sky130_fd_sc_hd__and2b_2 _20422_ (.A_N(decoder_pseudo_trigger),
    .B(_17255_),
    .X(_17256_));
 sky130_vsdinv _20423_ (.A(_17256_),
    .Y(_17257_));
 sky130_fd_sc_hd__buf_1 _20424_ (.A(_17257_),
    .X(_17258_));
 sky130_fd_sc_hd__nor3_2 _20425_ (.A(_17251_),
    .B(_17254_),
    .C(_17258_),
    .Y(_17259_));
 sky130_fd_sc_hd__buf_1 _20426_ (.A(_17259_),
    .X(_17260_));
 sky130_fd_sc_hd__buf_1 _20427_ (.A(is_alu_reg_reg),
    .X(_17261_));
 sky130_fd_sc_hd__nand3b_2 _20428_ (.A_N(_17246_),
    .B(_17260_),
    .C(_17261_),
    .Y(_17262_));
 sky130_fd_sc_hd__buf_1 _20429_ (.A(decoder_pseudo_trigger),
    .X(_17263_));
 sky130_fd_sc_hd__buf_1 _20430_ (.A(_17263_),
    .X(_17264_));
 sky130_fd_sc_hd__buf_1 _20431_ (.A(_17264_),
    .X(_17265_));
 sky130_vsdinv _20432_ (.A(_16927_),
    .Y(_17266_));
 sky130_fd_sc_hd__buf_1 _20433_ (.A(_17266_),
    .X(_17267_));
 sky130_fd_sc_hd__buf_1 _20434_ (.A(_17267_),
    .X(_17268_));
 sky130_fd_sc_hd__buf_1 _20435_ (.A(instr_and),
    .X(_17269_));
 sky130_fd_sc_hd__buf_1 _20436_ (.A(_17269_),
    .X(_17270_));
 sky130_fd_sc_hd__o21ai_2 _20437_ (.A1(_17265_),
    .A2(_17268_),
    .B1(_17270_),
    .Y(_17271_));
 sky130_fd_sc_hd__a21oi_2 _20438_ (.A1(_17262_),
    .A2(_17271_),
    .B1(_17054_),
    .Y(_04018_));
 sky130_fd_sc_hd__buf_1 _20439_ (.A(\mem_rdata_q[14] ),
    .X(_17272_));
 sky130_fd_sc_hd__nand3b_2 _20440_ (.A_N(_17245_),
    .B(_17272_),
    .C(_17244_),
    .Y(_17273_));
 sky130_fd_sc_hd__nand3b_2 _20441_ (.A_N(_17273_),
    .B(_17260_),
    .C(_17261_),
    .Y(_17274_));
 sky130_fd_sc_hd__buf_1 _20442_ (.A(instr_or),
    .X(_17275_));
 sky130_fd_sc_hd__buf_1 _20443_ (.A(_17275_),
    .X(_17276_));
 sky130_fd_sc_hd__o21ai_2 _20444_ (.A1(_17265_),
    .A2(_17268_),
    .B1(_17276_),
    .Y(_17277_));
 sky130_fd_sc_hd__a21oi_2 _20445_ (.A1(_17274_),
    .A2(_17277_),
    .B1(_17054_),
    .Y(_04017_));
 sky130_fd_sc_hd__and4_2 _20446_ (.A(_17252_),
    .B(_17253_),
    .C(_17248_),
    .D(\mem_rdata_q[30] ),
    .X(_17278_));
 sky130_vsdinv _20447_ (.A(is_alu_reg_reg),
    .Y(_17279_));
 sky130_fd_sc_hd__nand3b_2 _20448_ (.A_N(_17243_),
    .B(_17241_),
    .C(_17245_),
    .Y(_17280_));
 sky130_fd_sc_hd__nor2_2 _20449_ (.A(_17279_),
    .B(_17280_),
    .Y(_17281_));
 sky130_fd_sc_hd__buf_1 _20450_ (.A(\mem_rdata_q[29] ),
    .X(_17282_));
 sky130_fd_sc_hd__buf_1 _20451_ (.A(decoder_pseudo_trigger),
    .X(_17283_));
 sky130_fd_sc_hd__buf_1 _20452_ (.A(_17255_),
    .X(_17284_));
 sky130_fd_sc_hd__nor3b_2 _20453_ (.A(_17282_),
    .B(_17283_),
    .C_N(_17284_),
    .Y(_17285_));
 sky130_fd_sc_hd__nand3_2 _20454_ (.A(_17278_),
    .B(_17281_),
    .C(_17285_),
    .Y(_17286_));
 sky130_fd_sc_hd__o21ai_2 _20455_ (.A1(_17265_),
    .A2(_17268_),
    .B1(instr_sra),
    .Y(_17287_));
 sky130_fd_sc_hd__a21oi_2 _20456_ (.A1(_17286_),
    .A2(_17287_),
    .B1(_17054_),
    .Y(_04016_));
 sky130_fd_sc_hd__nor2_2 _20457_ (.A(_17251_),
    .B(_17254_),
    .Y(_17288_));
 sky130_fd_sc_hd__buf_1 _20458_ (.A(_17256_),
    .X(_17289_));
 sky130_fd_sc_hd__buf_1 _20459_ (.A(_17289_),
    .X(_17290_));
 sky130_fd_sc_hd__buf_1 _20460_ (.A(_17290_),
    .X(_17291_));
 sky130_fd_sc_hd__nand3_2 _20461_ (.A(_17288_),
    .B(_17291_),
    .C(_17281_),
    .Y(_17292_));
 sky130_fd_sc_hd__buf_1 _20462_ (.A(_17263_),
    .X(_17293_));
 sky130_fd_sc_hd__buf_1 _20463_ (.A(_17293_),
    .X(_17294_));
 sky130_fd_sc_hd__o21ai_2 _20464_ (.A1(_17294_),
    .A2(_17268_),
    .B1(instr_srl),
    .Y(_17295_));
 sky130_fd_sc_hd__buf_1 _20465_ (.A(_17049_),
    .X(_17296_));
 sky130_fd_sc_hd__a21oi_2 _20466_ (.A1(_17292_),
    .A2(_17295_),
    .B1(_17296_),
    .Y(_04015_));
 sky130_fd_sc_hd__buf_1 _20467_ (.A(_17259_),
    .X(_17297_));
 sky130_fd_sc_hd__buf_1 _20468_ (.A(_17261_),
    .X(_17298_));
 sky130_fd_sc_hd__nor3b_2 _20469_ (.A(_17244_),
    .B(_17245_),
    .C_N(_17242_),
    .Y(_17299_));
 sky130_fd_sc_hd__nand3_2 _20470_ (.A(_17297_),
    .B(_17298_),
    .C(_17299_),
    .Y(_17300_));
 sky130_fd_sc_hd__buf_1 _20471_ (.A(_17266_),
    .X(_17301_));
 sky130_fd_sc_hd__buf_1 _20472_ (.A(_17301_),
    .X(_17302_));
 sky130_fd_sc_hd__buf_1 _20473_ (.A(instr_xor),
    .X(_17303_));
 sky130_fd_sc_hd__o21ai_2 _20474_ (.A1(_17294_),
    .A2(_17302_),
    .B1(_17303_),
    .Y(_17304_));
 sky130_fd_sc_hd__a21oi_2 _20475_ (.A1(_17300_),
    .A2(_17304_),
    .B1(_17296_),
    .Y(_04014_));
 sky130_fd_sc_hd__buf_1 _20476_ (.A(\mem_rdata_q[12] ),
    .X(_17305_));
 sky130_fd_sc_hd__nand2_2 _20477_ (.A(_17243_),
    .B(_17305_),
    .Y(_17306_));
 sky130_fd_sc_hd__nor2_2 _20478_ (.A(_17272_),
    .B(_17306_),
    .Y(_17307_));
 sky130_fd_sc_hd__nand3_2 _20479_ (.A(_17297_),
    .B(_17298_),
    .C(_17307_),
    .Y(_17308_));
 sky130_fd_sc_hd__o21ai_2 _20480_ (.A1(_17294_),
    .A2(_17302_),
    .B1(instr_sltu),
    .Y(_17309_));
 sky130_fd_sc_hd__a21oi_2 _20481_ (.A1(_17308_),
    .A2(_17309_),
    .B1(_17296_),
    .Y(_04013_));
 sky130_fd_sc_hd__nor3b_2 _20482_ (.A(\mem_rdata_q[14] ),
    .B(\mem_rdata_q[12] ),
    .C_N(\mem_rdata_q[13] ),
    .Y(_17310_));
 sky130_fd_sc_hd__nand3_2 _20483_ (.A(_17260_),
    .B(_17298_),
    .C(_17310_),
    .Y(_17311_));
 sky130_fd_sc_hd__o21ai_2 _20484_ (.A1(_17294_),
    .A2(_17302_),
    .B1(instr_slt),
    .Y(_17312_));
 sky130_fd_sc_hd__a21oi_2 _20485_ (.A1(_17311_),
    .A2(_17312_),
    .B1(_17296_),
    .Y(_04012_));
 sky130_fd_sc_hd__nor3b_2 _20486_ (.A(_17272_),
    .B(_17244_),
    .C_N(_17305_),
    .Y(_17313_));
 sky130_fd_sc_hd__nand3_2 _20487_ (.A(_17260_),
    .B(_17298_),
    .C(_17313_),
    .Y(_17314_));
 sky130_fd_sc_hd__buf_1 _20488_ (.A(_17293_),
    .X(_17315_));
 sky130_fd_sc_hd__buf_1 _20489_ (.A(instr_sll),
    .X(_17316_));
 sky130_fd_sc_hd__o21ai_2 _20490_ (.A1(_17315_),
    .A2(_17302_),
    .B1(_17316_),
    .Y(_17317_));
 sky130_fd_sc_hd__buf_1 _20491_ (.A(_17048_),
    .X(_17318_));
 sky130_fd_sc_hd__buf_1 _20492_ (.A(_17318_),
    .X(_17319_));
 sky130_fd_sc_hd__a21oi_2 _20493_ (.A1(_17314_),
    .A2(_17317_),
    .B1(_17319_),
    .Y(_04011_));
 sky130_fd_sc_hd__buf_1 _20494_ (.A(_17293_),
    .X(_17320_));
 sky130_fd_sc_hd__o21a_2 _20495_ (.A1(_17320_),
    .A2(_17267_),
    .B1(instr_sub),
    .X(_17321_));
 sky130_fd_sc_hd__or3_2 _20496_ (.A(_17241_),
    .B(\mem_rdata_q[13] ),
    .C(_17305_),
    .X(_17322_));
 sky130_fd_sc_hd__and4b_2 _20497_ (.A_N(_17322_),
    .B(_17278_),
    .C(is_alu_reg_reg),
    .D(_17285_),
    .X(_17323_));
 sky130_fd_sc_hd__buf_1 _20498_ (.A(_16854_),
    .X(_17324_));
 sky130_fd_sc_hd__buf_1 _20499_ (.A(_17324_),
    .X(_17325_));
 sky130_fd_sc_hd__buf_1 _20500_ (.A(_17325_),
    .X(_17326_));
 sky130_fd_sc_hd__o21a_2 _20501_ (.A1(_17321_),
    .A2(_17323_),
    .B1(_17326_),
    .X(_04010_));
 sky130_fd_sc_hd__nand3b_2 _20502_ (.A_N(_17322_),
    .B(_17259_),
    .C(_17261_),
    .Y(_17327_));
 sky130_fd_sc_hd__buf_1 _20503_ (.A(_17301_),
    .X(_17328_));
 sky130_fd_sc_hd__o21ai_2 _20504_ (.A1(_17315_),
    .A2(_17328_),
    .B1(instr_add),
    .Y(_17329_));
 sky130_fd_sc_hd__a21oi_2 _20505_ (.A1(_17327_),
    .A2(_17329_),
    .B1(_17319_),
    .Y(_04009_));
 sky130_fd_sc_hd__buf_1 _20506_ (.A(_17256_),
    .X(_17330_));
 sky130_fd_sc_hd__buf_1 _20507_ (.A(_17330_),
    .X(_17331_));
 sky130_fd_sc_hd__buf_1 _20508_ (.A(is_alu_reg_imm),
    .X(_17332_));
 sky130_fd_sc_hd__nand3b_2 _20509_ (.A_N(_17246_),
    .B(_17331_),
    .C(_17332_),
    .Y(_17333_));
 sky130_fd_sc_hd__buf_1 _20510_ (.A(instr_andi),
    .X(_17334_));
 sky130_fd_sc_hd__buf_1 _20511_ (.A(_17334_),
    .X(_17335_));
 sky130_fd_sc_hd__o21ai_2 _20512_ (.A1(_17315_),
    .A2(_17328_),
    .B1(_17335_),
    .Y(_17336_));
 sky130_fd_sc_hd__a21oi_2 _20513_ (.A1(_17333_),
    .A2(_17336_),
    .B1(_17319_),
    .Y(_04008_));
 sky130_fd_sc_hd__buf_1 _20514_ (.A(_17255_),
    .X(_17337_));
 sky130_fd_sc_hd__nand3b_2 _20515_ (.A_N(_17263_),
    .B(_17332_),
    .C(_17337_),
    .Y(_17338_));
 sky130_fd_sc_hd__buf_1 _20516_ (.A(instr_ori),
    .X(_17339_));
 sky130_fd_sc_hd__buf_1 _20517_ (.A(_17339_),
    .X(_17340_));
 sky130_fd_sc_hd__buf_1 _20518_ (.A(_17258_),
    .X(_17341_));
 sky130_fd_sc_hd__buf_1 _20519_ (.A(_17341_),
    .X(_17342_));
 sky130_fd_sc_hd__a2bb2oi_2 _20520_ (.A1_N(_17273_),
    .A2_N(_17338_),
    .B1(_17340_),
    .B2(_17342_),
    .Y(_17343_));
 sky130_fd_sc_hd__nor2_2 _20521_ (.A(_17050_),
    .B(_17343_),
    .Y(_04007_));
 sky130_fd_sc_hd__buf_1 _20522_ (.A(_17332_),
    .X(_17344_));
 sky130_fd_sc_hd__buf_1 _20523_ (.A(_17330_),
    .X(_17345_));
 sky130_fd_sc_hd__nand3_2 _20524_ (.A(_17299_),
    .B(_17344_),
    .C(_17345_),
    .Y(_17346_));
 sky130_fd_sc_hd__buf_1 _20525_ (.A(instr_xori),
    .X(_17347_));
 sky130_fd_sc_hd__o21ai_2 _20526_ (.A1(_17315_),
    .A2(_17328_),
    .B1(_17347_),
    .Y(_17348_));
 sky130_fd_sc_hd__a21oi_2 _20527_ (.A1(_17346_),
    .A2(_17348_),
    .B1(_17319_),
    .Y(_04006_));
 sky130_fd_sc_hd__nand3_2 _20528_ (.A(_17307_),
    .B(_17344_),
    .C(_17345_),
    .Y(_17349_));
 sky130_fd_sc_hd__buf_1 _20529_ (.A(_17293_),
    .X(_17350_));
 sky130_fd_sc_hd__o21ai_2 _20530_ (.A1(_17350_),
    .A2(_17328_),
    .B1(instr_sltiu),
    .Y(_17351_));
 sky130_fd_sc_hd__buf_1 _20531_ (.A(_17318_),
    .X(_17352_));
 sky130_fd_sc_hd__a21oi_2 _20532_ (.A1(_17349_),
    .A2(_17351_),
    .B1(_17352_),
    .Y(_04005_));
 sky130_fd_sc_hd__nand3_2 _20533_ (.A(_17310_),
    .B(_17344_),
    .C(_17291_),
    .Y(_17353_));
 sky130_fd_sc_hd__buf_1 _20534_ (.A(_17301_),
    .X(_17354_));
 sky130_fd_sc_hd__o21ai_2 _20535_ (.A1(_17350_),
    .A2(_17354_),
    .B1(instr_slti),
    .Y(_17355_));
 sky130_fd_sc_hd__a21oi_2 _20536_ (.A1(_17353_),
    .A2(_17355_),
    .B1(_17352_),
    .Y(_04004_));
 sky130_fd_sc_hd__o21a_2 _20537_ (.A1(_17320_),
    .A2(_17267_),
    .B1(instr_addi),
    .X(_17356_));
 sky130_fd_sc_hd__buf_1 _20538_ (.A(_17322_),
    .X(_17357_));
 sky130_fd_sc_hd__nor2_2 _20539_ (.A(_17338_),
    .B(_17357_),
    .Y(_17358_));
 sky130_fd_sc_hd__o21a_2 _20540_ (.A1(_17356_),
    .A2(_17358_),
    .B1(_17326_),
    .X(_04003_));
 sky130_fd_sc_hd__nand3b_2 _20541_ (.A_N(_17246_),
    .B(_17331_),
    .C(_17226_),
    .Y(_17359_));
 sky130_fd_sc_hd__o21ai_2 _20542_ (.A1(_17350_),
    .A2(_17354_),
    .B1(instr_bgeu),
    .Y(_17360_));
 sky130_fd_sc_hd__a21oi_2 _20543_ (.A1(_17359_),
    .A2(_17360_),
    .B1(_17352_),
    .Y(_04002_));
 sky130_fd_sc_hd__buf_1 _20544_ (.A(_17284_),
    .X(_17361_));
 sky130_fd_sc_hd__nand3b_2 _20545_ (.A_N(_17264_),
    .B(_16980_),
    .C(_17361_),
    .Y(_17362_));
 sky130_fd_sc_hd__a2bb2oi_2 _20546_ (.A1_N(_17273_),
    .A2_N(_17362_),
    .B1(instr_bltu),
    .B2(_17342_),
    .Y(_17363_));
 sky130_fd_sc_hd__nor2_2 _20547_ (.A(_17050_),
    .B(_17363_),
    .Y(_04001_));
 sky130_fd_sc_hd__a2bb2oi_2 _20548_ (.A1_N(_17280_),
    .A2_N(_17362_),
    .B1(instr_bge),
    .B2(_17342_),
    .Y(_17364_));
 sky130_fd_sc_hd__nor2_2 _20549_ (.A(_17050_),
    .B(_17364_),
    .Y(_04000_));
 sky130_fd_sc_hd__nand3_2 _20550_ (.A(_17299_),
    .B(_17226_),
    .C(_17291_),
    .Y(_17365_));
 sky130_fd_sc_hd__o21ai_2 _20551_ (.A1(_17350_),
    .A2(_17354_),
    .B1(instr_blt),
    .Y(_17366_));
 sky130_fd_sc_hd__a21oi_2 _20552_ (.A1(_17365_),
    .A2(_17366_),
    .B1(_17352_),
    .Y(_03999_));
 sky130_fd_sc_hd__buf_1 _20553_ (.A(_17313_),
    .X(_17367_));
 sky130_fd_sc_hd__nand3_2 _20554_ (.A(_17367_),
    .B(_17226_),
    .C(_17291_),
    .Y(_17368_));
 sky130_fd_sc_hd__o21ai_2 _20555_ (.A1(_17320_),
    .A2(_17354_),
    .B1(instr_bne),
    .Y(_17369_));
 sky130_fd_sc_hd__buf_1 _20556_ (.A(_17318_),
    .X(_17370_));
 sky130_fd_sc_hd__a21oi_2 _20557_ (.A1(_17368_),
    .A2(_17369_),
    .B1(_17370_),
    .Y(_03998_));
 sky130_fd_sc_hd__o21a_2 _20558_ (.A1(_17320_),
    .A2(_17267_),
    .B1(instr_beq),
    .X(_17371_));
 sky130_fd_sc_hd__nor2_2 _20559_ (.A(_17362_),
    .B(_17357_),
    .Y(_17372_));
 sky130_fd_sc_hd__o21a_2 _20560_ (.A1(_17371_),
    .A2(_17372_),
    .B1(_17326_),
    .X(_03997_));
 sky130_vsdinv _20561_ (.A(\pcpi_timeout_counter[3] ),
    .Y(_17373_));
 sky130_fd_sc_hd__nor3_2 _20562_ (.A(\pcpi_timeout_counter[2] ),
    .B(\pcpi_timeout_counter[1] ),
    .C(\pcpi_timeout_counter[0] ),
    .Y(_17374_));
 sky130_fd_sc_hd__o21ai_2 _20563_ (.A1(_17373_),
    .A2(_17374_),
    .B1(_16945_),
    .Y(_03996_));
 sky130_fd_sc_hd__nor2_2 _20564_ (.A(\pcpi_timeout_counter[1] ),
    .B(\pcpi_timeout_counter[0] ),
    .Y(_17375_));
 sky130_fd_sc_hd__nand3b_2 _20565_ (.A_N(\pcpi_timeout_counter[2] ),
    .B(_17375_),
    .C(\pcpi_timeout_counter[3] ),
    .Y(_17376_));
 sky130_fd_sc_hd__buf_1 _20566_ (.A(\pcpi_timeout_counter[0] ),
    .X(_17377_));
 sky130_fd_sc_hd__o21ai_2 _20567_ (.A1(\pcpi_timeout_counter[1] ),
    .A2(_17377_),
    .B1(\pcpi_timeout_counter[2] ),
    .Y(_17378_));
 sky130_fd_sc_hd__nand3_2 _20568_ (.A(_17376_),
    .B(_16945_),
    .C(_17378_),
    .Y(_03995_));
 sky130_vsdinv _20569_ (.A(pcpi_valid),
    .Y(_17379_));
 sky130_fd_sc_hd__o21a_2 _20570_ (.A1(\pcpi_timeout_counter[3] ),
    .A2(\pcpi_timeout_counter[2] ),
    .B1(_17375_),
    .X(_17380_));
 sky130_fd_sc_hd__a2111o_2 _20571_ (.A1(\pcpi_timeout_counter[1] ),
    .A2(_17377_),
    .B1(_17109_),
    .C1(_17379_),
    .D1(_17380_),
    .X(_03994_));
 sky130_fd_sc_hd__a21o_2 _20572_ (.A1(_17374_),
    .A2(_17373_),
    .B1(_17377_),
    .X(_17381_));
 sky130_fd_sc_hd__nand3_2 _20573_ (.A(_17374_),
    .B(_17373_),
    .C(_17377_),
    .Y(_17382_));
 sky130_fd_sc_hd__nand3_2 _20574_ (.A(_17381_),
    .B(_16945_),
    .C(_17382_),
    .Y(_03993_));
 sky130_fd_sc_hd__and2b_2 _20575_ (.A_N(_17217_),
    .B(_16854_),
    .X(_17383_));
 sky130_fd_sc_hd__buf_1 _20576_ (.A(_16822_),
    .X(_17384_));
 sky130_fd_sc_hd__nand3_2 _20577_ (.A(_17383_),
    .B(_16985_),
    .C(_17384_),
    .Y(_17385_));
 sky130_fd_sc_hd__buf_1 _20578_ (.A(_16803_),
    .X(_17386_));
 sky130_fd_sc_hd__o21a_2 _20579_ (.A1(_16809_),
    .A2(_17386_),
    .B1(_16805_),
    .X(_17387_));
 sky130_fd_sc_hd__buf_1 _20580_ (.A(_17387_),
    .X(_00296_));
 sky130_fd_sc_hd__o32ai_2 _20581_ (.A1(_17076_),
    .A2(_17385_),
    .A3(_00296_),
    .B1(_00291_),
    .B2(_17056_),
    .Y(_03992_));
 sky130_fd_sc_hd__buf_1 _20582_ (.A(_16811_),
    .X(_17388_));
 sky130_fd_sc_hd__buf_1 _20583_ (.A(_16821_),
    .X(_17389_));
 sky130_fd_sc_hd__buf_1 _20584_ (.A(_17389_),
    .X(_17390_));
 sky130_fd_sc_hd__nand3b_2 _20585_ (.A_N(_17388_),
    .B(_17120_),
    .C(_17390_),
    .Y(_17391_));
 sky130_fd_sc_hd__o2bb2ai_2 _20586_ (.A1_N(_17388_),
    .A2_N(_17069_),
    .B1(_17391_),
    .B2(_00296_),
    .Y(_03991_));
 sky130_fd_sc_hd__buf_1 _20587_ (.A(_17044_),
    .X(_17392_));
 sky130_fd_sc_hd__buf_1 _20588_ (.A(_17026_),
    .X(_17393_));
 sky130_fd_sc_hd__buf_1 _20589_ (.A(_17393_),
    .X(_17394_));
 sky130_fd_sc_hd__or2_2 _20590_ (.A(\reg_next_pc[31] ),
    .B(_17394_),
    .X(_17395_));
 sky130_fd_sc_hd__o211a_2 _20591_ (.A1(_02530_),
    .A2(_17392_),
    .B1(_17227_),
    .C1(_17395_),
    .X(_03990_));
 sky130_fd_sc_hd__buf_1 _20592_ (.A(_17394_),
    .X(_17396_));
 sky130_fd_sc_hd__buf_1 _20593_ (.A(_17039_),
    .X(_17397_));
 sky130_fd_sc_hd__or2b_2 _20594_ (.A(_02529_),
    .B_N(_17397_),
    .X(_17398_));
 sky130_fd_sc_hd__o211a_2 _20595_ (.A1(_17396_),
    .A2(\reg_next_pc[30] ),
    .B1(_17227_),
    .C1(_17398_),
    .X(_03989_));
 sky130_fd_sc_hd__buf_1 _20596_ (.A(_17026_),
    .X(_17399_));
 sky130_fd_sc_hd__buf_1 _20597_ (.A(_17399_),
    .X(_17400_));
 sky130_fd_sc_hd__buf_1 _20598_ (.A(_17400_),
    .X(_17401_));
 sky130_fd_sc_hd__or2b_2 _20599_ (.A(_02527_),
    .B_N(_17397_),
    .X(_17402_));
 sky130_fd_sc_hd__o211a_2 _20600_ (.A1(_17401_),
    .A2(\reg_next_pc[29] ),
    .B1(_17227_),
    .C1(_17402_),
    .X(_03988_));
 sky130_fd_sc_hd__buf_1 _20601_ (.A(_17043_),
    .X(_17403_));
 sky130_fd_sc_hd__buf_1 _20602_ (.A(_17403_),
    .X(_00322_));
 sky130_fd_sc_hd__buf_1 _20603_ (.A(_16818_),
    .X(_17404_));
 sky130_fd_sc_hd__buf_1 _20604_ (.A(_17026_),
    .X(_17405_));
 sky130_fd_sc_hd__buf_1 _20605_ (.A(_17405_),
    .X(_17406_));
 sky130_fd_sc_hd__or2_2 _20606_ (.A(_17406_),
    .B(\reg_next_pc[28] ),
    .X(_17407_));
 sky130_fd_sc_hd__o211a_2 _20607_ (.A1(_00322_),
    .A2(_02526_),
    .B1(_17404_),
    .C1(_17407_),
    .X(_03987_));
 sky130_fd_sc_hd__or2b_2 _20608_ (.A(_02525_),
    .B_N(_17397_),
    .X(_17408_));
 sky130_fd_sc_hd__o211a_2 _20609_ (.A1(_17401_),
    .A2(\reg_next_pc[27] ),
    .B1(_17404_),
    .C1(_17408_),
    .X(_03986_));
 sky130_fd_sc_hd__buf_1 _20610_ (.A(_17403_),
    .X(_17409_));
 sky130_fd_sc_hd__or2_2 _20611_ (.A(_17406_),
    .B(\reg_next_pc[26] ),
    .X(_17410_));
 sky130_fd_sc_hd__o211a_2 _20612_ (.A1(_17409_),
    .A2(_02524_),
    .B1(_17404_),
    .C1(_17410_),
    .X(_03985_));
 sky130_fd_sc_hd__or2b_2 _20613_ (.A(_02523_),
    .B_N(_17397_),
    .X(_17411_));
 sky130_fd_sc_hd__o211a_2 _20614_ (.A1(_17401_),
    .A2(\reg_next_pc[25] ),
    .B1(_17404_),
    .C1(_17411_),
    .X(_03984_));
 sky130_fd_sc_hd__buf_1 _20615_ (.A(_16818_),
    .X(_17412_));
 sky130_fd_sc_hd__or2_2 _20616_ (.A(_17406_),
    .B(\reg_next_pc[24] ),
    .X(_17413_));
 sky130_fd_sc_hd__o211a_2 _20617_ (.A1(_17409_),
    .A2(_02522_),
    .B1(_17412_),
    .C1(_17413_),
    .X(_03983_));
 sky130_fd_sc_hd__buf_1 _20618_ (.A(_17027_),
    .X(_17414_));
 sky130_fd_sc_hd__buf_1 _20619_ (.A(_17414_),
    .X(_17415_));
 sky130_fd_sc_hd__or2b_2 _20620_ (.A(_02521_),
    .B_N(_17415_),
    .X(_17416_));
 sky130_fd_sc_hd__o211a_2 _20621_ (.A1(_17401_),
    .A2(\reg_next_pc[23] ),
    .B1(_17412_),
    .C1(_17416_),
    .X(_03982_));
 sky130_fd_sc_hd__buf_1 _20622_ (.A(_17400_),
    .X(_17417_));
 sky130_fd_sc_hd__or2b_2 _20623_ (.A(_02520_),
    .B_N(_17415_),
    .X(_17418_));
 sky130_fd_sc_hd__o211a_2 _20624_ (.A1(_17417_),
    .A2(\reg_next_pc[22] ),
    .B1(_17412_),
    .C1(_17418_),
    .X(_03981_));
 sky130_fd_sc_hd__or2_2 _20625_ (.A(_17406_),
    .B(\reg_next_pc[21] ),
    .X(_17419_));
 sky130_fd_sc_hd__o211a_2 _20626_ (.A1(_17409_),
    .A2(_02519_),
    .B1(_17412_),
    .C1(_17419_),
    .X(_03980_));
 sky130_fd_sc_hd__buf_1 _20627_ (.A(_16817_),
    .X(_17420_));
 sky130_fd_sc_hd__buf_1 _20628_ (.A(_17420_),
    .X(_17421_));
 sky130_fd_sc_hd__buf_1 _20629_ (.A(_17399_),
    .X(_17422_));
 sky130_fd_sc_hd__or2_2 _20630_ (.A(_17422_),
    .B(\reg_next_pc[20] ),
    .X(_17423_));
 sky130_fd_sc_hd__o211a_2 _20631_ (.A1(_17409_),
    .A2(_02518_),
    .B1(_17421_),
    .C1(_17423_),
    .X(_03979_));
 sky130_fd_sc_hd__buf_1 _20632_ (.A(_17043_),
    .X(_17424_));
 sky130_fd_sc_hd__buf_1 _20633_ (.A(_17424_),
    .X(_17425_));
 sky130_fd_sc_hd__or2_2 _20634_ (.A(_17422_),
    .B(\reg_next_pc[19] ),
    .X(_17426_));
 sky130_fd_sc_hd__o211a_2 _20635_ (.A1(_17425_),
    .A2(_02516_),
    .B1(_17421_),
    .C1(_17426_),
    .X(_03978_));
 sky130_fd_sc_hd__or2b_2 _20636_ (.A(_02515_),
    .B_N(_17415_),
    .X(_17427_));
 sky130_fd_sc_hd__o211a_2 _20637_ (.A1(_17417_),
    .A2(\reg_next_pc[18] ),
    .B1(_17421_),
    .C1(_17427_),
    .X(_03977_));
 sky130_fd_sc_hd__or2_2 _20638_ (.A(_17422_),
    .B(\reg_next_pc[17] ),
    .X(_17428_));
 sky130_fd_sc_hd__o211a_2 _20639_ (.A1(_17425_),
    .A2(_02514_),
    .B1(_17421_),
    .C1(_17428_),
    .X(_03976_));
 sky130_fd_sc_hd__buf_1 _20640_ (.A(_17420_),
    .X(_17429_));
 sky130_fd_sc_hd__or2b_2 _20641_ (.A(_02513_),
    .B_N(_17415_),
    .X(_17430_));
 sky130_fd_sc_hd__o211a_2 _20642_ (.A1(_17417_),
    .A2(\reg_next_pc[16] ),
    .B1(_17429_),
    .C1(_17430_),
    .X(_03975_));
 sky130_fd_sc_hd__or2_2 _20643_ (.A(_17422_),
    .B(\reg_next_pc[15] ),
    .X(_17431_));
 sky130_fd_sc_hd__o211a_2 _20644_ (.A1(_17425_),
    .A2(_02512_),
    .B1(_17429_),
    .C1(_17431_),
    .X(_03974_));
 sky130_fd_sc_hd__buf_1 _20645_ (.A(_17399_),
    .X(_17432_));
 sky130_fd_sc_hd__or2_2 _20646_ (.A(_17432_),
    .B(\reg_next_pc[14] ),
    .X(_17433_));
 sky130_fd_sc_hd__o211a_2 _20647_ (.A1(_17425_),
    .A2(_02511_),
    .B1(_17429_),
    .C1(_17433_),
    .X(_03973_));
 sky130_fd_sc_hd__buf_1 _20648_ (.A(_17424_),
    .X(_17434_));
 sky130_fd_sc_hd__or2_2 _20649_ (.A(_17432_),
    .B(\reg_next_pc[13] ),
    .X(_17435_));
 sky130_fd_sc_hd__o211a_2 _20650_ (.A1(_17434_),
    .A2(_02510_),
    .B1(_17429_),
    .C1(_17435_),
    .X(_03972_));
 sky130_fd_sc_hd__buf_1 _20651_ (.A(_17420_),
    .X(_17436_));
 sky130_fd_sc_hd__buf_1 _20652_ (.A(_17414_),
    .X(_17437_));
 sky130_fd_sc_hd__or2b_2 _20653_ (.A(_02509_),
    .B_N(_17437_),
    .X(_17438_));
 sky130_fd_sc_hd__o211a_2 _20654_ (.A1(_17417_),
    .A2(\reg_next_pc[12] ),
    .B1(_17436_),
    .C1(_17438_),
    .X(_03971_));
 sky130_fd_sc_hd__buf_1 _20655_ (.A(_17400_),
    .X(_17439_));
 sky130_fd_sc_hd__or2b_2 _20656_ (.A(_02508_),
    .B_N(_17437_),
    .X(_17440_));
 sky130_fd_sc_hd__o211a_2 _20657_ (.A1(_17439_),
    .A2(\reg_next_pc[11] ),
    .B1(_17436_),
    .C1(_17440_),
    .X(_03970_));
 sky130_fd_sc_hd__or2b_2 _20658_ (.A(_02507_),
    .B_N(_17437_),
    .X(_17441_));
 sky130_fd_sc_hd__o211a_2 _20659_ (.A1(_17439_),
    .A2(\reg_next_pc[10] ),
    .B1(_17436_),
    .C1(_17441_),
    .X(_03969_));
 sky130_fd_sc_hd__or2b_2 _20660_ (.A(_02537_),
    .B_N(_17437_),
    .X(_17442_));
 sky130_fd_sc_hd__o211a_2 _20661_ (.A1(_17439_),
    .A2(\reg_next_pc[9] ),
    .B1(_17436_),
    .C1(_17442_),
    .X(_03968_));
 sky130_fd_sc_hd__buf_1 _20662_ (.A(_17420_),
    .X(_17443_));
 sky130_fd_sc_hd__buf_1 _20663_ (.A(_17414_),
    .X(_17444_));
 sky130_fd_sc_hd__or2b_2 _20664_ (.A(_02536_),
    .B_N(_17444_),
    .X(_17445_));
 sky130_fd_sc_hd__o211a_2 _20665_ (.A1(_17439_),
    .A2(\reg_next_pc[8] ),
    .B1(_17443_),
    .C1(_17445_),
    .X(_03967_));
 sky130_fd_sc_hd__buf_1 _20666_ (.A(_17393_),
    .X(_17446_));
 sky130_fd_sc_hd__buf_1 _20667_ (.A(_17446_),
    .X(_17447_));
 sky130_fd_sc_hd__or2b_2 _20668_ (.A(_02535_),
    .B_N(_17444_),
    .X(_17448_));
 sky130_fd_sc_hd__o211a_2 _20669_ (.A1(_17447_),
    .A2(\reg_next_pc[7] ),
    .B1(_17443_),
    .C1(_17448_),
    .X(_03966_));
 sky130_fd_sc_hd__or2b_2 _20670_ (.A(_02534_),
    .B_N(_17444_),
    .X(_17449_));
 sky130_fd_sc_hd__o211a_2 _20671_ (.A1(_17447_),
    .A2(\reg_next_pc[6] ),
    .B1(_17443_),
    .C1(_17449_),
    .X(_03965_));
 sky130_fd_sc_hd__or2_2 _20672_ (.A(_17432_),
    .B(\reg_next_pc[5] ),
    .X(_17450_));
 sky130_fd_sc_hd__o211a_2 _20673_ (.A1(_17434_),
    .A2(_02533_),
    .B1(_17443_),
    .C1(_17450_),
    .X(_03964_));
 sky130_fd_sc_hd__buf_1 _20674_ (.A(_16816_),
    .X(_17451_));
 sky130_fd_sc_hd__buf_1 _20675_ (.A(_17451_),
    .X(_17452_));
 sky130_fd_sc_hd__buf_1 _20676_ (.A(_17452_),
    .X(_17453_));
 sky130_fd_sc_hd__or2b_2 _20677_ (.A(_02532_),
    .B_N(_17444_),
    .X(_17454_));
 sky130_fd_sc_hd__o211a_2 _20678_ (.A1(_17447_),
    .A2(\reg_next_pc[4] ),
    .B1(_17453_),
    .C1(_17454_),
    .X(_03963_));
 sky130_fd_sc_hd__buf_1 _20679_ (.A(_17414_),
    .X(_17455_));
 sky130_fd_sc_hd__or2b_2 _20680_ (.A(_02531_),
    .B_N(_17455_),
    .X(_17456_));
 sky130_fd_sc_hd__o211a_2 _20681_ (.A1(_17447_),
    .A2(\reg_next_pc[3] ),
    .B1(_17453_),
    .C1(_17456_),
    .X(_03962_));
 sky130_fd_sc_hd__buf_1 _20682_ (.A(_17446_),
    .X(_17457_));
 sky130_fd_sc_hd__or2b_2 _20683_ (.A(_02528_),
    .B_N(_17455_),
    .X(_17458_));
 sky130_fd_sc_hd__o211a_2 _20684_ (.A1(_17457_),
    .A2(\reg_next_pc[2] ),
    .B1(_17453_),
    .C1(_17458_),
    .X(_03961_));
 sky130_fd_sc_hd__or2b_2 _20685_ (.A(_02517_),
    .B_N(_17455_),
    .X(_17459_));
 sky130_fd_sc_hd__o211a_2 _20686_ (.A1(_17457_),
    .A2(\reg_next_pc[1] ),
    .B1(_17453_),
    .C1(_17459_),
    .X(_03960_));
 sky130_vsdinv _20687_ (.A(_02581_),
    .Y(_17460_));
 sky130_fd_sc_hd__buf_1 _20688_ (.A(_17039_),
    .X(_17461_));
 sky130_fd_sc_hd__nor2_2 _20689_ (.A(_17461_),
    .B(\reg_pc[31] ),
    .Y(_17462_));
 sky130_fd_sc_hd__a211oi_2 _20690_ (.A1(_17460_),
    .A2(_17396_),
    .B1(_16934_),
    .C1(_17462_),
    .Y(_03959_));
 sky130_fd_sc_hd__buf_1 _20691_ (.A(_02580_),
    .X(_17463_));
 sky130_vsdinv _20692_ (.A(_17463_),
    .Y(_17464_));
 sky130_fd_sc_hd__buf_1 _20693_ (.A(\reg_pc[30] ),
    .X(_17465_));
 sky130_fd_sc_hd__nor2_2 _20694_ (.A(_17461_),
    .B(_17465_),
    .Y(_17466_));
 sky130_fd_sc_hd__a211oi_2 _20695_ (.A1(_17464_),
    .A2(_17396_),
    .B1(_16934_),
    .C1(_17466_),
    .Y(_03958_));
 sky130_fd_sc_hd__buf_1 _20696_ (.A(\reg_pc[29] ),
    .X(_17467_));
 sky130_fd_sc_hd__buf_1 _20697_ (.A(_17452_),
    .X(_17468_));
 sky130_fd_sc_hd__buf_1 _20698_ (.A(_02579_),
    .X(_17469_));
 sky130_fd_sc_hd__or2b_2 _20699_ (.A(_17469_),
    .B_N(_17455_),
    .X(_17470_));
 sky130_fd_sc_hd__o211a_2 _20700_ (.A1(_17457_),
    .A2(_17467_),
    .B1(_17468_),
    .C1(_17470_),
    .X(_03957_));
 sky130_fd_sc_hd__buf_1 _20701_ (.A(\reg_pc[28] ),
    .X(_17471_));
 sky130_fd_sc_hd__buf_1 _20702_ (.A(_02578_),
    .X(_17472_));
 sky130_fd_sc_hd__buf_1 _20703_ (.A(_17405_),
    .X(_17473_));
 sky130_fd_sc_hd__or2b_2 _20704_ (.A(_17472_),
    .B_N(_17473_),
    .X(_17474_));
 sky130_fd_sc_hd__o211a_2 _20705_ (.A1(_17457_),
    .A2(_17471_),
    .B1(_17468_),
    .C1(_17474_),
    .X(_03956_));
 sky130_fd_sc_hd__buf_1 _20706_ (.A(_02577_),
    .X(_17475_));
 sky130_fd_sc_hd__buf_1 _20707_ (.A(\reg_pc[27] ),
    .X(_17476_));
 sky130_fd_sc_hd__or2_2 _20708_ (.A(_17432_),
    .B(_17476_),
    .X(_17477_));
 sky130_fd_sc_hd__o211a_2 _20709_ (.A1(_17434_),
    .A2(_17475_),
    .B1(_17468_),
    .C1(_17477_),
    .X(_03955_));
 sky130_fd_sc_hd__buf_1 _20710_ (.A(_02576_),
    .X(_17478_));
 sky130_fd_sc_hd__buf_1 _20711_ (.A(_17399_),
    .X(_17479_));
 sky130_fd_sc_hd__buf_1 _20712_ (.A(\reg_pc[26] ),
    .X(_17480_));
 sky130_fd_sc_hd__or2_2 _20713_ (.A(_17479_),
    .B(_17480_),
    .X(_17481_));
 sky130_fd_sc_hd__o211a_2 _20714_ (.A1(_17434_),
    .A2(_17478_),
    .B1(_17468_),
    .C1(_17481_),
    .X(_03954_));
 sky130_fd_sc_hd__buf_1 _20715_ (.A(_17446_),
    .X(_17482_));
 sky130_fd_sc_hd__buf_1 _20716_ (.A(\reg_pc[25] ),
    .X(_17483_));
 sky130_fd_sc_hd__buf_1 _20717_ (.A(_17483_),
    .X(_17484_));
 sky130_fd_sc_hd__buf_1 _20718_ (.A(_17452_),
    .X(_17485_));
 sky130_fd_sc_hd__buf_1 _20719_ (.A(_02575_),
    .X(_17486_));
 sky130_fd_sc_hd__buf_1 _20720_ (.A(_17486_),
    .X(_17487_));
 sky130_fd_sc_hd__or2b_2 _20721_ (.A(_17487_),
    .B_N(_17473_),
    .X(_17488_));
 sky130_fd_sc_hd__o211a_2 _20722_ (.A1(_17482_),
    .A2(_17484_),
    .B1(_17485_),
    .C1(_17488_),
    .X(_03953_));
 sky130_fd_sc_hd__buf_1 _20723_ (.A(\reg_pc[24] ),
    .X(_17489_));
 sky130_fd_sc_hd__buf_1 _20724_ (.A(_02574_),
    .X(_17490_));
 sky130_fd_sc_hd__or2b_2 _20725_ (.A(_17490_),
    .B_N(_17473_),
    .X(_17491_));
 sky130_fd_sc_hd__o211a_2 _20726_ (.A1(_17482_),
    .A2(_17489_),
    .B1(_17485_),
    .C1(_17491_),
    .X(_03952_));
 sky130_fd_sc_hd__buf_1 _20727_ (.A(\reg_pc[23] ),
    .X(_17492_));
 sky130_fd_sc_hd__buf_1 _20728_ (.A(_02573_),
    .X(_17493_));
 sky130_fd_sc_hd__buf_1 _20729_ (.A(_17493_),
    .X(_17494_));
 sky130_fd_sc_hd__or2b_2 _20730_ (.A(_17494_),
    .B_N(_17473_),
    .X(_17495_));
 sky130_fd_sc_hd__o211a_2 _20731_ (.A1(_17482_),
    .A2(_17492_),
    .B1(_17485_),
    .C1(_17495_),
    .X(_03951_));
 sky130_fd_sc_hd__buf_1 _20732_ (.A(_17424_),
    .X(_17496_));
 sky130_fd_sc_hd__buf_1 _20733_ (.A(_02572_),
    .X(_17497_));
 sky130_vsdinv _20734_ (.A(\reg_pc[22] ),
    .Y(_17498_));
 sky130_fd_sc_hd__nand2_2 _20735_ (.A(_17392_),
    .B(_17498_),
    .Y(_17499_));
 sky130_fd_sc_hd__o211a_2 _20736_ (.A1(_17496_),
    .A2(_17497_),
    .B1(_17485_),
    .C1(_17499_),
    .X(_03950_));
 sky130_fd_sc_hd__buf_1 _20737_ (.A(_02570_),
    .X(_17500_));
 sky130_fd_sc_hd__buf_1 _20738_ (.A(_17500_),
    .X(_17501_));
 sky130_fd_sc_hd__buf_1 _20739_ (.A(_17452_),
    .X(_17502_));
 sky130_fd_sc_hd__buf_1 _20740_ (.A(\reg_pc[21] ),
    .X(_17503_));
 sky130_fd_sc_hd__or2_2 _20741_ (.A(_17479_),
    .B(_17503_),
    .X(_17504_));
 sky130_fd_sc_hd__o211a_2 _20742_ (.A1(_17496_),
    .A2(_17501_),
    .B1(_17502_),
    .C1(_17504_),
    .X(_03949_));
 sky130_fd_sc_hd__buf_1 _20743_ (.A(_02569_),
    .X(_17505_));
 sky130_fd_sc_hd__buf_1 _20744_ (.A(_17505_),
    .X(_17506_));
 sky130_vsdinv _20745_ (.A(\reg_pc[20] ),
    .Y(_17507_));
 sky130_fd_sc_hd__nand2_2 _20746_ (.A(_17392_),
    .B(_17507_),
    .Y(_17508_));
 sky130_fd_sc_hd__o211a_2 _20747_ (.A1(_17496_),
    .A2(_17506_),
    .B1(_17502_),
    .C1(_17508_),
    .X(_03948_));
 sky130_fd_sc_hd__buf_1 _20748_ (.A(\reg_pc[19] ),
    .X(_17509_));
 sky130_fd_sc_hd__buf_1 _20749_ (.A(_17509_),
    .X(_17510_));
 sky130_fd_sc_hd__buf_1 _20750_ (.A(_02568_),
    .X(_17511_));
 sky130_fd_sc_hd__buf_1 _20751_ (.A(_17405_),
    .X(_17512_));
 sky130_fd_sc_hd__or2b_2 _20752_ (.A(_17511_),
    .B_N(_17512_),
    .X(_17513_));
 sky130_fd_sc_hd__o211a_2 _20753_ (.A1(_17482_),
    .A2(_17510_),
    .B1(_17502_),
    .C1(_17513_),
    .X(_03947_));
 sky130_fd_sc_hd__buf_1 _20754_ (.A(_17446_),
    .X(_17514_));
 sky130_fd_sc_hd__buf_1 _20755_ (.A(\reg_pc[18] ),
    .X(_17515_));
 sky130_fd_sc_hd__buf_1 _20756_ (.A(_17515_),
    .X(_17516_));
 sky130_fd_sc_hd__buf_1 _20757_ (.A(_02567_),
    .X(_17517_));
 sky130_fd_sc_hd__buf_1 _20758_ (.A(_17517_),
    .X(_17518_));
 sky130_fd_sc_hd__or2b_2 _20759_ (.A(_17518_),
    .B_N(_17512_),
    .X(_17519_));
 sky130_fd_sc_hd__o211a_2 _20760_ (.A1(_17514_),
    .A2(_17516_),
    .B1(_17502_),
    .C1(_17519_),
    .X(_03946_));
 sky130_fd_sc_hd__buf_1 _20761_ (.A(_02566_),
    .X(_17520_));
 sky130_fd_sc_hd__buf_1 _20762_ (.A(_17451_),
    .X(_17521_));
 sky130_fd_sc_hd__buf_1 _20763_ (.A(_17521_),
    .X(_17522_));
 sky130_fd_sc_hd__buf_1 _20764_ (.A(\reg_pc[17] ),
    .X(_17523_));
 sky130_fd_sc_hd__buf_1 _20765_ (.A(_17523_),
    .X(_17524_));
 sky130_fd_sc_hd__or2_2 _20766_ (.A(_17479_),
    .B(_17524_),
    .X(_17525_));
 sky130_fd_sc_hd__o211a_2 _20767_ (.A1(_17496_),
    .A2(_17520_),
    .B1(_17522_),
    .C1(_17525_),
    .X(_03945_));
 sky130_fd_sc_hd__buf_1 _20768_ (.A(\reg_pc[16] ),
    .X(_17526_));
 sky130_fd_sc_hd__buf_1 _20769_ (.A(_02565_),
    .X(_17527_));
 sky130_fd_sc_hd__or2b_2 _20770_ (.A(_17527_),
    .B_N(_17512_),
    .X(_17528_));
 sky130_fd_sc_hd__o211a_2 _20771_ (.A1(_17514_),
    .A2(_17526_),
    .B1(_17522_),
    .C1(_17528_),
    .X(_03944_));
 sky130_fd_sc_hd__buf_1 _20772_ (.A(\reg_pc[15] ),
    .X(_17529_));
 sky130_fd_sc_hd__buf_1 _20773_ (.A(_17529_),
    .X(_17530_));
 sky130_fd_sc_hd__buf_1 _20774_ (.A(_02564_),
    .X(_17531_));
 sky130_fd_sc_hd__or2b_2 _20775_ (.A(_17531_),
    .B_N(_17512_),
    .X(_17532_));
 sky130_fd_sc_hd__o211a_2 _20776_ (.A1(_17514_),
    .A2(_17530_),
    .B1(_17522_),
    .C1(_17532_),
    .X(_03943_));
 sky130_fd_sc_hd__buf_1 _20777_ (.A(_17424_),
    .X(_17533_));
 sky130_fd_sc_hd__buf_1 _20778_ (.A(_02563_),
    .X(_17534_));
 sky130_fd_sc_hd__buf_1 _20779_ (.A(\reg_pc[14] ),
    .X(_17535_));
 sky130_fd_sc_hd__buf_1 _20780_ (.A(_17535_),
    .X(_17536_));
 sky130_fd_sc_hd__or2_2 _20781_ (.A(_17479_),
    .B(_17536_),
    .X(_17537_));
 sky130_fd_sc_hd__o211a_2 _20782_ (.A1(_17533_),
    .A2(_17534_),
    .B1(_17522_),
    .C1(_17537_),
    .X(_03942_));
 sky130_fd_sc_hd__buf_1 _20783_ (.A(\reg_pc[13] ),
    .X(_17538_));
 sky130_fd_sc_hd__buf_1 _20784_ (.A(_17538_),
    .X(_17539_));
 sky130_fd_sc_hd__buf_1 _20785_ (.A(_17521_),
    .X(_17540_));
 sky130_fd_sc_hd__buf_1 _20786_ (.A(_02562_),
    .X(_17541_));
 sky130_fd_sc_hd__buf_1 _20787_ (.A(_17405_),
    .X(_17542_));
 sky130_fd_sc_hd__or2b_2 _20788_ (.A(_17541_),
    .B_N(_17542_),
    .X(_17543_));
 sky130_fd_sc_hd__o211a_2 _20789_ (.A1(_17514_),
    .A2(_17539_),
    .B1(_17540_),
    .C1(_17543_),
    .X(_03941_));
 sky130_fd_sc_hd__buf_1 _20790_ (.A(_02561_),
    .X(_17544_));
 sky130_fd_sc_hd__buf_1 _20791_ (.A(\reg_pc[12] ),
    .X(_17545_));
 sky130_fd_sc_hd__inv_2 _20792_ (.A(_17545_),
    .Y(_17546_));
 sky130_fd_sc_hd__nand2_2 _20793_ (.A(_17045_),
    .B(_17546_),
    .Y(_17547_));
 sky130_fd_sc_hd__o211a_2 _20794_ (.A1(_17533_),
    .A2(_17544_),
    .B1(_17540_),
    .C1(_17547_),
    .X(_03940_));
 sky130_fd_sc_hd__buf_1 _20795_ (.A(_17394_),
    .X(_17548_));
 sky130_fd_sc_hd__buf_1 _20796_ (.A(\reg_pc[11] ),
    .X(_17549_));
 sky130_fd_sc_hd__buf_1 _20797_ (.A(_02589_),
    .X(_17550_));
 sky130_fd_sc_hd__or2b_2 _20798_ (.A(_17550_),
    .B_N(_17542_),
    .X(_17551_));
 sky130_fd_sc_hd__o211a_2 _20799_ (.A1(_17548_),
    .A2(_17549_),
    .B1(_17540_),
    .C1(_17551_),
    .X(_03939_));
 sky130_fd_sc_hd__buf_1 _20800_ (.A(\reg_pc[10] ),
    .X(_17552_));
 sky130_fd_sc_hd__buf_1 _20801_ (.A(_17552_),
    .X(_17553_));
 sky130_fd_sc_hd__buf_1 _20802_ (.A(_02588_),
    .X(_17554_));
 sky130_fd_sc_hd__buf_1 _20803_ (.A(_17554_),
    .X(_17555_));
 sky130_fd_sc_hd__or2b_2 _20804_ (.A(_17555_),
    .B_N(_17542_),
    .X(_17556_));
 sky130_fd_sc_hd__o211a_2 _20805_ (.A1(_17548_),
    .A2(_17553_),
    .B1(_17540_),
    .C1(_17556_),
    .X(_03938_));
 sky130_fd_sc_hd__buf_1 _20806_ (.A(\reg_pc[9] ),
    .X(_17557_));
 sky130_fd_sc_hd__buf_1 _20807_ (.A(_17557_),
    .X(_17558_));
 sky130_fd_sc_hd__buf_1 _20808_ (.A(_17521_),
    .X(_17559_));
 sky130_vsdinv _20809_ (.A(_02587_),
    .Y(_17560_));
 sky130_fd_sc_hd__buf_1 _20810_ (.A(_17039_),
    .X(_17561_));
 sky130_fd_sc_hd__nand2_2 _20811_ (.A(_17560_),
    .B(_17561_),
    .Y(_17562_));
 sky130_fd_sc_hd__o211a_2 _20812_ (.A1(_17548_),
    .A2(_17558_),
    .B1(_17559_),
    .C1(_17562_),
    .X(_03937_));
 sky130_fd_sc_hd__buf_1 _20813_ (.A(_02586_),
    .X(_17563_));
 sky130_fd_sc_hd__buf_1 _20814_ (.A(_17563_),
    .X(_17564_));
 sky130_fd_sc_hd__inv_2 _20815_ (.A(\reg_pc[8] ),
    .Y(_17565_));
 sky130_fd_sc_hd__nand2_2 _20816_ (.A(_17045_),
    .B(_17565_),
    .Y(_17566_));
 sky130_fd_sc_hd__o211a_2 _20817_ (.A1(_17533_),
    .A2(_17564_),
    .B1(_17559_),
    .C1(_17566_),
    .X(_03936_));
 sky130_fd_sc_hd__buf_1 _20818_ (.A(\reg_pc[7] ),
    .X(_17567_));
 sky130_vsdinv _20819_ (.A(_02585_),
    .Y(_17568_));
 sky130_fd_sc_hd__nand2_2 _20820_ (.A(_17568_),
    .B(_17561_),
    .Y(_17569_));
 sky130_fd_sc_hd__o211a_2 _20821_ (.A1(_17548_),
    .A2(_17567_),
    .B1(_17559_),
    .C1(_17569_),
    .X(_03935_));
 sky130_fd_sc_hd__buf_1 _20822_ (.A(_17394_),
    .X(_17570_));
 sky130_fd_sc_hd__buf_1 _20823_ (.A(\reg_pc[6] ),
    .X(_17571_));
 sky130_fd_sc_hd__buf_1 _20824_ (.A(_02584_),
    .X(_17572_));
 sky130_fd_sc_hd__or2b_2 _20825_ (.A(_17572_),
    .B_N(_17542_),
    .X(_17573_));
 sky130_fd_sc_hd__o211a_2 _20826_ (.A1(_17570_),
    .A2(_17571_),
    .B1(_17559_),
    .C1(_17573_),
    .X(_03934_));
 sky130_fd_sc_hd__buf_1 _20827_ (.A(\reg_pc[5] ),
    .X(_17574_));
 sky130_fd_sc_hd__buf_1 _20828_ (.A(_17574_),
    .X(_17575_));
 sky130_fd_sc_hd__buf_1 _20829_ (.A(_17521_),
    .X(_17576_));
 sky130_vsdinv _20830_ (.A(_02583_),
    .Y(_17577_));
 sky130_fd_sc_hd__nand2_2 _20831_ (.A(_17577_),
    .B(_17561_),
    .Y(_17578_));
 sky130_fd_sc_hd__o211a_2 _20832_ (.A1(_17570_),
    .A2(_17575_),
    .B1(_17576_),
    .C1(_17578_),
    .X(_03933_));
 sky130_fd_sc_hd__buf_1 _20833_ (.A(_01475_),
    .X(_17579_));
 sky130_fd_sc_hd__buf_1 _20834_ (.A(\reg_pc[4] ),
    .X(_17580_));
 sky130_fd_sc_hd__buf_1 _20835_ (.A(_17580_),
    .X(_17581_));
 sky130_fd_sc_hd__nor2_2 _20836_ (.A(_17461_),
    .B(_17581_),
    .Y(_17582_));
 sky130_fd_sc_hd__a211oi_2 _20837_ (.A1(_17396_),
    .A2(_17579_),
    .B1(_16934_),
    .C1(_17582_),
    .Y(_03932_));
 sky130_vsdinv _20838_ (.A(_01475_),
    .Y(_17583_));
 sky130_fd_sc_hd__buf_1 _20839_ (.A(_17583_),
    .X(_02582_));
 sky130_fd_sc_hd__buf_1 _20840_ (.A(\reg_pc[3] ),
    .X(_17584_));
 sky130_fd_sc_hd__buf_1 _20841_ (.A(_17584_),
    .X(_17585_));
 sky130_fd_sc_hd__buf_1 _20842_ (.A(_02571_),
    .X(_17586_));
 sky130_fd_sc_hd__buf_1 _20843_ (.A(_17586_),
    .X(_17587_));
 sky130_vsdinv _20844_ (.A(_17587_),
    .Y(_17588_));
 sky130_fd_sc_hd__nand2_2 _20845_ (.A(_17588_),
    .B(_17561_),
    .Y(_17589_));
 sky130_fd_sc_hd__o211a_2 _20846_ (.A1(_17570_),
    .A2(_17585_),
    .B1(_17576_),
    .C1(_17589_),
    .X(_03931_));
 sky130_fd_sc_hd__buf_1 _20847_ (.A(\reg_pc[2] ),
    .X(_17590_));
 sky130_fd_sc_hd__buf_1 _20848_ (.A(_17590_),
    .X(_17591_));
 sky130_fd_sc_hd__buf_1 _20849_ (.A(_02560_),
    .X(_17592_));
 sky130_fd_sc_hd__inv_2 _20850_ (.A(_17592_),
    .Y(_01561_));
 sky130_fd_sc_hd__nand2_2 _20851_ (.A(_01561_),
    .B(_17461_),
    .Y(_17593_));
 sky130_fd_sc_hd__o211a_2 _20852_ (.A1(_17570_),
    .A2(_17591_),
    .B1(_17576_),
    .C1(_17593_),
    .X(_03930_));
 sky130_fd_sc_hd__buf_1 _20853_ (.A(\reg_pc[1] ),
    .X(_17594_));
 sky130_fd_sc_hd__or2_2 _20854_ (.A(_17400_),
    .B(_17594_),
    .X(_17595_));
 sky130_fd_sc_hd__o211a_2 _20855_ (.A1(_17533_),
    .A2(_02590_),
    .B1(_17576_),
    .C1(_17595_),
    .X(_03929_));
 sky130_vsdinv _20856_ (.A(\count_instr[62] ),
    .Y(_17596_));
 sky130_vsdinv _20857_ (.A(\count_instr[59] ),
    .Y(_17597_));
 sky130_vsdinv _20858_ (.A(\count_instr[58] ),
    .Y(_17598_));
 sky130_vsdinv _20859_ (.A(\count_instr[53] ),
    .Y(_17599_));
 sky130_fd_sc_hd__nand2_2 _20860_ (.A(\count_instr[55] ),
    .B(\count_instr[54] ),
    .Y(_17600_));
 sky130_vsdinv _20861_ (.A(\count_instr[50] ),
    .Y(_17601_));
 sky130_vsdinv _20862_ (.A(\count_instr[49] ),
    .Y(_17602_));
 sky130_vsdinv _20863_ (.A(\count_instr[43] ),
    .Y(_17603_));
 sky130_vsdinv _20864_ (.A(\count_instr[42] ),
    .Y(_17604_));
 sky130_vsdinv _20865_ (.A(\count_instr[37] ),
    .Y(_17605_));
 sky130_fd_sc_hd__nand2_2 _20866_ (.A(\count_instr[39] ),
    .B(\count_instr[38] ),
    .Y(_17606_));
 sky130_vsdinv _20867_ (.A(\count_instr[34] ),
    .Y(_17607_));
 sky130_vsdinv _20868_ (.A(\count_instr[33] ),
    .Y(_17608_));
 sky130_vsdinv _20869_ (.A(\count_instr[24] ),
    .Y(_17609_));
 sky130_fd_sc_hd__nand2_2 _20870_ (.A(\count_instr[23] ),
    .B(\count_instr[22] ),
    .Y(_17610_));
 sky130_fd_sc_hd__nand3_2 _20871_ (.A(\count_instr[4] ),
    .B(\count_instr[3] ),
    .C(\count_instr[0] ),
    .Y(_17611_));
 sky130_fd_sc_hd__nand2_2 _20872_ (.A(\count_instr[6] ),
    .B(\count_instr[5] ),
    .Y(_17612_));
 sky130_fd_sc_hd__nand3b_2 _20873_ (.A_N(_17612_),
    .B(\count_instr[8] ),
    .C(\count_instr[7] ),
    .Y(_17613_));
 sky130_fd_sc_hd__and4_2 _20874_ (.A(\count_instr[12] ),
    .B(\count_instr[11] ),
    .C(\count_instr[10] ),
    .D(\count_instr[9] ),
    .X(_17614_));
 sky130_fd_sc_hd__nand3_2 _20875_ (.A(_17614_),
    .B(\count_instr[2] ),
    .C(\count_instr[1] ),
    .Y(_17615_));
 sky130_fd_sc_hd__nor3_2 _20876_ (.A(_17611_),
    .B(_17613_),
    .C(_17615_),
    .Y(_17616_));
 sky130_vsdinv _20877_ (.A(_17616_),
    .Y(_17617_));
 sky130_fd_sc_hd__nor2_2 _20878_ (.A(_17617_),
    .B(_16928_),
    .Y(_17618_));
 sky130_fd_sc_hd__and2_2 _20879_ (.A(\count_instr[15] ),
    .B(\count_instr[14] ),
    .X(_17619_));
 sky130_fd_sc_hd__and4_2 _20880_ (.A(_17618_),
    .B(\count_instr[16] ),
    .C(\count_instr[13] ),
    .D(_17619_),
    .X(_17620_));
 sky130_fd_sc_hd__and4_2 _20881_ (.A(_17620_),
    .B(\count_instr[19] ),
    .C(\count_instr[18] ),
    .D(\count_instr[17] ),
    .X(_17621_));
 sky130_fd_sc_hd__nand3_2 _20882_ (.A(_17621_),
    .B(\count_instr[21] ),
    .C(\count_instr[20] ),
    .Y(_17622_));
 sky130_fd_sc_hd__nor3_2 _20883_ (.A(_17609_),
    .B(_17610_),
    .C(_17622_),
    .Y(_17623_));
 sky130_fd_sc_hd__and4_2 _20884_ (.A(_17623_),
    .B(\count_instr[27] ),
    .C(\count_instr[26] ),
    .D(\count_instr[25] ),
    .X(_17624_));
 sky130_fd_sc_hd__and4_2 _20885_ (.A(\count_instr[31] ),
    .B(\count_instr[30] ),
    .C(\count_instr[29] ),
    .D(\count_instr[28] ),
    .X(_17625_));
 sky130_fd_sc_hd__nand3_2 _20886_ (.A(_17624_),
    .B(\count_instr[32] ),
    .C(_17625_),
    .Y(_17626_));
 sky130_fd_sc_hd__nor3_2 _20887_ (.A(_17607_),
    .B(_17608_),
    .C(_17626_),
    .Y(_17627_));
 sky130_fd_sc_hd__nand3_2 _20888_ (.A(_17627_),
    .B(\count_instr[36] ),
    .C(\count_instr[35] ),
    .Y(_17628_));
 sky130_fd_sc_hd__nor3_2 _20889_ (.A(_17605_),
    .B(_17606_),
    .C(_17628_),
    .Y(_17629_));
 sky130_fd_sc_hd__nand3_2 _20890_ (.A(_17629_),
    .B(\count_instr[41] ),
    .C(\count_instr[40] ),
    .Y(_17630_));
 sky130_fd_sc_hd__nor3_2 _20891_ (.A(_17603_),
    .B(_17604_),
    .C(_17630_),
    .Y(_17631_));
 sky130_fd_sc_hd__and4_2 _20892_ (.A(\count_instr[47] ),
    .B(\count_instr[46] ),
    .C(\count_instr[45] ),
    .D(\count_instr[44] ),
    .X(_17632_));
 sky130_fd_sc_hd__nand3_2 _20893_ (.A(_17631_),
    .B(\count_instr[48] ),
    .C(_17632_),
    .Y(_17633_));
 sky130_fd_sc_hd__nor3_2 _20894_ (.A(_17601_),
    .B(_17602_),
    .C(_17633_),
    .Y(_17634_));
 sky130_fd_sc_hd__nand3_2 _20895_ (.A(_17634_),
    .B(\count_instr[52] ),
    .C(\count_instr[51] ),
    .Y(_17635_));
 sky130_fd_sc_hd__nor3_2 _20896_ (.A(_17599_),
    .B(_17600_),
    .C(_17635_),
    .Y(_17636_));
 sky130_fd_sc_hd__nand3_2 _20897_ (.A(_17636_),
    .B(\count_instr[57] ),
    .C(\count_instr[56] ),
    .Y(_17637_));
 sky130_fd_sc_hd__nor3_2 _20898_ (.A(_17597_),
    .B(_17598_),
    .C(_17637_),
    .Y(_17638_));
 sky130_fd_sc_hd__nand3_2 _20899_ (.A(_17638_),
    .B(\count_instr[61] ),
    .C(\count_instr[60] ),
    .Y(_17639_));
 sky130_fd_sc_hd__nor3b_2 _20900_ (.A(_17596_),
    .B(_17639_),
    .C_N(\count_instr[63] ),
    .Y(_17640_));
 sky130_fd_sc_hd__nor2_2 _20901_ (.A(_17596_),
    .B(_17639_),
    .Y(_17641_));
 sky130_fd_sc_hd__o21bai_2 _20902_ (.A1(\count_instr[63] ),
    .A2(_17641_),
    .B1_N(_16933_),
    .Y(_17642_));
 sky130_fd_sc_hd__nor2_2 _20903_ (.A(_17640_),
    .B(_17642_),
    .Y(_03928_));
 sky130_fd_sc_hd__buf_1 _20904_ (.A(_17638_),
    .X(_17643_));
 sky130_fd_sc_hd__buf_1 _20905_ (.A(\count_instr[61] ),
    .X(_17644_));
 sky130_fd_sc_hd__a31oi_2 _20906_ (.A1(_17643_),
    .A2(_17644_),
    .A3(\count_instr[60] ),
    .B1(\count_instr[62] ),
    .Y(_17645_));
 sky130_fd_sc_hd__nor3_2 _20907_ (.A(_17370_),
    .B(_17645_),
    .C(_17641_),
    .Y(_03927_));
 sky130_fd_sc_hd__buf_1 _20908_ (.A(_17637_),
    .X(_17646_));
 sky130_fd_sc_hd__nor2_2 _20909_ (.A(_17598_),
    .B(_17646_),
    .Y(_17647_));
 sky130_fd_sc_hd__buf_1 _20910_ (.A(\count_instr[59] ),
    .X(_17648_));
 sky130_fd_sc_hd__and3_2 _20911_ (.A(_17647_),
    .B(\count_instr[60] ),
    .C(_17648_),
    .X(_17649_));
 sky130_fd_sc_hd__buf_1 _20912_ (.A(\count_instr[60] ),
    .X(_17650_));
 sky130_fd_sc_hd__buf_1 _20913_ (.A(_17148_),
    .X(_17651_));
 sky130_fd_sc_hd__a31oi_2 _20914_ (.A1(_17643_),
    .A2(_17644_),
    .A3(_17650_),
    .B1(_17651_),
    .Y(_17652_));
 sky130_fd_sc_hd__o21a_2 _20915_ (.A1(_17644_),
    .A2(_17649_),
    .B1(_17652_),
    .X(_03926_));
 sky130_fd_sc_hd__a31oi_2 _20916_ (.A1(_17647_),
    .A2(_17650_),
    .A3(_17648_),
    .B1(_17651_),
    .Y(_17653_));
 sky130_fd_sc_hd__o21a_2 _20917_ (.A1(_17650_),
    .A2(_17643_),
    .B1(_17653_),
    .X(_03925_));
 sky130_fd_sc_hd__buf_1 _20918_ (.A(_17318_),
    .X(_17654_));
 sky130_fd_sc_hd__buf_1 _20919_ (.A(_17636_),
    .X(_17655_));
 sky130_fd_sc_hd__a41oi_2 _20920_ (.A1(\count_instr[58] ),
    .A2(_17655_),
    .A3(\count_instr[57] ),
    .A4(\count_instr[56] ),
    .B1(_17648_),
    .Y(_17656_));
 sky130_fd_sc_hd__nor3_2 _20921_ (.A(_17654_),
    .B(_17656_),
    .C(_17643_),
    .Y(_03924_));
 sky130_fd_sc_hd__buf_1 _20922_ (.A(_16932_),
    .X(_17657_));
 sky130_fd_sc_hd__o21bai_2 _20923_ (.A1(_17598_),
    .A2(_17646_),
    .B1_N(_17657_),
    .Y(_17658_));
 sky130_fd_sc_hd__a21oi_2 _20924_ (.A1(_17598_),
    .A2(_17646_),
    .B1(_17658_),
    .Y(_03923_));
 sky130_fd_sc_hd__buf_1 _20925_ (.A(\count_instr[56] ),
    .X(_17659_));
 sky130_fd_sc_hd__a21oi_2 _20926_ (.A1(_17655_),
    .A2(_17659_),
    .B1(\count_instr[57] ),
    .Y(_17660_));
 sky130_vsdinv _20927_ (.A(_17646_),
    .Y(_17661_));
 sky130_fd_sc_hd__nor3_2 _20928_ (.A(_17654_),
    .B(_17660_),
    .C(_17661_),
    .Y(_03922_));
 sky130_fd_sc_hd__a21oi_2 _20929_ (.A1(_17655_),
    .A2(_17659_),
    .B1(_17197_),
    .Y(_17662_));
 sky130_fd_sc_hd__o21a_2 _20930_ (.A1(_17659_),
    .A2(_17655_),
    .B1(_17662_),
    .X(_03921_));
 sky130_fd_sc_hd__buf_1 _20931_ (.A(_17599_),
    .X(_17663_));
 sky130_fd_sc_hd__buf_1 _20932_ (.A(_17635_),
    .X(_17664_));
 sky130_fd_sc_hd__nor2_2 _20933_ (.A(_17663_),
    .B(_17664_),
    .Y(_17665_));
 sky130_fd_sc_hd__buf_1 _20934_ (.A(\count_instr[54] ),
    .X(_17666_));
 sky130_fd_sc_hd__and3_2 _20935_ (.A(_17665_),
    .B(\count_instr[55] ),
    .C(_17666_),
    .X(_17667_));
 sky130_fd_sc_hd__nor3b_2 _20936_ (.A(_17663_),
    .B(_17664_),
    .C_N(_17666_),
    .Y(_17668_));
 sky130_fd_sc_hd__o21bai_2 _20937_ (.A1(\count_instr[55] ),
    .A2(_17668_),
    .B1_N(_16933_),
    .Y(_17669_));
 sky130_fd_sc_hd__nor2_2 _20938_ (.A(_17667_),
    .B(_17669_),
    .Y(_03920_));
 sky130_fd_sc_hd__buf_1 _20939_ (.A(_17634_),
    .X(_17670_));
 sky130_fd_sc_hd__buf_1 _20940_ (.A(\count_instr[52] ),
    .X(_17671_));
 sky130_fd_sc_hd__a41oi_2 _20941_ (.A1(\count_instr[53] ),
    .A2(_17670_),
    .A3(_17671_),
    .A4(\count_instr[51] ),
    .B1(_17666_),
    .Y(_17672_));
 sky130_fd_sc_hd__nor3_2 _20942_ (.A(_17654_),
    .B(_17672_),
    .C(_17668_),
    .Y(_03919_));
 sky130_fd_sc_hd__o21bai_2 _20943_ (.A1(_17663_),
    .A2(_17664_),
    .B1_N(_17657_),
    .Y(_17673_));
 sky130_fd_sc_hd__a21oi_2 _20944_ (.A1(_17663_),
    .A2(_17664_),
    .B1(_17673_),
    .Y(_03918_));
 sky130_fd_sc_hd__nor2_2 _20945_ (.A(_17602_),
    .B(_17633_),
    .Y(_17674_));
 sky130_fd_sc_hd__buf_1 _20946_ (.A(\count_instr[50] ),
    .X(_17675_));
 sky130_fd_sc_hd__and3_2 _20947_ (.A(_17674_),
    .B(\count_instr[51] ),
    .C(_17675_),
    .X(_17676_));
 sky130_fd_sc_hd__buf_1 _20948_ (.A(\count_instr[51] ),
    .X(_17677_));
 sky130_fd_sc_hd__a31oi_2 _20949_ (.A1(_17670_),
    .A2(_17671_),
    .A3(_17677_),
    .B1(_17651_),
    .Y(_17678_));
 sky130_fd_sc_hd__o21a_2 _20950_ (.A1(_17671_),
    .A2(_17676_),
    .B1(_17678_),
    .X(_03917_));
 sky130_fd_sc_hd__a31oi_2 _20951_ (.A1(_17674_),
    .A2(_17677_),
    .A3(_17675_),
    .B1(_17651_),
    .Y(_17679_));
 sky130_fd_sc_hd__o21a_2 _20952_ (.A1(_17677_),
    .A2(_17670_),
    .B1(_17679_),
    .X(_03916_));
 sky130_fd_sc_hd__buf_1 _20953_ (.A(_17631_),
    .X(_17680_));
 sky130_fd_sc_hd__buf_1 _20954_ (.A(\count_instr[48] ),
    .X(_17681_));
 sky130_fd_sc_hd__a41oi_2 _20955_ (.A1(\count_instr[49] ),
    .A2(_17680_),
    .A3(_17681_),
    .A4(_17632_),
    .B1(_17675_),
    .Y(_17682_));
 sky130_fd_sc_hd__nor3_2 _20956_ (.A(_17654_),
    .B(_17682_),
    .C(_17670_),
    .Y(_03915_));
 sky130_fd_sc_hd__buf_1 _20957_ (.A(_16932_),
    .X(_17683_));
 sky130_fd_sc_hd__o21bai_2 _20958_ (.A1(_17602_),
    .A2(_17633_),
    .B1_N(_17683_),
    .Y(_17684_));
 sky130_fd_sc_hd__a21oi_2 _20959_ (.A1(_17602_),
    .A2(_17633_),
    .B1(_17684_),
    .Y(_03914_));
 sky130_fd_sc_hd__nor2_2 _20960_ (.A(_17604_),
    .B(_17630_),
    .Y(_17685_));
 sky130_fd_sc_hd__buf_1 _20961_ (.A(\count_instr[43] ),
    .X(_17686_));
 sky130_fd_sc_hd__and3_2 _20962_ (.A(_17685_),
    .B(_17686_),
    .C(_17632_),
    .X(_17687_));
 sky130_fd_sc_hd__buf_1 _20963_ (.A(_17147_),
    .X(_17688_));
 sky130_fd_sc_hd__buf_1 _20964_ (.A(_17688_),
    .X(_17689_));
 sky130_fd_sc_hd__a31oi_2 _20965_ (.A1(_17680_),
    .A2(_17681_),
    .A3(_17632_),
    .B1(_17689_),
    .Y(_17690_));
 sky130_fd_sc_hd__o21a_2 _20966_ (.A1(_17681_),
    .A2(_17687_),
    .B1(_17690_),
    .X(_03913_));
 sky130_vsdinv _20967_ (.A(\count_instr[46] ),
    .Y(_17691_));
 sky130_fd_sc_hd__buf_1 _20968_ (.A(\count_instr[44] ),
    .X(_17692_));
 sky130_fd_sc_hd__nand3_2 _20969_ (.A(_17631_),
    .B(\count_instr[45] ),
    .C(_17692_),
    .Y(_17693_));
 sky130_fd_sc_hd__nor3b_2 _20970_ (.A(_17691_),
    .B(_17693_),
    .C_N(\count_instr[47] ),
    .Y(_17694_));
 sky130_fd_sc_hd__nor2_2 _20971_ (.A(_17691_),
    .B(_17693_),
    .Y(_17695_));
 sky130_fd_sc_hd__buf_1 _20972_ (.A(_16931_),
    .X(_17696_));
 sky130_fd_sc_hd__buf_1 _20973_ (.A(_17696_),
    .X(_17697_));
 sky130_fd_sc_hd__o21bai_2 _20974_ (.A1(\count_instr[47] ),
    .A2(_17695_),
    .B1_N(_17697_),
    .Y(_17698_));
 sky130_fd_sc_hd__nor2_2 _20975_ (.A(_17694_),
    .B(_17698_),
    .Y(_03912_));
 sky130_fd_sc_hd__buf_1 _20976_ (.A(_17696_),
    .X(_17699_));
 sky130_fd_sc_hd__buf_1 _20977_ (.A(_17699_),
    .X(_17700_));
 sky130_fd_sc_hd__buf_1 _20978_ (.A(\count_instr[45] ),
    .X(_17701_));
 sky130_fd_sc_hd__buf_1 _20979_ (.A(_17692_),
    .X(_17702_));
 sky130_fd_sc_hd__a31oi_2 _20980_ (.A1(_17680_),
    .A2(_17701_),
    .A3(_17702_),
    .B1(\count_instr[46] ),
    .Y(_17703_));
 sky130_fd_sc_hd__nor3_2 _20981_ (.A(_17700_),
    .B(_17703_),
    .C(_17695_),
    .Y(_03911_));
 sky130_fd_sc_hd__buf_1 _20982_ (.A(_17685_),
    .X(_17704_));
 sky130_fd_sc_hd__a31oi_2 _20983_ (.A1(_17704_),
    .A2(_17692_),
    .A3(_17686_),
    .B1(_17701_),
    .Y(_17705_));
 sky130_fd_sc_hd__and4_2 _20984_ (.A(_17685_),
    .B(_17701_),
    .C(_17692_),
    .D(\count_instr[43] ),
    .X(_17706_));
 sky130_fd_sc_hd__nor3_2 _20985_ (.A(_17700_),
    .B(_17705_),
    .C(_17706_),
    .Y(_03910_));
 sky130_fd_sc_hd__a31oi_2 _20986_ (.A1(_17704_),
    .A2(_17702_),
    .A3(_17686_),
    .B1(_17689_),
    .Y(_17707_));
 sky130_fd_sc_hd__o21a_2 _20987_ (.A1(_17702_),
    .A2(_17680_),
    .B1(_17707_),
    .X(_03909_));
 sky130_vsdinv _20988_ (.A(_17704_),
    .Y(_17708_));
 sky130_fd_sc_hd__o31ai_2 _20989_ (.A1(_17603_),
    .A2(_17604_),
    .A3(_17630_),
    .B1(_17120_),
    .Y(_17709_));
 sky130_fd_sc_hd__a21oi_2 _20990_ (.A1(_17708_),
    .A2(_17603_),
    .B1(_17709_),
    .Y(_03908_));
 sky130_fd_sc_hd__buf_1 _20991_ (.A(\count_instr[41] ),
    .X(_17710_));
 sky130_fd_sc_hd__buf_1 _20992_ (.A(\count_instr[40] ),
    .X(_17711_));
 sky130_fd_sc_hd__a31oi_2 _20993_ (.A1(_17629_),
    .A2(_17710_),
    .A3(_17711_),
    .B1(\count_instr[42] ),
    .Y(_17712_));
 sky130_fd_sc_hd__nor3_2 _20994_ (.A(_17700_),
    .B(_17712_),
    .C(_17704_),
    .Y(_03907_));
 sky130_vsdinv _20995_ (.A(_17711_),
    .Y(_17713_));
 sky130_fd_sc_hd__nor2_2 _20996_ (.A(_17605_),
    .B(_17628_),
    .Y(_17714_));
 sky130_fd_sc_hd__nor3b_2 _20997_ (.A(_17713_),
    .B(_17606_),
    .C_N(_17714_),
    .Y(_17715_));
 sky130_fd_sc_hd__a31oi_2 _20998_ (.A1(_17629_),
    .A2(_17710_),
    .A3(_17711_),
    .B1(_17689_),
    .Y(_17716_));
 sky130_fd_sc_hd__o21a_2 _20999_ (.A1(_17710_),
    .A2(_17715_),
    .B1(_17716_),
    .X(_03906_));
 sky130_vsdinv _21000_ (.A(_17629_),
    .Y(_17717_));
 sky130_fd_sc_hd__buf_1 _21001_ (.A(_16838_),
    .X(_17718_));
 sky130_fd_sc_hd__o41ai_2 _21002_ (.A1(_17713_),
    .A2(_17605_),
    .A3(_17606_),
    .A4(_17628_),
    .B1(_17718_),
    .Y(_17719_));
 sky130_fd_sc_hd__a21oi_2 _21003_ (.A1(_17717_),
    .A2(_17713_),
    .B1(_17719_),
    .Y(_03905_));
 sky130_fd_sc_hd__buf_1 _21004_ (.A(\count_instr[38] ),
    .X(_17720_));
 sky130_fd_sc_hd__and3_2 _21005_ (.A(_17714_),
    .B(\count_instr[39] ),
    .C(_17720_),
    .X(_17721_));
 sky130_vsdinv _21006_ (.A(_17720_),
    .Y(_17722_));
 sky130_fd_sc_hd__nor3_2 _21007_ (.A(_17722_),
    .B(_17605_),
    .C(_17628_),
    .Y(_17723_));
 sky130_fd_sc_hd__o21bai_2 _21008_ (.A1(\count_instr[39] ),
    .A2(_17723_),
    .B1_N(_17697_),
    .Y(_17724_));
 sky130_fd_sc_hd__nor2_2 _21009_ (.A(_17721_),
    .B(_17724_),
    .Y(_03904_));
 sky130_fd_sc_hd__buf_1 _21010_ (.A(_17627_),
    .X(_17725_));
 sky130_fd_sc_hd__buf_1 _21011_ (.A(\count_instr[36] ),
    .X(_17726_));
 sky130_fd_sc_hd__buf_1 _21012_ (.A(\count_instr[35] ),
    .X(_17727_));
 sky130_fd_sc_hd__a41oi_2 _21013_ (.A1(\count_instr[37] ),
    .A2(_17725_),
    .A3(_17726_),
    .A4(_17727_),
    .B1(_17720_),
    .Y(_17728_));
 sky130_fd_sc_hd__nor3_2 _21014_ (.A(_17700_),
    .B(_17728_),
    .C(_17723_),
    .Y(_03903_));
 sky130_fd_sc_hd__buf_1 _21015_ (.A(_17699_),
    .X(_17729_));
 sky130_fd_sc_hd__a31oi_2 _21016_ (.A1(_17725_),
    .A2(_17726_),
    .A3(_17727_),
    .B1(\count_instr[37] ),
    .Y(_17730_));
 sky130_fd_sc_hd__nor3_2 _21017_ (.A(_17729_),
    .B(_17730_),
    .C(_17714_),
    .Y(_03902_));
 sky130_vsdinv _21018_ (.A(\count_instr[35] ),
    .Y(_17731_));
 sky130_fd_sc_hd__buf_1 _21019_ (.A(_17607_),
    .X(_17732_));
 sky130_vsdinv _21020_ (.A(\count_instr[26] ),
    .Y(_17733_));
 sky130_fd_sc_hd__buf_1 _21021_ (.A(_17622_),
    .X(_17734_));
 sky130_fd_sc_hd__nor2_2 _21022_ (.A(_17610_),
    .B(_17734_),
    .Y(_17735_));
 sky130_fd_sc_hd__nand3_2 _21023_ (.A(_17735_),
    .B(\count_instr[25] ),
    .C(\count_instr[24] ),
    .Y(_17736_));
 sky130_fd_sc_hd__nor2_2 _21024_ (.A(_17733_),
    .B(_17736_),
    .Y(_17737_));
 sky130_fd_sc_hd__and3_2 _21025_ (.A(_17737_),
    .B(\count_instr[27] ),
    .C(_17625_),
    .X(_17738_));
 sky130_fd_sc_hd__nand3_2 _21026_ (.A(_17738_),
    .B(\count_instr[33] ),
    .C(\count_instr[32] ),
    .Y(_17739_));
 sky130_fd_sc_hd__nor3_2 _21027_ (.A(_17731_),
    .B(_17732_),
    .C(_17739_),
    .Y(_17740_));
 sky130_fd_sc_hd__a31oi_2 _21028_ (.A1(_17725_),
    .A2(_17726_),
    .A3(_17727_),
    .B1(_17689_),
    .Y(_17741_));
 sky130_fd_sc_hd__o21a_2 _21029_ (.A1(_17726_),
    .A2(_17740_),
    .B1(_17741_),
    .X(_03901_));
 sky130_vsdinv _21030_ (.A(_17725_),
    .Y(_17742_));
 sky130_fd_sc_hd__buf_1 _21031_ (.A(_17608_),
    .X(_17743_));
 sky130_fd_sc_hd__o41ai_2 _21032_ (.A1(_17731_),
    .A2(_17732_),
    .A3(_17743_),
    .A4(_17626_),
    .B1(_17718_),
    .Y(_17744_));
 sky130_fd_sc_hd__a21oi_2 _21033_ (.A1(_17731_),
    .A2(_17742_),
    .B1(_17744_),
    .Y(_03900_));
 sky130_fd_sc_hd__buf_1 _21034_ (.A(_17626_),
    .X(_17745_));
 sky130_fd_sc_hd__o31ai_2 _21035_ (.A1(_17732_),
    .A2(_17743_),
    .A3(_17745_),
    .B1(_17120_),
    .Y(_17746_));
 sky130_fd_sc_hd__a21oi_2 _21036_ (.A1(_17732_),
    .A2(_17739_),
    .B1(_17746_),
    .Y(_03899_));
 sky130_fd_sc_hd__o21bai_2 _21037_ (.A1(_17743_),
    .A2(_17745_),
    .B1_N(_17683_),
    .Y(_17747_));
 sky130_fd_sc_hd__a21oi_2 _21038_ (.A1(_17743_),
    .A2(_17745_),
    .B1(_17747_),
    .Y(_03898_));
 sky130_fd_sc_hd__buf_1 _21039_ (.A(_17696_),
    .X(_17748_));
 sky130_fd_sc_hd__buf_1 _21040_ (.A(_17748_),
    .X(_17749_));
 sky130_fd_sc_hd__buf_1 _21041_ (.A(_17737_),
    .X(_17750_));
 sky130_fd_sc_hd__buf_1 _21042_ (.A(\count_instr[27] ),
    .X(_17751_));
 sky130_fd_sc_hd__a31oi_2 _21043_ (.A1(_17750_),
    .A2(_17751_),
    .A3(_17625_),
    .B1(\count_instr[32] ),
    .Y(_17752_));
 sky130_fd_sc_hd__nor3b_2 _21044_ (.A(_17749_),
    .B(_17752_),
    .C_N(_17745_),
    .Y(_03897_));
 sky130_fd_sc_hd__buf_1 _21045_ (.A(\count_instr[28] ),
    .X(_17753_));
 sky130_fd_sc_hd__and4_2 _21046_ (.A(_17737_),
    .B(\count_instr[29] ),
    .C(_17753_),
    .D(_17751_),
    .X(_17754_));
 sky130_fd_sc_hd__buf_1 _21047_ (.A(\count_instr[30] ),
    .X(_17755_));
 sky130_fd_sc_hd__and3_2 _21048_ (.A(_17754_),
    .B(\count_instr[31] ),
    .C(_17755_),
    .X(_17756_));
 sky130_fd_sc_hd__buf_1 _21049_ (.A(\count_instr[29] ),
    .X(_17757_));
 sky130_fd_sc_hd__and4_2 _21050_ (.A(_17624_),
    .B(_17755_),
    .C(_17757_),
    .D(_17753_),
    .X(_17758_));
 sky130_fd_sc_hd__o21bai_2 _21051_ (.A1(\count_instr[31] ),
    .A2(_17758_),
    .B1_N(_17697_),
    .Y(_17759_));
 sky130_fd_sc_hd__nor2_2 _21052_ (.A(_17756_),
    .B(_17759_),
    .Y(_03896_));
 sky130_fd_sc_hd__buf_1 _21053_ (.A(_17753_),
    .X(_17760_));
 sky130_fd_sc_hd__a31oi_2 _21054_ (.A1(_17624_),
    .A2(_17757_),
    .A3(_17760_),
    .B1(_17755_),
    .Y(_17761_));
 sky130_fd_sc_hd__nor3_2 _21055_ (.A(_17729_),
    .B(_17761_),
    .C(_17758_),
    .Y(_03895_));
 sky130_fd_sc_hd__a31oi_2 _21056_ (.A1(_17750_),
    .A2(_17753_),
    .A3(_17751_),
    .B1(_17757_),
    .Y(_17762_));
 sky130_fd_sc_hd__nor3_2 _21057_ (.A(_17729_),
    .B(_17762_),
    .C(_17754_),
    .Y(_03894_));
 sky130_fd_sc_hd__buf_1 _21058_ (.A(_17751_),
    .X(_17763_));
 sky130_fd_sc_hd__buf_1 _21059_ (.A(_17688_),
    .X(_17764_));
 sky130_fd_sc_hd__a31oi_2 _21060_ (.A1(_17750_),
    .A2(_17760_),
    .A3(_17763_),
    .B1(_17764_),
    .Y(_17765_));
 sky130_fd_sc_hd__o21a_2 _21061_ (.A1(_17760_),
    .A2(_17624_),
    .B1(_17765_),
    .X(_03893_));
 sky130_fd_sc_hd__buf_1 _21062_ (.A(_17623_),
    .X(_17766_));
 sky130_fd_sc_hd__buf_1 _21063_ (.A(\count_instr[26] ),
    .X(_17767_));
 sky130_fd_sc_hd__buf_1 _21064_ (.A(_17147_),
    .X(_17768_));
 sky130_fd_sc_hd__buf_1 _21065_ (.A(_17768_),
    .X(_17769_));
 sky130_fd_sc_hd__a41oi_2 _21066_ (.A1(_17763_),
    .A2(_17766_),
    .A3(_17767_),
    .A4(\count_instr[25] ),
    .B1(_17769_),
    .Y(_17770_));
 sky130_fd_sc_hd__o21a_2 _21067_ (.A1(_17763_),
    .A2(_17750_),
    .B1(_17770_),
    .X(_03892_));
 sky130_vsdinv _21068_ (.A(_17736_),
    .Y(_17771_));
 sky130_fd_sc_hd__buf_1 _21069_ (.A(\count_instr[25] ),
    .X(_17772_));
 sky130_fd_sc_hd__a31oi_2 _21070_ (.A1(_17766_),
    .A2(_17767_),
    .A3(_17772_),
    .B1(_17764_),
    .Y(_17773_));
 sky130_fd_sc_hd__o21a_2 _21071_ (.A1(_17767_),
    .A2(_17771_),
    .B1(_17773_),
    .X(_03891_));
 sky130_fd_sc_hd__a31oi_2 _21072_ (.A1(_17735_),
    .A2(_17772_),
    .A3(\count_instr[24] ),
    .B1(_17764_),
    .Y(_17774_));
 sky130_fd_sc_hd__o21a_2 _21073_ (.A1(_17772_),
    .A2(_17766_),
    .B1(_17774_),
    .X(_03890_));
 sky130_fd_sc_hd__o21a_2 _21074_ (.A1(_17610_),
    .A2(_17734_),
    .B1(_17609_),
    .X(_17775_));
 sky130_fd_sc_hd__nor3_2 _21075_ (.A(_17729_),
    .B(_17766_),
    .C(_17775_),
    .Y(_03889_));
 sky130_vsdinv _21076_ (.A(\count_instr[22] ),
    .Y(_17776_));
 sky130_fd_sc_hd__buf_1 _21077_ (.A(_17734_),
    .X(_17777_));
 sky130_fd_sc_hd__nor3b_2 _21078_ (.A(_17776_),
    .B(_17777_),
    .C_N(\count_instr[23] ),
    .Y(_17778_));
 sky130_fd_sc_hd__nor2_2 _21079_ (.A(_17776_),
    .B(_17734_),
    .Y(_17779_));
 sky130_fd_sc_hd__o21bai_2 _21080_ (.A1(\count_instr[23] ),
    .A2(_17779_),
    .B1_N(_17697_),
    .Y(_17780_));
 sky130_fd_sc_hd__nor2_2 _21081_ (.A(_17778_),
    .B(_17780_),
    .Y(_03888_));
 sky130_fd_sc_hd__o21bai_2 _21082_ (.A1(_17776_),
    .A2(_17777_),
    .B1_N(_17683_),
    .Y(_17781_));
 sky130_fd_sc_hd__a21oi_2 _21083_ (.A1(_17776_),
    .A2(_17777_),
    .B1(_17781_),
    .Y(_03887_));
 sky130_fd_sc_hd__buf_1 _21084_ (.A(_16933_),
    .X(_17782_));
 sky130_fd_sc_hd__buf_1 _21085_ (.A(\count_instr[20] ),
    .X(_17783_));
 sky130_fd_sc_hd__nor3b_2 _21086_ (.A(_17617_),
    .B(_16928_),
    .C_N(\count_instr[13] ),
    .Y(_17784_));
 sky130_fd_sc_hd__buf_1 _21087_ (.A(_17619_),
    .X(_17785_));
 sky130_fd_sc_hd__and4_2 _21088_ (.A(_17784_),
    .B(\count_instr[17] ),
    .C(\count_instr[16] ),
    .D(_17785_),
    .X(_17786_));
 sky130_fd_sc_hd__buf_1 _21089_ (.A(\count_instr[19] ),
    .X(_17787_));
 sky130_fd_sc_hd__a41oi_2 _21090_ (.A1(_17783_),
    .A2(_17786_),
    .A3(_17787_),
    .A4(\count_instr[18] ),
    .B1(\count_instr[21] ),
    .Y(_17788_));
 sky130_fd_sc_hd__nor3b_2 _21091_ (.A(_17782_),
    .B(_17788_),
    .C_N(_17777_),
    .Y(_03886_));
 sky130_fd_sc_hd__buf_1 _21092_ (.A(\count_instr[18] ),
    .X(_17789_));
 sky130_fd_sc_hd__a41oi_2 _21093_ (.A1(_17783_),
    .A2(_17786_),
    .A3(_17787_),
    .A4(_17789_),
    .B1(_17769_),
    .Y(_17790_));
 sky130_fd_sc_hd__o21a_2 _21094_ (.A1(_17783_),
    .A2(_17621_),
    .B1(_17790_),
    .X(_03885_));
 sky130_fd_sc_hd__buf_1 _21095_ (.A(_17699_),
    .X(_17791_));
 sky130_fd_sc_hd__buf_1 _21096_ (.A(\count_instr[17] ),
    .X(_17792_));
 sky130_fd_sc_hd__a31oi_2 _21097_ (.A1(_17620_),
    .A2(\count_instr[18] ),
    .A3(_17792_),
    .B1(_17787_),
    .Y(_17793_));
 sky130_fd_sc_hd__nor3_2 _21098_ (.A(_17791_),
    .B(_17793_),
    .C(_17621_),
    .Y(_03884_));
 sky130_fd_sc_hd__a31oi_2 _21099_ (.A1(_17620_),
    .A2(_17789_),
    .A3(_17792_),
    .B1(_17764_),
    .Y(_17794_));
 sky130_fd_sc_hd__o21a_2 _21100_ (.A1(_17789_),
    .A2(_17786_),
    .B1(_17794_),
    .X(_03883_));
 sky130_fd_sc_hd__buf_1 _21101_ (.A(\count_instr[16] ),
    .X(_17795_));
 sky130_fd_sc_hd__buf_1 _21102_ (.A(_17618_),
    .X(_17796_));
 sky130_fd_sc_hd__buf_1 _21103_ (.A(\count_instr[13] ),
    .X(_17797_));
 sky130_fd_sc_hd__buf_1 _21104_ (.A(_17797_),
    .X(_17798_));
 sky130_fd_sc_hd__a41oi_2 _21105_ (.A1(_17795_),
    .A2(_17796_),
    .A3(_17798_),
    .A4(_17785_),
    .B1(_17792_),
    .Y(_17799_));
 sky130_fd_sc_hd__nor3_2 _21106_ (.A(_17791_),
    .B(_17799_),
    .C(_17786_),
    .Y(_03882_));
 sky130_fd_sc_hd__and3_2 _21107_ (.A(_17796_),
    .B(_17797_),
    .C(_17785_),
    .X(_17800_));
 sky130_fd_sc_hd__a41oi_2 _21108_ (.A1(_17795_),
    .A2(_17796_),
    .A3(_17798_),
    .A4(_17785_),
    .B1(_17769_),
    .Y(_17801_));
 sky130_fd_sc_hd__o21a_2 _21109_ (.A1(_17795_),
    .A2(_17800_),
    .B1(_17801_),
    .X(_03881_));
 sky130_fd_sc_hd__a31o_2 _21110_ (.A1(_17618_),
    .A2(\count_instr[14] ),
    .A3(_17797_),
    .B1(\count_instr[15] ),
    .X(_17802_));
 sky130_fd_sc_hd__buf_1 _21111_ (.A(_16854_),
    .X(_17803_));
 sky130_fd_sc_hd__buf_1 _21112_ (.A(_17803_),
    .X(_17804_));
 sky130_fd_sc_hd__buf_1 _21113_ (.A(\count_instr[14] ),
    .X(_17805_));
 sky130_fd_sc_hd__nand3_2 _21114_ (.A(_17784_),
    .B(\count_instr[15] ),
    .C(_17805_),
    .Y(_17806_));
 sky130_fd_sc_hd__nand3_2 _21115_ (.A(_17802_),
    .B(_17804_),
    .C(_17806_),
    .Y(_17807_));
 sky130_vsdinv _21116_ (.A(_17807_),
    .Y(_03880_));
 sky130_fd_sc_hd__buf_1 _21117_ (.A(_17688_),
    .X(_17808_));
 sky130_fd_sc_hd__a31oi_2 _21118_ (.A1(_17796_),
    .A2(_17805_),
    .A3(_17798_),
    .B1(_17808_),
    .Y(_17809_));
 sky130_fd_sc_hd__o21a_2 _21119_ (.A1(_17805_),
    .A2(_17784_),
    .B1(_17809_),
    .X(_03879_));
 sky130_fd_sc_hd__buf_1 _21120_ (.A(_17337_),
    .X(_17810_));
 sky130_fd_sc_hd__a41oi_2 _21121_ (.A1(_17040_),
    .A2(_16926_),
    .A3(_17810_),
    .A4(_17616_),
    .B1(_17798_),
    .Y(_17811_));
 sky130_fd_sc_hd__nor3_2 _21122_ (.A(_17791_),
    .B(_17811_),
    .C(_17784_),
    .Y(_03878_));
 sky130_fd_sc_hd__buf_1 _21123_ (.A(\count_instr[9] ),
    .X(_17812_));
 sky130_vsdinv _21124_ (.A(_17812_),
    .Y(_17813_));
 sky130_fd_sc_hd__buf_1 _21125_ (.A(\count_instr[0] ),
    .X(_17814_));
 sky130_vsdinv _21126_ (.A(_17814_),
    .Y(_17815_));
 sky130_fd_sc_hd__nor2_2 _21127_ (.A(_17815_),
    .B(_16928_),
    .Y(_17816_));
 sky130_fd_sc_hd__and4_2 _21128_ (.A(_17816_),
    .B(\count_instr[3] ),
    .C(\count_instr[2] ),
    .D(\count_instr[1] ),
    .X(_17817_));
 sky130_fd_sc_hd__buf_1 _21129_ (.A(\count_instr[6] ),
    .X(_17818_));
 sky130_fd_sc_hd__buf_1 _21130_ (.A(\count_instr[4] ),
    .X(_17819_));
 sky130_fd_sc_hd__and4_2 _21131_ (.A(_17817_),
    .B(_17818_),
    .C(\count_instr[5] ),
    .D(_17819_),
    .X(_17820_));
 sky130_fd_sc_hd__nand3_2 _21132_ (.A(_17820_),
    .B(\count_instr[8] ),
    .C(\count_instr[7] ),
    .Y(_17821_));
 sky130_fd_sc_hd__nor2_2 _21133_ (.A(_17813_),
    .B(_17821_),
    .Y(_17822_));
 sky130_fd_sc_hd__buf_1 _21134_ (.A(\count_instr[10] ),
    .X(_17823_));
 sky130_fd_sc_hd__a31o_2 _21135_ (.A1(_17822_),
    .A2(\count_instr[11] ),
    .A3(_17823_),
    .B1(\count_instr[12] ),
    .X(_17824_));
 sky130_fd_sc_hd__nor3b_2 _21136_ (.A(_17813_),
    .B(_17821_),
    .C_N(\count_instr[10] ),
    .Y(_17825_));
 sky130_fd_sc_hd__buf_1 _21137_ (.A(\count_instr[11] ),
    .X(_17826_));
 sky130_fd_sc_hd__nand3_2 _21138_ (.A(_17825_),
    .B(\count_instr[12] ),
    .C(_17826_),
    .Y(_17827_));
 sky130_fd_sc_hd__nand3_2 _21139_ (.A(_17824_),
    .B(_17718_),
    .C(_17827_),
    .Y(_17828_));
 sky130_vsdinv _21140_ (.A(_17828_),
    .Y(_03877_));
 sky130_fd_sc_hd__a31oi_2 _21141_ (.A1(_17822_),
    .A2(_17826_),
    .A3(_17823_),
    .B1(_17808_),
    .Y(_17829_));
 sky130_fd_sc_hd__o21a_2 _21142_ (.A1(_17826_),
    .A2(_17825_),
    .B1(_17829_),
    .X(_03876_));
 sky130_fd_sc_hd__buf_1 _21143_ (.A(\count_instr[8] ),
    .X(_17830_));
 sky130_fd_sc_hd__buf_1 _21144_ (.A(\count_instr[7] ),
    .X(_17831_));
 sky130_fd_sc_hd__a41oi_2 _21145_ (.A1(_17812_),
    .A2(_17820_),
    .A3(_17830_),
    .A4(_17831_),
    .B1(_17823_),
    .Y(_17832_));
 sky130_fd_sc_hd__nor3_2 _21146_ (.A(_17791_),
    .B(_17832_),
    .C(_17825_),
    .Y(_03875_));
 sky130_fd_sc_hd__buf_1 _21147_ (.A(_17699_),
    .X(_17833_));
 sky130_fd_sc_hd__buf_1 _21148_ (.A(_17820_),
    .X(_17834_));
 sky130_fd_sc_hd__a31oi_2 _21149_ (.A1(_17834_),
    .A2(_17830_),
    .A3(_17831_),
    .B1(_17812_),
    .Y(_17835_));
 sky130_fd_sc_hd__nor3_2 _21150_ (.A(_17833_),
    .B(_17835_),
    .C(_17822_),
    .Y(_03874_));
 sky130_fd_sc_hd__and2_2 _21151_ (.A(_17820_),
    .B(_17831_),
    .X(_17836_));
 sky130_fd_sc_hd__buf_1 _21152_ (.A(_17831_),
    .X(_17837_));
 sky130_fd_sc_hd__a31oi_2 _21153_ (.A1(_17834_),
    .A2(_17830_),
    .A3(_17837_),
    .B1(_17808_),
    .Y(_17838_));
 sky130_fd_sc_hd__o21a_2 _21154_ (.A1(_17830_),
    .A2(_17836_),
    .B1(_17838_),
    .X(_03873_));
 sky130_fd_sc_hd__a21oi_2 _21155_ (.A1(_17834_),
    .A2(_17837_),
    .B1(_17197_),
    .Y(_17839_));
 sky130_fd_sc_hd__o21a_2 _21156_ (.A1(_17837_),
    .A2(_17834_),
    .B1(_17839_),
    .X(_03872_));
 sky130_fd_sc_hd__buf_1 _21157_ (.A(\count_instr[5] ),
    .X(_17840_));
 sky130_fd_sc_hd__and3_2 _21158_ (.A(_17817_),
    .B(_17840_),
    .C(_17819_),
    .X(_17841_));
 sky130_fd_sc_hd__a41oi_2 _21159_ (.A1(_17818_),
    .A2(_17817_),
    .A3(_17840_),
    .A4(_17819_),
    .B1(_17769_),
    .Y(_17842_));
 sky130_fd_sc_hd__o21a_2 _21160_ (.A1(_17818_),
    .A2(_17841_),
    .B1(_17842_),
    .X(_03871_));
 sky130_fd_sc_hd__buf_1 _21161_ (.A(_17817_),
    .X(_17843_));
 sky130_fd_sc_hd__buf_1 _21162_ (.A(_17819_),
    .X(_17844_));
 sky130_fd_sc_hd__a21oi_2 _21163_ (.A1(_17843_),
    .A2(_17844_),
    .B1(_17840_),
    .Y(_17845_));
 sky130_fd_sc_hd__nor3_2 _21164_ (.A(_17833_),
    .B(_17845_),
    .C(_17841_),
    .Y(_03870_));
 sky130_fd_sc_hd__a21oi_2 _21165_ (.A1(_17843_),
    .A2(_17844_),
    .B1(_17197_),
    .Y(_17846_));
 sky130_fd_sc_hd__o21a_2 _21166_ (.A1(_17844_),
    .A2(_17843_),
    .B1(_17846_),
    .X(_03869_));
 sky130_fd_sc_hd__buf_1 _21167_ (.A(\count_instr[2] ),
    .X(_17847_));
 sky130_fd_sc_hd__buf_1 _21168_ (.A(\count_instr[1] ),
    .X(_17848_));
 sky130_fd_sc_hd__a31oi_2 _21169_ (.A1(_17816_),
    .A2(_17847_),
    .A3(_17848_),
    .B1(\count_instr[3] ),
    .Y(_17849_));
 sky130_fd_sc_hd__nor3_2 _21170_ (.A(_17833_),
    .B(_17849_),
    .C(_17843_),
    .Y(_03868_));
 sky130_fd_sc_hd__nor3b_2 _21171_ (.A(_17815_),
    .B(_16929_),
    .C_N(_17848_),
    .Y(_17850_));
 sky130_fd_sc_hd__buf_1 _21172_ (.A(_17451_),
    .X(_17851_));
 sky130_fd_sc_hd__buf_1 _21173_ (.A(_17851_),
    .X(_17852_));
 sky130_fd_sc_hd__and3_2 _21174_ (.A(_17816_),
    .B(_17847_),
    .C(\count_instr[1] ),
    .X(_17853_));
 sky130_vsdinv _21175_ (.A(_17853_),
    .Y(_17854_));
 sky130_fd_sc_hd__o211a_2 _21176_ (.A1(_17847_),
    .A2(_17850_),
    .B1(_17852_),
    .C1(_17854_),
    .X(_03867_));
 sky130_fd_sc_hd__a41oi_2 _21177_ (.A1(_17040_),
    .A2(_16926_),
    .A3(_17814_),
    .A4(_17810_),
    .B1(_17848_),
    .Y(_17855_));
 sky130_fd_sc_hd__nor3_2 _21178_ (.A(_17833_),
    .B(_17855_),
    .C(_17850_),
    .Y(_03866_));
 sky130_fd_sc_hd__buf_1 _21179_ (.A(_17696_),
    .X(_17856_));
 sky130_fd_sc_hd__buf_1 _21180_ (.A(_17856_),
    .X(_17857_));
 sky130_fd_sc_hd__a31oi_2 _21181_ (.A1(_16926_),
    .A2(_17040_),
    .A3(_17810_),
    .B1(_17814_),
    .Y(_17858_));
 sky130_fd_sc_hd__nor3_2 _21182_ (.A(_17857_),
    .B(_17858_),
    .C(_17816_),
    .Y(_03865_));
 sky130_fd_sc_hd__buf_1 _21183_ (.A(_16829_),
    .X(_17859_));
 sky130_fd_sc_hd__buf_1 _21184_ (.A(_17859_),
    .X(_17860_));
 sky130_fd_sc_hd__buf_1 _21185_ (.A(\irq_pending[31] ),
    .X(_17861_));
 sky130_fd_sc_hd__nor3b_2 _21186_ (.A(_17088_),
    .B(_17860_),
    .C_N(_17861_),
    .Y(_17862_));
 sky130_fd_sc_hd__nor2_2 _21187_ (.A(_17025_),
    .B(\cpu_state[2] ),
    .Y(_00315_));
 sky130_fd_sc_hd__and2b_2 _21188_ (.A_N(_17033_),
    .B(_17025_),
    .X(_17863_));
 sky130_fd_sc_hd__a211o_2 _21189_ (.A1(_17007_),
    .A2(_17019_),
    .B1(_00315_),
    .C1(_17863_),
    .X(_17864_));
 sky130_fd_sc_hd__buf_1 _21190_ (.A(_17864_),
    .X(_17865_));
 sky130_fd_sc_hd__buf_1 _21191_ (.A(_17865_),
    .X(_17866_));
 sky130_fd_sc_hd__buf_1 _21192_ (.A(_17864_),
    .X(_17867_));
 sky130_fd_sc_hd__buf_1 _21193_ (.A(_17867_),
    .X(_17868_));
 sky130_fd_sc_hd__or2b_2 _21194_ (.A(eoi[31]),
    .B_N(_17868_),
    .X(_17869_));
 sky130_fd_sc_hd__o211a_2 _21195_ (.A1(_17862_),
    .A2(_17866_),
    .B1(_17852_),
    .C1(_17869_),
    .X(_03864_));
 sky130_fd_sc_hd__buf_1 _21196_ (.A(\irq_pending[30] ),
    .X(_17870_));
 sky130_fd_sc_hd__nor3b_2 _21197_ (.A(_17108_),
    .B(_17860_),
    .C_N(_17870_),
    .Y(_17871_));
 sky130_fd_sc_hd__or2b_2 _21198_ (.A(eoi[30]),
    .B_N(_17868_),
    .X(_17872_));
 sky130_fd_sc_hd__o211a_2 _21199_ (.A1(_17871_),
    .A2(_17866_),
    .B1(_17852_),
    .C1(_17872_),
    .X(_03863_));
 sky130_fd_sc_hd__buf_1 _21200_ (.A(\irq_pending[29] ),
    .X(_17873_));
 sky130_fd_sc_hd__nor3b_2 _21201_ (.A(_17113_),
    .B(_17860_),
    .C_N(_17873_),
    .Y(_17874_));
 sky130_fd_sc_hd__or2b_2 _21202_ (.A(eoi[29]),
    .B_N(_17868_),
    .X(_17875_));
 sky130_fd_sc_hd__o211a_2 _21203_ (.A1(_17874_),
    .A2(_17866_),
    .B1(_17852_),
    .C1(_17875_),
    .X(_03862_));
 sky130_fd_sc_hd__buf_1 _21204_ (.A(\irq_pending[28] ),
    .X(_17876_));
 sky130_fd_sc_hd__nor3b_2 _21205_ (.A(_17116_),
    .B(_17860_),
    .C_N(_17876_),
    .Y(_17877_));
 sky130_fd_sc_hd__buf_1 _21206_ (.A(_17851_),
    .X(_17878_));
 sky130_fd_sc_hd__or2b_2 _21207_ (.A(eoi[28]),
    .B_N(_17868_),
    .X(_17879_));
 sky130_fd_sc_hd__o211a_2 _21208_ (.A1(_17877_),
    .A2(_17866_),
    .B1(_17878_),
    .C1(_17879_),
    .X(_03861_));
 sky130_fd_sc_hd__buf_1 _21209_ (.A(_17859_),
    .X(_17880_));
 sky130_fd_sc_hd__buf_1 _21210_ (.A(\irq_pending[27] ),
    .X(_17881_));
 sky130_fd_sc_hd__nor3b_2 _21211_ (.A(\irq_mask[27] ),
    .B(_17880_),
    .C_N(_17881_),
    .Y(_17882_));
 sky130_fd_sc_hd__buf_1 _21212_ (.A(_17865_),
    .X(_17883_));
 sky130_fd_sc_hd__buf_1 _21213_ (.A(_17867_),
    .X(_17884_));
 sky130_fd_sc_hd__or2b_2 _21214_ (.A(eoi[27]),
    .B_N(_17884_),
    .X(_17885_));
 sky130_fd_sc_hd__o211a_2 _21215_ (.A1(_17882_),
    .A2(_17883_),
    .B1(_17878_),
    .C1(_17885_),
    .X(_03860_));
 sky130_fd_sc_hd__buf_1 _21216_ (.A(\irq_pending[26] ),
    .X(_17886_));
 sky130_fd_sc_hd__nor3b_2 _21217_ (.A(_17126_),
    .B(_17880_),
    .C_N(_17886_),
    .Y(_17887_));
 sky130_fd_sc_hd__or2b_2 _21218_ (.A(eoi[26]),
    .B_N(_17884_),
    .X(_17888_));
 sky130_fd_sc_hd__o211a_2 _21219_ (.A1(_17887_),
    .A2(_17883_),
    .B1(_17878_),
    .C1(_17888_),
    .X(_03859_));
 sky130_fd_sc_hd__buf_1 _21220_ (.A(\irq_pending[25] ),
    .X(_17889_));
 sky130_fd_sc_hd__nor3b_2 _21221_ (.A(_17129_),
    .B(_17880_),
    .C_N(_17889_),
    .Y(_17890_));
 sky130_fd_sc_hd__or2b_2 _21222_ (.A(eoi[25]),
    .B_N(_17884_),
    .X(_17891_));
 sky130_fd_sc_hd__o211a_2 _21223_ (.A1(_17890_),
    .A2(_17883_),
    .B1(_17878_),
    .C1(_17891_),
    .X(_03858_));
 sky130_fd_sc_hd__buf_1 _21224_ (.A(\irq_pending[24] ),
    .X(_17892_));
 sky130_fd_sc_hd__nor3b_2 _21225_ (.A(_17134_),
    .B(_17880_),
    .C_N(_17892_),
    .Y(_17893_));
 sky130_fd_sc_hd__buf_1 _21226_ (.A(_17851_),
    .X(_17894_));
 sky130_fd_sc_hd__or2b_2 _21227_ (.A(eoi[24]),
    .B_N(_17884_),
    .X(_17895_));
 sky130_fd_sc_hd__o211a_2 _21228_ (.A1(_17893_),
    .A2(_17883_),
    .B1(_17894_),
    .C1(_17895_),
    .X(_03857_));
 sky130_fd_sc_hd__buf_1 _21229_ (.A(\irq_mask[23] ),
    .X(_17896_));
 sky130_fd_sc_hd__buf_1 _21230_ (.A(_16829_),
    .X(_17897_));
 sky130_fd_sc_hd__buf_1 _21231_ (.A(_17897_),
    .X(_17898_));
 sky130_fd_sc_hd__buf_1 _21232_ (.A(\irq_pending[23] ),
    .X(_17899_));
 sky130_fd_sc_hd__nor3b_2 _21233_ (.A(_17896_),
    .B(_17898_),
    .C_N(_17899_),
    .Y(_17900_));
 sky130_fd_sc_hd__buf_1 _21234_ (.A(_17865_),
    .X(_17901_));
 sky130_fd_sc_hd__buf_1 _21235_ (.A(_17867_),
    .X(_17902_));
 sky130_fd_sc_hd__or2b_2 _21236_ (.A(eoi[23]),
    .B_N(_17902_),
    .X(_17903_));
 sky130_fd_sc_hd__o211a_2 _21237_ (.A1(_17900_),
    .A2(_17901_),
    .B1(_17894_),
    .C1(_17903_),
    .X(_03856_));
 sky130_fd_sc_hd__buf_1 _21238_ (.A(\irq_pending[22] ),
    .X(_17904_));
 sky130_fd_sc_hd__nor3b_2 _21239_ (.A(_17143_),
    .B(_17898_),
    .C_N(_17904_),
    .Y(_17905_));
 sky130_fd_sc_hd__or2b_2 _21240_ (.A(eoi[22]),
    .B_N(_17902_),
    .X(_17906_));
 sky130_fd_sc_hd__o211a_2 _21241_ (.A1(_17905_),
    .A2(_17901_),
    .B1(_17894_),
    .C1(_17906_),
    .X(_03855_));
 sky130_fd_sc_hd__buf_1 _21242_ (.A(\irq_pending[21] ),
    .X(_17907_));
 sky130_fd_sc_hd__nor3b_2 _21243_ (.A(_17146_),
    .B(_17898_),
    .C_N(_17907_),
    .Y(_17908_));
 sky130_fd_sc_hd__or2b_2 _21244_ (.A(eoi[21]),
    .B_N(_17902_),
    .X(_17909_));
 sky130_fd_sc_hd__o211a_2 _21245_ (.A1(_17908_),
    .A2(_17901_),
    .B1(_17894_),
    .C1(_17909_),
    .X(_03854_));
 sky130_fd_sc_hd__buf_1 _21246_ (.A(\irq_pending[20] ),
    .X(_17910_));
 sky130_fd_sc_hd__nor3b_2 _21247_ (.A(_17151_),
    .B(_17898_),
    .C_N(_17910_),
    .Y(_17911_));
 sky130_fd_sc_hd__buf_1 _21248_ (.A(_17851_),
    .X(_17912_));
 sky130_fd_sc_hd__or2b_2 _21249_ (.A(eoi[20]),
    .B_N(_17902_),
    .X(_17913_));
 sky130_fd_sc_hd__o211a_2 _21250_ (.A1(_17911_),
    .A2(_17901_),
    .B1(_17912_),
    .C1(_17913_),
    .X(_03853_));
 sky130_fd_sc_hd__buf_1 _21251_ (.A(_17897_),
    .X(_17914_));
 sky130_fd_sc_hd__buf_1 _21252_ (.A(\irq_pending[19] ),
    .X(_17915_));
 sky130_fd_sc_hd__nor3b_2 _21253_ (.A(_17154_),
    .B(_17914_),
    .C_N(_17915_),
    .Y(_17916_));
 sky130_fd_sc_hd__buf_1 _21254_ (.A(_17865_),
    .X(_17917_));
 sky130_fd_sc_hd__buf_1 _21255_ (.A(_17867_),
    .X(_17918_));
 sky130_fd_sc_hd__or2b_2 _21256_ (.A(eoi[19]),
    .B_N(_17918_),
    .X(_17919_));
 sky130_fd_sc_hd__o211a_2 _21257_ (.A1(_17916_),
    .A2(_17917_),
    .B1(_17912_),
    .C1(_17919_),
    .X(_03852_));
 sky130_fd_sc_hd__buf_1 _21258_ (.A(\irq_pending[18] ),
    .X(_17920_));
 sky130_fd_sc_hd__nor3b_2 _21259_ (.A(_17157_),
    .B(_17914_),
    .C_N(_17920_),
    .Y(_17921_));
 sky130_fd_sc_hd__or2b_2 _21260_ (.A(eoi[18]),
    .B_N(_17918_),
    .X(_17922_));
 sky130_fd_sc_hd__o211a_2 _21261_ (.A1(_17921_),
    .A2(_17917_),
    .B1(_17912_),
    .C1(_17922_),
    .X(_03851_));
 sky130_fd_sc_hd__buf_1 _21262_ (.A(\irq_pending[17] ),
    .X(_17923_));
 sky130_fd_sc_hd__nor3b_2 _21263_ (.A(_17159_),
    .B(_17914_),
    .C_N(_17923_),
    .Y(_17924_));
 sky130_fd_sc_hd__or2b_2 _21264_ (.A(eoi[17]),
    .B_N(_17918_),
    .X(_17925_));
 sky130_fd_sc_hd__o211a_2 _21265_ (.A1(_17924_),
    .A2(_17917_),
    .B1(_17912_),
    .C1(_17925_),
    .X(_03850_));
 sky130_fd_sc_hd__buf_1 _21266_ (.A(\irq_pending[16] ),
    .X(_17926_));
 sky130_fd_sc_hd__nor3b_2 _21267_ (.A(_17162_),
    .B(_17914_),
    .C_N(_17926_),
    .Y(_17927_));
 sky130_fd_sc_hd__buf_1 _21268_ (.A(_17451_),
    .X(_17928_));
 sky130_fd_sc_hd__buf_1 _21269_ (.A(_17928_),
    .X(_17929_));
 sky130_fd_sc_hd__or2b_2 _21270_ (.A(eoi[16]),
    .B_N(_17918_),
    .X(_17930_));
 sky130_fd_sc_hd__o211a_2 _21271_ (.A1(_17927_),
    .A2(_17917_),
    .B1(_17929_),
    .C1(_17930_),
    .X(_03849_));
 sky130_fd_sc_hd__buf_1 _21272_ (.A(\irq_mask[15] ),
    .X(_17931_));
 sky130_fd_sc_hd__buf_1 _21273_ (.A(_17897_),
    .X(_17932_));
 sky130_fd_sc_hd__buf_1 _21274_ (.A(\irq_pending[15] ),
    .X(_17933_));
 sky130_fd_sc_hd__nor3b_2 _21275_ (.A(_17931_),
    .B(_17932_),
    .C_N(_17933_),
    .Y(_17934_));
 sky130_fd_sc_hd__buf_1 _21276_ (.A(_17864_),
    .X(_17935_));
 sky130_fd_sc_hd__buf_1 _21277_ (.A(_17935_),
    .X(_17936_));
 sky130_fd_sc_hd__buf_1 _21278_ (.A(_17864_),
    .X(_17937_));
 sky130_fd_sc_hd__buf_1 _21279_ (.A(_17937_),
    .X(_17938_));
 sky130_fd_sc_hd__or2b_2 _21280_ (.A(eoi[15]),
    .B_N(_17938_),
    .X(_17939_));
 sky130_fd_sc_hd__o211a_2 _21281_ (.A1(_17934_),
    .A2(_17936_),
    .B1(_17929_),
    .C1(_17939_),
    .X(_03848_));
 sky130_fd_sc_hd__buf_1 _21282_ (.A(\irq_pending[14] ),
    .X(_17940_));
 sky130_fd_sc_hd__nor3b_2 _21283_ (.A(_17166_),
    .B(_17932_),
    .C_N(_17940_),
    .Y(_17941_));
 sky130_fd_sc_hd__or2b_2 _21284_ (.A(eoi[14]),
    .B_N(_17938_),
    .X(_17942_));
 sky130_fd_sc_hd__o211a_2 _21285_ (.A1(_17941_),
    .A2(_17936_),
    .B1(_17929_),
    .C1(_17942_),
    .X(_03847_));
 sky130_fd_sc_hd__buf_1 _21286_ (.A(\irq_pending[13] ),
    .X(_17943_));
 sky130_fd_sc_hd__nor3b_2 _21287_ (.A(_17170_),
    .B(_17932_),
    .C_N(_17943_),
    .Y(_17944_));
 sky130_fd_sc_hd__or2b_2 _21288_ (.A(eoi[13]),
    .B_N(_17938_),
    .X(_17945_));
 sky130_fd_sc_hd__o211a_2 _21289_ (.A1(_17944_),
    .A2(_17936_),
    .B1(_17929_),
    .C1(_17945_),
    .X(_03846_));
 sky130_fd_sc_hd__buf_1 _21290_ (.A(\irq_pending[12] ),
    .X(_17946_));
 sky130_fd_sc_hd__nor3b_2 _21291_ (.A(_17176_),
    .B(_17932_),
    .C_N(_17946_),
    .Y(_17947_));
 sky130_fd_sc_hd__buf_1 _21292_ (.A(_17928_),
    .X(_17948_));
 sky130_fd_sc_hd__or2b_2 _21293_ (.A(eoi[12]),
    .B_N(_17938_),
    .X(_17949_));
 sky130_fd_sc_hd__o211a_2 _21294_ (.A1(_17947_),
    .A2(_17936_),
    .B1(_17948_),
    .C1(_17949_),
    .X(_03845_));
 sky130_fd_sc_hd__buf_1 _21295_ (.A(_17897_),
    .X(_17950_));
 sky130_fd_sc_hd__buf_1 _21296_ (.A(\irq_pending[11] ),
    .X(_17951_));
 sky130_fd_sc_hd__nor3b_2 _21297_ (.A(\irq_mask[11] ),
    .B(_17950_),
    .C_N(_17951_),
    .Y(_17952_));
 sky130_fd_sc_hd__buf_1 _21298_ (.A(_17935_),
    .X(_17953_));
 sky130_fd_sc_hd__buf_1 _21299_ (.A(_17937_),
    .X(_17954_));
 sky130_fd_sc_hd__or2b_2 _21300_ (.A(eoi[11]),
    .B_N(_17954_),
    .X(_17955_));
 sky130_fd_sc_hd__o211a_2 _21301_ (.A1(_17952_),
    .A2(_17953_),
    .B1(_17948_),
    .C1(_17955_),
    .X(_03844_));
 sky130_fd_sc_hd__buf_1 _21302_ (.A(\irq_pending[10] ),
    .X(_17956_));
 sky130_fd_sc_hd__nor3b_2 _21303_ (.A(_17180_),
    .B(_17950_),
    .C_N(_17956_),
    .Y(_17957_));
 sky130_fd_sc_hd__or2b_2 _21304_ (.A(eoi[10]),
    .B_N(_17954_),
    .X(_17958_));
 sky130_fd_sc_hd__o211a_2 _21305_ (.A1(_17957_),
    .A2(_17953_),
    .B1(_17948_),
    .C1(_17958_),
    .X(_03843_));
 sky130_fd_sc_hd__buf_1 _21306_ (.A(\irq_pending[9] ),
    .X(_17959_));
 sky130_fd_sc_hd__nor3b_2 _21307_ (.A(_17183_),
    .B(_17950_),
    .C_N(_17959_),
    .Y(_17960_));
 sky130_fd_sc_hd__or2b_2 _21308_ (.A(eoi[9]),
    .B_N(_17954_),
    .X(_17961_));
 sky130_fd_sc_hd__o211a_2 _21309_ (.A1(_17960_),
    .A2(_17953_),
    .B1(_17948_),
    .C1(_17961_),
    .X(_03842_));
 sky130_fd_sc_hd__buf_1 _21310_ (.A(\irq_pending[8] ),
    .X(_17962_));
 sky130_fd_sc_hd__nor3b_2 _21311_ (.A(_17187_),
    .B(_17950_),
    .C_N(_17962_),
    .Y(_17963_));
 sky130_fd_sc_hd__buf_1 _21312_ (.A(_17928_),
    .X(_17964_));
 sky130_fd_sc_hd__or2b_2 _21313_ (.A(eoi[8]),
    .B_N(_17954_),
    .X(_17965_));
 sky130_fd_sc_hd__o211a_2 _21314_ (.A1(_17963_),
    .A2(_17953_),
    .B1(_17964_),
    .C1(_17965_),
    .X(_03841_));
 sky130_fd_sc_hd__buf_1 _21315_ (.A(_16828_),
    .X(_17966_));
 sky130_fd_sc_hd__buf_1 _21316_ (.A(_17966_),
    .X(_17967_));
 sky130_fd_sc_hd__buf_1 _21317_ (.A(\irq_pending[7] ),
    .X(_17968_));
 sky130_fd_sc_hd__nor3b_2 _21318_ (.A(\irq_mask[7] ),
    .B(_17967_),
    .C_N(_17968_),
    .Y(_17969_));
 sky130_fd_sc_hd__buf_1 _21319_ (.A(_17935_),
    .X(_17970_));
 sky130_fd_sc_hd__buf_1 _21320_ (.A(_17937_),
    .X(_17971_));
 sky130_fd_sc_hd__or2b_2 _21321_ (.A(eoi[7]),
    .B_N(_17971_),
    .X(_17972_));
 sky130_fd_sc_hd__o211a_2 _21322_ (.A1(_17969_),
    .A2(_17970_),
    .B1(_17964_),
    .C1(_17972_),
    .X(_03840_));
 sky130_fd_sc_hd__buf_1 _21323_ (.A(\irq_pending[6] ),
    .X(_17973_));
 sky130_fd_sc_hd__nor3b_2 _21324_ (.A(_17196_),
    .B(_17967_),
    .C_N(_17973_),
    .Y(_17974_));
 sky130_fd_sc_hd__or2b_2 _21325_ (.A(eoi[6]),
    .B_N(_17971_),
    .X(_17975_));
 sky130_fd_sc_hd__o211a_2 _21326_ (.A1(_17974_),
    .A2(_17970_),
    .B1(_17964_),
    .C1(_17975_),
    .X(_03839_));
 sky130_fd_sc_hd__buf_1 _21327_ (.A(\irq_pending[5] ),
    .X(_17976_));
 sky130_fd_sc_hd__nor3b_2 _21328_ (.A(_17199_),
    .B(_17967_),
    .C_N(_17976_),
    .Y(_17977_));
 sky130_fd_sc_hd__or2b_2 _21329_ (.A(eoi[5]),
    .B_N(_17971_),
    .X(_17978_));
 sky130_fd_sc_hd__o211a_2 _21330_ (.A1(_17977_),
    .A2(_17970_),
    .B1(_17964_),
    .C1(_17978_),
    .X(_03838_));
 sky130_fd_sc_hd__buf_1 _21331_ (.A(\irq_pending[4] ),
    .X(_17979_));
 sky130_fd_sc_hd__nor3b_2 _21332_ (.A(_17202_),
    .B(_17967_),
    .C_N(_17979_),
    .Y(_17980_));
 sky130_fd_sc_hd__buf_1 _21333_ (.A(_17928_),
    .X(_17981_));
 sky130_fd_sc_hd__or2b_2 _21334_ (.A(eoi[4]),
    .B_N(_17971_),
    .X(_17982_));
 sky130_fd_sc_hd__o211a_2 _21335_ (.A1(_17980_),
    .A2(_17970_),
    .B1(_17981_),
    .C1(_17982_),
    .X(_03837_));
 sky130_fd_sc_hd__buf_1 _21336_ (.A(_17966_),
    .X(_17983_));
 sky130_fd_sc_hd__buf_1 _21337_ (.A(\irq_pending[3] ),
    .X(_17984_));
 sky130_fd_sc_hd__nor3b_2 _21338_ (.A(_17205_),
    .B(_17983_),
    .C_N(_17984_),
    .Y(_17985_));
 sky130_fd_sc_hd__buf_1 _21339_ (.A(_17935_),
    .X(_17986_));
 sky130_fd_sc_hd__buf_1 _21340_ (.A(_17937_),
    .X(_17987_));
 sky130_fd_sc_hd__or2b_2 _21341_ (.A(eoi[3]),
    .B_N(_17987_),
    .X(_17988_));
 sky130_fd_sc_hd__o211a_2 _21342_ (.A1(_17985_),
    .A2(_17986_),
    .B1(_17981_),
    .C1(_17988_),
    .X(_03836_));
 sky130_fd_sc_hd__buf_1 _21343_ (.A(\irq_mask[2] ),
    .X(_17989_));
 sky130_fd_sc_hd__buf_1 _21344_ (.A(_17989_),
    .X(_17990_));
 sky130_fd_sc_hd__buf_1 _21345_ (.A(\irq_pending[2] ),
    .X(_17991_));
 sky130_fd_sc_hd__nor3b_2 _21346_ (.A(_17990_),
    .B(_17983_),
    .C_N(_17991_),
    .Y(_17992_));
 sky130_fd_sc_hd__or2b_2 _21347_ (.A(eoi[2]),
    .B_N(_17987_),
    .X(_17993_));
 sky130_fd_sc_hd__o211a_2 _21348_ (.A1(_17992_),
    .A2(_17986_),
    .B1(_17981_),
    .C1(_17993_),
    .X(_03835_));
 sky130_fd_sc_hd__buf_1 _21349_ (.A(\irq_pending[1] ),
    .X(_17994_));
 sky130_fd_sc_hd__nor3b_2 _21350_ (.A(_17210_),
    .B(_17983_),
    .C_N(_17994_),
    .Y(_17995_));
 sky130_fd_sc_hd__or2b_2 _21351_ (.A(eoi[1]),
    .B_N(_17987_),
    .X(_17996_));
 sky130_fd_sc_hd__o211a_2 _21352_ (.A1(_17995_),
    .A2(_17986_),
    .B1(_17981_),
    .C1(_17996_),
    .X(_03834_));
 sky130_fd_sc_hd__nor3b_2 _21353_ (.A(_17214_),
    .B(_17983_),
    .C_N(\irq_pending[0] ),
    .Y(_17997_));
 sky130_fd_sc_hd__buf_1 _21354_ (.A(_16838_),
    .X(_17998_));
 sky130_fd_sc_hd__or2b_2 _21355_ (.A(eoi[0]),
    .B_N(_17987_),
    .X(_17999_));
 sky130_fd_sc_hd__o211a_2 _21356_ (.A1(_17997_),
    .A2(_17986_),
    .B1(_17998_),
    .C1(_17999_),
    .X(_03833_));
 sky130_fd_sc_hd__nand3_2 _21357_ (.A(_17003_),
    .B(_17017_),
    .C(_17014_),
    .Y(_18000_));
 sky130_fd_sc_hd__buf_1 _21358_ (.A(_17189_),
    .X(_18001_));
 sky130_fd_sc_hd__nor2_2 _21359_ (.A(instr_ecall_ebreak),
    .B(pcpi_timeout),
    .Y(_00311_));
 sky130_vsdinv _21360_ (.A(_00311_),
    .Y(_18002_));
 sky130_fd_sc_hd__buf_1 _21361_ (.A(_17065_),
    .X(_18003_));
 sky130_fd_sc_hd__o2111a_2 _21362_ (.A1(\pcpi_mul.active[1] ),
    .A2(_18002_),
    .B1(_18003_),
    .C1(_17015_),
    .D1(_17004_),
    .X(_18004_));
 sky130_fd_sc_hd__a211oi_2 _21363_ (.A1(_17379_),
    .A2(_18000_),
    .B1(_18001_),
    .C1(_18004_),
    .Y(_03832_));
 sky130_fd_sc_hd__buf_1 _21364_ (.A(mem_valid),
    .X(_18005_));
 sky130_fd_sc_hd__o21bai_2 _21365_ (.A1(_18005_),
    .A2(_16850_),
    .B1_N(_16802_),
    .Y(_18006_));
 sky130_fd_sc_hd__nand3_2 _21366_ (.A(_16835_),
    .B(_16844_),
    .C(_18005_),
    .Y(_18007_));
 sky130_fd_sc_hd__a21o_2 _21367_ (.A1(_18006_),
    .A2(_18007_),
    .B1(_16836_),
    .X(_18008_));
 sky130_fd_sc_hd__or2b_2 _21368_ (.A(_16800_),
    .B_N(_18005_),
    .X(_18009_));
 sky130_fd_sc_hd__a21oi_2 _21369_ (.A1(_18008_),
    .A2(_18009_),
    .B1(_17370_),
    .Y(_03831_));
 sky130_fd_sc_hd__or4_2 _21370_ (.A(_17907_),
    .B(_17910_),
    .C(\irq_pending[23] ),
    .D(_17904_),
    .X(_18010_));
 sky130_fd_sc_hd__or4_2 _21371_ (.A(_17923_),
    .B(_17926_),
    .C(_17915_),
    .D(_17920_),
    .X(_18011_));
 sky130_fd_sc_hd__or4_2 _21372_ (.A(_17873_),
    .B(_17876_),
    .C(_17861_),
    .D(_17870_),
    .X(_18012_));
 sky130_fd_sc_hd__or4_2 _21373_ (.A(_17889_),
    .B(_17892_),
    .C(\irq_pending[27] ),
    .D(_17886_),
    .X(_18013_));
 sky130_fd_sc_hd__or4_2 _21374_ (.A(_18010_),
    .B(_18011_),
    .C(_18012_),
    .D(_18013_),
    .X(_18014_));
 sky130_fd_sc_hd__or4_2 _21375_ (.A(_17976_),
    .B(_17979_),
    .C(\irq_pending[7] ),
    .D(_17973_),
    .X(_18015_));
 sky130_fd_sc_hd__or4_2 _21376_ (.A(_17994_),
    .B(\irq_pending[0] ),
    .C(_17984_),
    .D(\irq_pending[2] ),
    .X(_18016_));
 sky130_fd_sc_hd__or4_2 _21377_ (.A(_17943_),
    .B(_17946_),
    .C(\irq_pending[15] ),
    .D(_17940_),
    .X(_18017_));
 sky130_fd_sc_hd__or4_2 _21378_ (.A(_17959_),
    .B(_17962_),
    .C(\irq_pending[11] ),
    .D(_17956_),
    .X(_18018_));
 sky130_fd_sc_hd__or4_2 _21379_ (.A(_18015_),
    .B(_18016_),
    .C(_18017_),
    .D(_18018_),
    .X(_18019_));
 sky130_fd_sc_hd__nor2_2 _21380_ (.A(_18014_),
    .B(_18019_),
    .Y(_02410_));
 sky130_vsdinv _21381_ (.A(_02410_),
    .Y(_18020_));
 sky130_fd_sc_hd__and4_2 _21382_ (.A(_16902_),
    .B(_16913_),
    .C(_16918_),
    .D(_16923_),
    .X(_18021_));
 sky130_fd_sc_hd__buf_1 _21383_ (.A(_16881_),
    .X(_18022_));
 sky130_fd_sc_hd__o21a_2 _21384_ (.A1(_17255_),
    .A2(do_waitirq),
    .B1(instr_waitirq),
    .X(_18023_));
 sky130_fd_sc_hd__o2111ai_2 _21385_ (.A1(_16924_),
    .A2(_18021_),
    .B1(_16815_),
    .C1(_18022_),
    .D1(_18023_),
    .Y(_18024_));
 sky130_fd_sc_hd__nor3_2 _21386_ (.A(_00322_),
    .B(_18020_),
    .C(_18024_),
    .Y(_03830_));
 sky130_fd_sc_hd__nor3_2 _21387_ (.A(_16981_),
    .B(instr_sltu),
    .C(instr_slt),
    .Y(_18025_));
 sky130_fd_sc_hd__buf_1 _21388_ (.A(_17289_),
    .X(_18026_));
 sky130_fd_sc_hd__buf_1 _21389_ (.A(_18026_),
    .X(_18027_));
 sky130_fd_sc_hd__a211oi_2 _21390_ (.A1(_18025_),
    .A2(_17011_),
    .B1(_18001_),
    .C1(_18027_),
    .Y(_03829_));
 sky130_fd_sc_hd__buf_1 _21391_ (.A(_16823_),
    .X(_18028_));
 sky130_vsdinv _21392_ (.A(\cpu_state[5] ),
    .Y(_18029_));
 sky130_fd_sc_hd__buf_1 _21393_ (.A(_18029_),
    .X(_18030_));
 sky130_fd_sc_hd__a2111oi_2 _21394_ (.A1(_18028_),
    .A2(_18030_),
    .B1(_17211_),
    .C1(_17080_),
    .D1(_17386_),
    .Y(_03828_));
 sky130_fd_sc_hd__and3_2 _21395_ (.A(_17374_),
    .B(_17804_),
    .C(_17373_),
    .X(_03827_));
 sky130_fd_sc_hd__and2_2 _21396_ (.A(_17194_),
    .B(_02435_),
    .X(_03826_));
 sky130_fd_sc_hd__buf_1 _21397_ (.A(_17325_),
    .X(_18031_));
 sky130_fd_sc_hd__and2_2 _21398_ (.A(_18031_),
    .B(_02434_),
    .X(_03825_));
 sky130_fd_sc_hd__and2_2 _21399_ (.A(_18031_),
    .B(_02432_),
    .X(_03824_));
 sky130_fd_sc_hd__and2_2 _21400_ (.A(_18031_),
    .B(_02431_),
    .X(_03823_));
 sky130_fd_sc_hd__and2_2 _21401_ (.A(_18031_),
    .B(_02430_),
    .X(_03822_));
 sky130_fd_sc_hd__buf_1 _21402_ (.A(_17325_),
    .X(_18032_));
 sky130_fd_sc_hd__and2_2 _21403_ (.A(_18032_),
    .B(_02429_),
    .X(_03821_));
 sky130_fd_sc_hd__and2_2 _21404_ (.A(_18032_),
    .B(_02428_),
    .X(_03820_));
 sky130_fd_sc_hd__and2_2 _21405_ (.A(_18032_),
    .B(_02427_),
    .X(_03819_));
 sky130_fd_sc_hd__and2_2 _21406_ (.A(_18032_),
    .B(_02426_),
    .X(_03818_));
 sky130_fd_sc_hd__buf_1 _21407_ (.A(_17324_),
    .X(_18033_));
 sky130_fd_sc_hd__buf_1 _21408_ (.A(_18033_),
    .X(_18034_));
 sky130_fd_sc_hd__and2_2 _21409_ (.A(_18034_),
    .B(_02425_),
    .X(_03817_));
 sky130_fd_sc_hd__and2_2 _21410_ (.A(_18034_),
    .B(_02424_),
    .X(_03816_));
 sky130_fd_sc_hd__and2_2 _21411_ (.A(_18034_),
    .B(_02423_),
    .X(_03815_));
 sky130_fd_sc_hd__and2_2 _21412_ (.A(_18034_),
    .B(_02421_),
    .X(_03814_));
 sky130_fd_sc_hd__buf_1 _21413_ (.A(_18033_),
    .X(_18035_));
 sky130_fd_sc_hd__and2_2 _21414_ (.A(_18035_),
    .B(_02420_),
    .X(_03813_));
 sky130_fd_sc_hd__and2_2 _21415_ (.A(_18035_),
    .B(_02419_),
    .X(_03812_));
 sky130_fd_sc_hd__and2_2 _21416_ (.A(_18035_),
    .B(_02418_),
    .X(_03811_));
 sky130_fd_sc_hd__and2_2 _21417_ (.A(_18035_),
    .B(_02417_),
    .X(_03810_));
 sky130_fd_sc_hd__buf_1 _21418_ (.A(_18033_),
    .X(_18036_));
 sky130_fd_sc_hd__and2_2 _21419_ (.A(_18036_),
    .B(_02416_),
    .X(_03809_));
 sky130_fd_sc_hd__and2_2 _21420_ (.A(_18036_),
    .B(_02415_),
    .X(_03808_));
 sky130_fd_sc_hd__and2_2 _21421_ (.A(_18036_),
    .B(_02414_),
    .X(_03807_));
 sky130_fd_sc_hd__and2_2 _21422_ (.A(_18036_),
    .B(_02413_),
    .X(_03806_));
 sky130_fd_sc_hd__buf_1 _21423_ (.A(_18033_),
    .X(_18037_));
 sky130_fd_sc_hd__and2_2 _21424_ (.A(_18037_),
    .B(_02412_),
    .X(_03805_));
 sky130_fd_sc_hd__and2_2 _21425_ (.A(_18037_),
    .B(_02442_),
    .X(_03804_));
 sky130_fd_sc_hd__and2_2 _21426_ (.A(_18037_),
    .B(_02441_),
    .X(_03803_));
 sky130_fd_sc_hd__and2_2 _21427_ (.A(_18037_),
    .B(_02440_),
    .X(_03802_));
 sky130_fd_sc_hd__buf_1 _21428_ (.A(_17324_),
    .X(_18038_));
 sky130_fd_sc_hd__buf_1 _21429_ (.A(_18038_),
    .X(_18039_));
 sky130_fd_sc_hd__and2_2 _21430_ (.A(_18039_),
    .B(_02439_),
    .X(_03801_));
 sky130_fd_sc_hd__and2_2 _21431_ (.A(_18039_),
    .B(_02438_),
    .X(_03800_));
 sky130_fd_sc_hd__and2_2 _21432_ (.A(_18039_),
    .B(_02437_),
    .X(_03799_));
 sky130_fd_sc_hd__and2_2 _21433_ (.A(_18039_),
    .B(_02436_),
    .X(_03798_));
 sky130_fd_sc_hd__buf_1 _21434_ (.A(_18038_),
    .X(_18040_));
 sky130_fd_sc_hd__and2_2 _21435_ (.A(_18040_),
    .B(_02433_),
    .X(_03797_));
 sky130_fd_sc_hd__and2_2 _21436_ (.A(_18040_),
    .B(_02422_),
    .X(_03796_));
 sky130_fd_sc_hd__and2_2 _21437_ (.A(_18040_),
    .B(_02411_),
    .X(_03795_));
 sky130_fd_sc_hd__inv_2 _21438_ (.A(\count_cycle[18] ),
    .Y(_01938_));
 sky130_fd_sc_hd__inv_2 _21439_ (.A(\count_cycle[11] ),
    .Y(_01859_));
 sky130_fd_sc_hd__inv_2 _21440_ (.A(\count_cycle[8] ),
    .Y(_01820_));
 sky130_fd_sc_hd__inv_2 _21441_ (.A(\count_cycle[3] ),
    .Y(_01754_));
 sky130_fd_sc_hd__nand3_2 _21442_ (.A(\count_cycle[0] ),
    .B(\count_cycle[1] ),
    .C(\count_cycle[2] ),
    .Y(_18041_));
 sky130_fd_sc_hd__nor2_2 _21443_ (.A(_01754_),
    .B(_18041_),
    .Y(_18042_));
 sky130_fd_sc_hd__and3_2 _21444_ (.A(_18042_),
    .B(\count_cycle[4] ),
    .C(\count_cycle[5] ),
    .X(_18043_));
 sky130_fd_sc_hd__nand3_2 _21445_ (.A(_18043_),
    .B(\count_cycle[6] ),
    .C(\count_cycle[7] ),
    .Y(_18044_));
 sky130_fd_sc_hd__nor2_2 _21446_ (.A(_01820_),
    .B(_18044_),
    .Y(_18045_));
 sky130_fd_sc_hd__nand3_2 _21447_ (.A(_18045_),
    .B(\count_cycle[9] ),
    .C(\count_cycle[10] ),
    .Y(_18046_));
 sky130_fd_sc_hd__nor2_2 _21448_ (.A(_01859_),
    .B(_18046_),
    .Y(_18047_));
 sky130_fd_sc_hd__and2_2 _21449_ (.A(\count_cycle[14] ),
    .B(\count_cycle[15] ),
    .X(_18048_));
 sky130_fd_sc_hd__and4_2 _21450_ (.A(_18047_),
    .B(\count_cycle[12] ),
    .C(\count_cycle[13] ),
    .D(_18048_),
    .X(_18049_));
 sky130_fd_sc_hd__nand3_2 _21451_ (.A(_18049_),
    .B(\count_cycle[16] ),
    .C(\count_cycle[17] ),
    .Y(_18050_));
 sky130_fd_sc_hd__nor2_2 _21452_ (.A(_01938_),
    .B(_18050_),
    .Y(_18051_));
 sky130_fd_sc_hd__and4_2 _21453_ (.A(_18051_),
    .B(\count_cycle[19] ),
    .C(\count_cycle[20] ),
    .D(\count_cycle[21] ),
    .X(_18052_));
 sky130_fd_sc_hd__buf_1 _21454_ (.A(\count_cycle[24] ),
    .X(_18053_));
 sky130_fd_sc_hd__and2_2 _21455_ (.A(\count_cycle[22] ),
    .B(\count_cycle[23] ),
    .X(_18054_));
 sky130_fd_sc_hd__and4_2 _21456_ (.A(_18052_),
    .B(_18053_),
    .C(\count_cycle[25] ),
    .D(_18054_),
    .X(_18055_));
 sky130_fd_sc_hd__and4_2 _21457_ (.A(\count_cycle[28] ),
    .B(\count_cycle[29] ),
    .C(\count_cycle[30] ),
    .D(\count_cycle[31] ),
    .X(_18056_));
 sky130_fd_sc_hd__and4_2 _21458_ (.A(_18055_),
    .B(\count_cycle[26] ),
    .C(\count_cycle[27] ),
    .D(_18056_),
    .X(_18057_));
 sky130_fd_sc_hd__buf_1 _21459_ (.A(\count_cycle[32] ),
    .X(_18058_));
 sky130_fd_sc_hd__buf_1 _21460_ (.A(\count_cycle[33] ),
    .X(_18059_));
 sky130_fd_sc_hd__and4_2 _21461_ (.A(_18057_),
    .B(_18058_),
    .C(_18059_),
    .D(\count_cycle[34] ),
    .X(_18060_));
 sky130_fd_sc_hd__and4_2 _21462_ (.A(_18060_),
    .B(\count_cycle[35] ),
    .C(\count_cycle[36] ),
    .D(\count_cycle[37] ),
    .X(_18061_));
 sky130_fd_sc_hd__buf_1 _21463_ (.A(\count_cycle[40] ),
    .X(_18062_));
 sky130_fd_sc_hd__and2_2 _21464_ (.A(\count_cycle[38] ),
    .B(\count_cycle[39] ),
    .X(_18063_));
 sky130_fd_sc_hd__buf_1 _21465_ (.A(_18063_),
    .X(_18064_));
 sky130_fd_sc_hd__and4_2 _21466_ (.A(_18061_),
    .B(_18062_),
    .C(\count_cycle[41] ),
    .D(_18064_),
    .X(_18065_));
 sky130_fd_sc_hd__and4_2 _21467_ (.A(\count_cycle[44] ),
    .B(\count_cycle[45] ),
    .C(\count_cycle[46] ),
    .D(\count_cycle[47] ),
    .X(_18066_));
 sky130_fd_sc_hd__and4_2 _21468_ (.A(_18065_),
    .B(\count_cycle[42] ),
    .C(\count_cycle[43] ),
    .D(_18066_),
    .X(_18067_));
 sky130_fd_sc_hd__and4_2 _21469_ (.A(_18067_),
    .B(\count_cycle[48] ),
    .C(\count_cycle[49] ),
    .D(\count_cycle[50] ),
    .X(_18068_));
 sky130_fd_sc_hd__and4_2 _21470_ (.A(_18068_),
    .B(\count_cycle[51] ),
    .C(\count_cycle[52] ),
    .D(\count_cycle[53] ),
    .X(_18069_));
 sky130_fd_sc_hd__buf_1 _21471_ (.A(\count_cycle[56] ),
    .X(_18070_));
 sky130_fd_sc_hd__and2_2 _21472_ (.A(\count_cycle[54] ),
    .B(\count_cycle[55] ),
    .X(_18071_));
 sky130_fd_sc_hd__and4_2 _21473_ (.A(_18069_),
    .B(_18070_),
    .C(\count_cycle[57] ),
    .D(_18071_),
    .X(_18072_));
 sky130_fd_sc_hd__buf_1 _21474_ (.A(\count_cycle[59] ),
    .X(_18073_));
 sky130_fd_sc_hd__and4_2 _21475_ (.A(_18072_),
    .B(\count_cycle[58] ),
    .C(_18073_),
    .D(\count_cycle[60] ),
    .X(_18074_));
 sky130_fd_sc_hd__buf_1 _21476_ (.A(\count_cycle[61] ),
    .X(_18075_));
 sky130_fd_sc_hd__and4_2 _21477_ (.A(_18074_),
    .B(_18075_),
    .C(\count_cycle[62] ),
    .D(\count_cycle[63] ),
    .X(_18076_));
 sky130_vsdinv _21478_ (.A(\count_cycle[32] ),
    .Y(_18077_));
 sky130_fd_sc_hd__inv_2 _21479_ (.A(\count_cycle[19] ),
    .Y(_01947_));
 sky130_fd_sc_hd__nor3_2 _21480_ (.A(_01938_),
    .B(_01947_),
    .C(_18050_),
    .Y(_18078_));
 sky130_fd_sc_hd__and4_2 _21481_ (.A(_18078_),
    .B(\count_cycle[20] ),
    .C(\count_cycle[21] ),
    .D(_18054_),
    .X(_18079_));
 sky130_fd_sc_hd__and4_2 _21482_ (.A(_18079_),
    .B(\count_cycle[24] ),
    .C(\count_cycle[25] ),
    .D(\count_cycle[26] ),
    .X(_18080_));
 sky130_fd_sc_hd__nand3_2 _21483_ (.A(_18080_),
    .B(\count_cycle[27] ),
    .C(_18056_),
    .Y(_18081_));
 sky130_fd_sc_hd__nor3b_2 _21484_ (.A(_18077_),
    .B(_18081_),
    .C_N(\count_cycle[33] ),
    .Y(_18082_));
 sky130_fd_sc_hd__and4_2 _21485_ (.A(_18082_),
    .B(\count_cycle[34] ),
    .C(\count_cycle[35] ),
    .D(\count_cycle[36] ),
    .X(_18083_));
 sky130_fd_sc_hd__and4_2 _21486_ (.A(_18083_),
    .B(\count_cycle[37] ),
    .C(\count_cycle[40] ),
    .D(_18063_),
    .X(_18084_));
 sky130_fd_sc_hd__and4_2 _21487_ (.A(_18084_),
    .B(\count_cycle[41] ),
    .C(\count_cycle[42] ),
    .D(\count_cycle[43] ),
    .X(_18085_));
 sky130_fd_sc_hd__buf_1 _21488_ (.A(_18066_),
    .X(_18086_));
 sky130_fd_sc_hd__and4_2 _21489_ (.A(_18085_),
    .B(\count_cycle[48] ),
    .C(\count_cycle[49] ),
    .D(_18086_),
    .X(_18087_));
 sky130_fd_sc_hd__buf_1 _21490_ (.A(\count_cycle[50] ),
    .X(_18088_));
 sky130_fd_sc_hd__and4_2 _21491_ (.A(_18087_),
    .B(_18088_),
    .C(\count_cycle[51] ),
    .D(\count_cycle[52] ),
    .X(_18089_));
 sky130_fd_sc_hd__and4_2 _21492_ (.A(_18089_),
    .B(\count_cycle[53] ),
    .C(\count_cycle[56] ),
    .D(_18071_),
    .X(_18090_));
 sky130_fd_sc_hd__buf_1 _21493_ (.A(\count_cycle[57] ),
    .X(_18091_));
 sky130_fd_sc_hd__and4_2 _21494_ (.A(_18090_),
    .B(_18091_),
    .C(\count_cycle[58] ),
    .D(\count_cycle[59] ),
    .X(_18092_));
 sky130_fd_sc_hd__buf_1 _21495_ (.A(\count_cycle[60] ),
    .X(_18093_));
 sky130_fd_sc_hd__and4_2 _21496_ (.A(_18092_),
    .B(_18093_),
    .C(\count_cycle[61] ),
    .D(\count_cycle[62] ),
    .X(_18094_));
 sky130_fd_sc_hd__buf_1 _21497_ (.A(_16932_),
    .X(_18095_));
 sky130_fd_sc_hd__o21bai_2 _21498_ (.A1(\count_cycle[63] ),
    .A2(_18094_),
    .B1_N(_18095_),
    .Y(_18096_));
 sky130_fd_sc_hd__nor2_2 _21499_ (.A(_18076_),
    .B(_18096_),
    .Y(_03794_));
 sky130_fd_sc_hd__buf_1 _21500_ (.A(_18073_),
    .X(_18097_));
 sky130_fd_sc_hd__nor2_2 _21501_ (.A(_18077_),
    .B(_18081_),
    .Y(_18098_));
 sky130_fd_sc_hd__buf_1 _21502_ (.A(\count_cycle[34] ),
    .X(_18099_));
 sky130_fd_sc_hd__and4_2 _21503_ (.A(_18098_),
    .B(_18059_),
    .C(_18099_),
    .D(\count_cycle[35] ),
    .X(_18100_));
 sky130_fd_sc_hd__buf_1 _21504_ (.A(\count_cycle[36] ),
    .X(_18101_));
 sky130_fd_sc_hd__and4_2 _21505_ (.A(_18100_),
    .B(_18101_),
    .C(\count_cycle[37] ),
    .D(_18064_),
    .X(_18102_));
 sky130_fd_sc_hd__and4_2 _21506_ (.A(_18102_),
    .B(_18062_),
    .C(\count_cycle[41] ),
    .D(\count_cycle[42] ),
    .X(_18103_));
 sky130_fd_sc_hd__and4_2 _21507_ (.A(_18103_),
    .B(\count_cycle[43] ),
    .C(\count_cycle[48] ),
    .D(_18086_),
    .X(_18104_));
 sky130_fd_sc_hd__buf_1 _21508_ (.A(\count_cycle[49] ),
    .X(_18105_));
 sky130_fd_sc_hd__and4_2 _21509_ (.A(_18104_),
    .B(_18105_),
    .C(_18088_),
    .D(\count_cycle[51] ),
    .X(_18106_));
 sky130_fd_sc_hd__buf_1 _21510_ (.A(\count_cycle[52] ),
    .X(_18107_));
 sky130_fd_sc_hd__and4_2 _21511_ (.A(_18106_),
    .B(_18107_),
    .C(\count_cycle[53] ),
    .D(_18071_),
    .X(_18108_));
 sky130_fd_sc_hd__and4_2 _21512_ (.A(_18108_),
    .B(_18070_),
    .C(_18091_),
    .D(\count_cycle[58] ),
    .X(_18109_));
 sky130_fd_sc_hd__buf_1 _21513_ (.A(_18093_),
    .X(_18110_));
 sky130_fd_sc_hd__a41oi_2 _21514_ (.A1(_18097_),
    .A2(_18109_),
    .A3(_18110_),
    .A4(_18075_),
    .B1(\count_cycle[62] ),
    .Y(_18111_));
 sky130_fd_sc_hd__nor3_2 _21515_ (.A(_17857_),
    .B(_18111_),
    .C(_18094_),
    .Y(_03793_));
 sky130_fd_sc_hd__a31oi_2 _21516_ (.A1(_18109_),
    .A2(_18097_),
    .A3(_18110_),
    .B1(_18075_),
    .Y(_18112_));
 sky130_fd_sc_hd__and4_2 _21517_ (.A(_18109_),
    .B(_18073_),
    .C(_18093_),
    .D(\count_cycle[61] ),
    .X(_18113_));
 sky130_fd_sc_hd__nor3_2 _21518_ (.A(_17857_),
    .B(_18112_),
    .C(_18113_),
    .Y(_03792_));
 sky130_fd_sc_hd__a31oi_2 _21519_ (.A1(_18109_),
    .A2(_18097_),
    .A3(_18110_),
    .B1(_17808_),
    .Y(_18114_));
 sky130_fd_sc_hd__o21a_2 _21520_ (.A1(_18110_),
    .A2(_18092_),
    .B1(_18114_),
    .X(_03791_));
 sky130_fd_sc_hd__buf_1 _21521_ (.A(_18070_),
    .X(_18115_));
 sky130_fd_sc_hd__buf_1 _21522_ (.A(_18091_),
    .X(_18116_));
 sky130_fd_sc_hd__buf_1 _21523_ (.A(\count_cycle[58] ),
    .X(_18117_));
 sky130_fd_sc_hd__a41oi_2 _21524_ (.A1(_18115_),
    .A2(_18108_),
    .A3(_18116_),
    .A4(_18117_),
    .B1(_18097_),
    .Y(_18118_));
 sky130_fd_sc_hd__nor3_2 _21525_ (.A(_17857_),
    .B(_18118_),
    .C(_18092_),
    .Y(_03790_));
 sky130_fd_sc_hd__buf_1 _21526_ (.A(_17768_),
    .X(_18119_));
 sky130_fd_sc_hd__a41oi_2 _21527_ (.A1(_18115_),
    .A2(_18108_),
    .A3(_18116_),
    .A4(_18117_),
    .B1(_18119_),
    .Y(_18120_));
 sky130_fd_sc_hd__o21a_2 _21528_ (.A1(_18117_),
    .A2(_18072_),
    .B1(_18120_),
    .X(_03789_));
 sky130_fd_sc_hd__buf_1 _21529_ (.A(_17688_),
    .X(_18121_));
 sky130_fd_sc_hd__a31oi_2 _21530_ (.A1(_18108_),
    .A2(_18115_),
    .A3(_18116_),
    .B1(_18121_),
    .Y(_18122_));
 sky130_fd_sc_hd__o21a_2 _21531_ (.A1(_18116_),
    .A2(_18090_),
    .B1(_18122_),
    .X(_03788_));
 sky130_fd_sc_hd__buf_1 _21532_ (.A(_17856_),
    .X(_18123_));
 sky130_fd_sc_hd__buf_1 _21533_ (.A(_18107_),
    .X(_18124_));
 sky130_fd_sc_hd__buf_1 _21534_ (.A(_18106_),
    .X(_18125_));
 sky130_fd_sc_hd__buf_1 _21535_ (.A(\count_cycle[53] ),
    .X(_18126_));
 sky130_fd_sc_hd__buf_1 _21536_ (.A(_18126_),
    .X(_18127_));
 sky130_fd_sc_hd__a41oi_2 _21537_ (.A1(_18124_),
    .A2(_18125_),
    .A3(_18127_),
    .A4(_18071_),
    .B1(_18115_),
    .Y(_18128_));
 sky130_fd_sc_hd__nor3_2 _21538_ (.A(_18123_),
    .B(_18128_),
    .C(_18090_),
    .Y(_03787_));
 sky130_fd_sc_hd__buf_1 _21539_ (.A(\count_cycle[54] ),
    .X(_18129_));
 sky130_fd_sc_hd__and4_2 _21540_ (.A(_18089_),
    .B(_18126_),
    .C(_18129_),
    .D(\count_cycle[55] ),
    .X(_18130_));
 sky130_fd_sc_hd__and4_2 _21541_ (.A(_18125_),
    .B(_18107_),
    .C(_18126_),
    .D(_18129_),
    .X(_18131_));
 sky130_fd_sc_hd__o21bai_2 _21542_ (.A1(\count_cycle[55] ),
    .A2(_18131_),
    .B1_N(_18095_),
    .Y(_18132_));
 sky130_fd_sc_hd__nor2_2 _21543_ (.A(_18130_),
    .B(_18132_),
    .Y(_03786_));
 sky130_fd_sc_hd__a31oi_2 _21544_ (.A1(_18125_),
    .A2(_18107_),
    .A3(_18127_),
    .B1(_18129_),
    .Y(_18133_));
 sky130_fd_sc_hd__nor3_2 _21545_ (.A(_18123_),
    .B(_18133_),
    .C(_18131_),
    .Y(_03785_));
 sky130_fd_sc_hd__a31oi_2 _21546_ (.A1(_18125_),
    .A2(_18124_),
    .A3(_18127_),
    .B1(_18121_),
    .Y(_18134_));
 sky130_fd_sc_hd__o21a_2 _21547_ (.A1(_18127_),
    .A2(_18089_),
    .B1(_18134_),
    .X(_03784_));
 sky130_fd_sc_hd__buf_1 _21548_ (.A(_18104_),
    .X(_18135_));
 sky130_fd_sc_hd__buf_1 _21549_ (.A(\count_cycle[51] ),
    .X(_18136_));
 sky130_fd_sc_hd__a41oi_2 _21550_ (.A1(_18105_),
    .A2(_18135_),
    .A3(_18088_),
    .A4(_18136_),
    .B1(_18124_),
    .Y(_18137_));
 sky130_fd_sc_hd__nor3_2 _21551_ (.A(_18123_),
    .B(_18137_),
    .C(_18089_),
    .Y(_03783_));
 sky130_fd_sc_hd__buf_1 _21552_ (.A(_18105_),
    .X(_18138_));
 sky130_fd_sc_hd__buf_1 _21553_ (.A(_18088_),
    .X(_18139_));
 sky130_fd_sc_hd__a41oi_2 _21554_ (.A1(_18138_),
    .A2(_18135_),
    .A3(_18139_),
    .A4(_18136_),
    .B1(_18119_),
    .Y(_18140_));
 sky130_fd_sc_hd__o21a_2 _21555_ (.A1(_18136_),
    .A2(_18068_),
    .B1(_18140_),
    .X(_03782_));
 sky130_fd_sc_hd__a31oi_2 _21556_ (.A1(_18135_),
    .A2(_18138_),
    .A3(_18139_),
    .B1(_18121_),
    .Y(_18141_));
 sky130_fd_sc_hd__o21a_2 _21557_ (.A1(_18139_),
    .A2(_18087_),
    .B1(_18141_),
    .X(_03781_));
 sky130_fd_sc_hd__buf_1 _21558_ (.A(\count_cycle[48] ),
    .X(_18142_));
 sky130_fd_sc_hd__buf_1 _21559_ (.A(_18085_),
    .X(_18143_));
 sky130_fd_sc_hd__a41oi_2 _21560_ (.A1(_18142_),
    .A2(_18143_),
    .A3(_18105_),
    .A4(_18086_),
    .B1(_18119_),
    .Y(_18144_));
 sky130_fd_sc_hd__o21a_2 _21561_ (.A1(_18138_),
    .A2(_18135_),
    .B1(_18144_),
    .X(_03780_));
 sky130_fd_sc_hd__buf_1 _21562_ (.A(\count_cycle[43] ),
    .X(_18145_));
 sky130_fd_sc_hd__buf_1 _21563_ (.A(_18145_),
    .X(_18146_));
 sky130_fd_sc_hd__buf_1 _21564_ (.A(_18103_),
    .X(_18147_));
 sky130_fd_sc_hd__a41oi_2 _21565_ (.A1(_18146_),
    .A2(_18147_),
    .A3(_18142_),
    .A4(_18086_),
    .B1(_18119_),
    .Y(_18148_));
 sky130_fd_sc_hd__o21a_2 _21566_ (.A1(_18142_),
    .A2(_18067_),
    .B1(_18148_),
    .X(_03779_));
 sky130_fd_sc_hd__buf_1 _21567_ (.A(\count_cycle[42] ),
    .X(_18149_));
 sky130_fd_sc_hd__buf_1 _21568_ (.A(\count_cycle[44] ),
    .X(_18150_));
 sky130_fd_sc_hd__and4_2 _21569_ (.A(_18065_),
    .B(_18149_),
    .C(_18145_),
    .D(_18150_),
    .X(_18151_));
 sky130_fd_sc_hd__buf_1 _21570_ (.A(\count_cycle[46] ),
    .X(_18152_));
 sky130_fd_sc_hd__and4_2 _21571_ (.A(_18151_),
    .B(\count_cycle[45] ),
    .C(_18152_),
    .D(\count_cycle[47] ),
    .X(_18153_));
 sky130_fd_sc_hd__and4_2 _21572_ (.A(_18143_),
    .B(_18150_),
    .C(\count_cycle[45] ),
    .D(_18152_),
    .X(_18154_));
 sky130_fd_sc_hd__o21bai_2 _21573_ (.A1(\count_cycle[47] ),
    .A2(_18154_),
    .B1_N(_18095_),
    .Y(_18155_));
 sky130_fd_sc_hd__nor2_2 _21574_ (.A(_18153_),
    .B(_18155_),
    .Y(_03778_));
 sky130_fd_sc_hd__buf_1 _21575_ (.A(_18150_),
    .X(_18156_));
 sky130_fd_sc_hd__buf_1 _21576_ (.A(\count_cycle[45] ),
    .X(_18157_));
 sky130_fd_sc_hd__a41oi_2 _21577_ (.A1(_18145_),
    .A2(_18103_),
    .A3(_18156_),
    .A4(_18157_),
    .B1(_18152_),
    .Y(_18158_));
 sky130_fd_sc_hd__nor3_2 _21578_ (.A(_18123_),
    .B(_18158_),
    .C(_18154_),
    .Y(_03777_));
 sky130_fd_sc_hd__buf_1 _21579_ (.A(_17768_),
    .X(_18159_));
 sky130_fd_sc_hd__a41oi_2 _21580_ (.A1(_18146_),
    .A2(_18147_),
    .A3(_18156_),
    .A4(_18157_),
    .B1(_18159_),
    .Y(_18160_));
 sky130_fd_sc_hd__o21a_2 _21581_ (.A1(_18157_),
    .A2(_18151_),
    .B1(_18160_),
    .X(_03776_));
 sky130_fd_sc_hd__a31oi_2 _21582_ (.A1(_18147_),
    .A2(_18145_),
    .A3(_18156_),
    .B1(_18121_),
    .Y(_18161_));
 sky130_fd_sc_hd__o21a_2 _21583_ (.A1(_18156_),
    .A2(_18143_),
    .B1(_18161_),
    .X(_03775_));
 sky130_fd_sc_hd__buf_1 _21584_ (.A(_17856_),
    .X(_18162_));
 sky130_fd_sc_hd__buf_1 _21585_ (.A(_18062_),
    .X(_18163_));
 sky130_fd_sc_hd__buf_1 _21586_ (.A(\count_cycle[41] ),
    .X(_18164_));
 sky130_fd_sc_hd__a41oi_2 _21587_ (.A1(_18163_),
    .A2(_18102_),
    .A3(_18164_),
    .A4(_18149_),
    .B1(_18146_),
    .Y(_18165_));
 sky130_fd_sc_hd__nor3_2 _21588_ (.A(_18162_),
    .B(_18165_),
    .C(_18143_),
    .Y(_03774_));
 sky130_fd_sc_hd__a31oi_2 _21589_ (.A1(_18102_),
    .A2(_18163_),
    .A3(_18164_),
    .B1(_18149_),
    .Y(_18166_));
 sky130_fd_sc_hd__nor3_2 _21590_ (.A(_18162_),
    .B(_18166_),
    .C(_18147_),
    .Y(_03773_));
 sky130_fd_sc_hd__buf_1 _21591_ (.A(\count_cycle[37] ),
    .X(_18167_));
 sky130_fd_sc_hd__buf_1 _21592_ (.A(_18167_),
    .X(_18168_));
 sky130_fd_sc_hd__a41oi_2 _21593_ (.A1(_18168_),
    .A2(_18083_),
    .A3(_18062_),
    .A4(_18064_),
    .B1(_18164_),
    .Y(_18169_));
 sky130_fd_sc_hd__nor3_2 _21594_ (.A(_18162_),
    .B(_18169_),
    .C(_18065_),
    .Y(_03772_));
 sky130_fd_sc_hd__buf_1 _21595_ (.A(_18101_),
    .X(_18170_));
 sky130_fd_sc_hd__buf_1 _21596_ (.A(_18100_),
    .X(_18171_));
 sky130_fd_sc_hd__a41oi_2 _21597_ (.A1(_18170_),
    .A2(_18171_),
    .A3(_18168_),
    .A4(_18064_),
    .B1(_18163_),
    .Y(_18172_));
 sky130_fd_sc_hd__nor3_2 _21598_ (.A(_18162_),
    .B(_18172_),
    .C(_18084_),
    .Y(_03771_));
 sky130_fd_sc_hd__buf_1 _21599_ (.A(\count_cycle[38] ),
    .X(_18173_));
 sky130_fd_sc_hd__and4_2 _21600_ (.A(_18083_),
    .B(_18167_),
    .C(_18173_),
    .D(\count_cycle[39] ),
    .X(_18174_));
 sky130_fd_sc_hd__and4_2 _21601_ (.A(_18171_),
    .B(_18101_),
    .C(_18167_),
    .D(_18173_),
    .X(_18175_));
 sky130_fd_sc_hd__o21bai_2 _21602_ (.A1(\count_cycle[39] ),
    .A2(_18175_),
    .B1_N(_18095_),
    .Y(_18176_));
 sky130_fd_sc_hd__nor2_2 _21603_ (.A(_18174_),
    .B(_18176_),
    .Y(_03770_));
 sky130_fd_sc_hd__buf_1 _21604_ (.A(_17856_),
    .X(_18177_));
 sky130_fd_sc_hd__a31oi_2 _21605_ (.A1(_18171_),
    .A2(_18170_),
    .A3(_18168_),
    .B1(_18173_),
    .Y(_18178_));
 sky130_fd_sc_hd__nor3_2 _21606_ (.A(_18177_),
    .B(_18178_),
    .C(_18175_),
    .Y(_03769_));
 sky130_fd_sc_hd__buf_1 _21607_ (.A(_18099_),
    .X(_18179_));
 sky130_fd_sc_hd__buf_1 _21608_ (.A(\count_cycle[35] ),
    .X(_18180_));
 sky130_fd_sc_hd__a41oi_2 _21609_ (.A1(_18179_),
    .A2(_18082_),
    .A3(_18180_),
    .A4(_18101_),
    .B1(_18168_),
    .Y(_18181_));
 sky130_fd_sc_hd__nor3_2 _21610_ (.A(_18177_),
    .B(_18181_),
    .C(_18061_),
    .Y(_03768_));
 sky130_fd_sc_hd__buf_1 _21611_ (.A(_18059_),
    .X(_18182_));
 sky130_fd_sc_hd__buf_1 _21612_ (.A(_18098_),
    .X(_18183_));
 sky130_fd_sc_hd__a41oi_2 _21613_ (.A1(_18182_),
    .A2(_18183_),
    .A3(_18099_),
    .A4(_18180_),
    .B1(_18170_),
    .Y(_18184_));
 sky130_fd_sc_hd__nor3_2 _21614_ (.A(_18177_),
    .B(_18184_),
    .C(_18083_),
    .Y(_03767_));
 sky130_fd_sc_hd__a31oi_2 _21615_ (.A1(_18183_),
    .A2(_18059_),
    .A3(_18179_),
    .B1(_18180_),
    .Y(_18185_));
 sky130_fd_sc_hd__nor3_2 _21616_ (.A(_18177_),
    .B(_18185_),
    .C(_18171_),
    .Y(_03766_));
 sky130_fd_sc_hd__buf_1 _21617_ (.A(_17768_),
    .X(_18186_));
 sky130_fd_sc_hd__a31oi_2 _21618_ (.A1(_18183_),
    .A2(_18182_),
    .A3(_18179_),
    .B1(_18186_),
    .Y(_18187_));
 sky130_fd_sc_hd__o21a_2 _21619_ (.A1(_18179_),
    .A2(_18082_),
    .B1(_18187_),
    .X(_03765_));
 sky130_fd_sc_hd__buf_1 _21620_ (.A(_17748_),
    .X(_18188_));
 sky130_fd_sc_hd__buf_1 _21621_ (.A(_18080_),
    .X(_18189_));
 sky130_fd_sc_hd__buf_1 _21622_ (.A(\count_cycle[27] ),
    .X(_18190_));
 sky130_fd_sc_hd__buf_1 _21623_ (.A(_18190_),
    .X(_18191_));
 sky130_fd_sc_hd__a41oi_2 _21624_ (.A1(_18058_),
    .A2(_18189_),
    .A3(_18191_),
    .A4(_18056_),
    .B1(_18182_),
    .Y(_18192_));
 sky130_fd_sc_hd__nor3_2 _21625_ (.A(_18188_),
    .B(_18192_),
    .C(_18082_),
    .Y(_03764_));
 sky130_fd_sc_hd__a31oi_2 _21626_ (.A1(_18189_),
    .A2(_18191_),
    .A3(_18056_),
    .B1(_18058_),
    .Y(_18193_));
 sky130_fd_sc_hd__nor3_2 _21627_ (.A(_18188_),
    .B(_18193_),
    .C(_18183_),
    .Y(_03763_));
 sky130_fd_sc_hd__buf_1 _21628_ (.A(_18055_),
    .X(_18194_));
 sky130_fd_sc_hd__buf_1 _21629_ (.A(\count_cycle[26] ),
    .X(_18195_));
 sky130_fd_sc_hd__and4_2 _21630_ (.A(_18194_),
    .B(_18195_),
    .C(_18190_),
    .D(\count_cycle[28] ),
    .X(_18196_));
 sky130_fd_sc_hd__and4_2 _21631_ (.A(_18196_),
    .B(\count_cycle[29] ),
    .C(\count_cycle[30] ),
    .D(\count_cycle[31] ),
    .X(_18197_));
 sky130_fd_sc_hd__inv_2 _21632_ (.A(\count_cycle[30] ),
    .Y(_02046_));
 sky130_fd_sc_hd__and3_2 _21633_ (.A(_18055_),
    .B(_18195_),
    .C(_18190_),
    .X(_18198_));
 sky130_fd_sc_hd__nand3_2 _21634_ (.A(_18198_),
    .B(\count_cycle[28] ),
    .C(\count_cycle[29] ),
    .Y(_18199_));
 sky130_fd_sc_hd__nor2_2 _21635_ (.A(_02046_),
    .B(_18199_),
    .Y(_18200_));
 sky130_fd_sc_hd__o21bai_2 _21636_ (.A1(\count_cycle[31] ),
    .A2(_18200_),
    .B1_N(_17657_),
    .Y(_18201_));
 sky130_fd_sc_hd__nor2_2 _21637_ (.A(_18197_),
    .B(_18201_),
    .Y(_03762_));
 sky130_fd_sc_hd__buf_1 _21638_ (.A(\count_cycle[28] ),
    .X(_18202_));
 sky130_fd_sc_hd__buf_1 _21639_ (.A(\count_cycle[29] ),
    .X(_18203_));
 sky130_fd_sc_hd__a41oi_2 _21640_ (.A1(_18191_),
    .A2(_18080_),
    .A3(_18202_),
    .A4(_18203_),
    .B1(\count_cycle[30] ),
    .Y(_18204_));
 sky130_fd_sc_hd__nor3_2 _21641_ (.A(_18188_),
    .B(_18204_),
    .C(_18200_),
    .Y(_03761_));
 sky130_fd_sc_hd__buf_1 _21642_ (.A(_18190_),
    .X(_18205_));
 sky130_fd_sc_hd__a41oi_2 _21643_ (.A1(_18205_),
    .A2(_18189_),
    .A3(_18202_),
    .A4(_18203_),
    .B1(_18159_),
    .Y(_18206_));
 sky130_fd_sc_hd__o21a_2 _21644_ (.A1(_18203_),
    .A2(_18196_),
    .B1(_18206_),
    .X(_03760_));
 sky130_fd_sc_hd__a31oi_2 _21645_ (.A1(_18194_),
    .A2(_18195_),
    .A3(_18191_),
    .B1(_18202_),
    .Y(_18207_));
 sky130_fd_sc_hd__nor3_2 _21646_ (.A(_18188_),
    .B(_18207_),
    .C(_18196_),
    .Y(_03759_));
 sky130_fd_sc_hd__buf_1 _21647_ (.A(_18195_),
    .X(_18208_));
 sky130_fd_sc_hd__a31oi_2 _21648_ (.A1(_18194_),
    .A2(_18208_),
    .A3(_18205_),
    .B1(_18186_),
    .Y(_18209_));
 sky130_fd_sc_hd__o21a_2 _21649_ (.A1(_18205_),
    .A2(_18189_),
    .B1(_18209_),
    .X(_03758_));
 sky130_fd_sc_hd__buf_1 _21650_ (.A(_18053_),
    .X(_18210_));
 sky130_fd_sc_hd__buf_1 _21651_ (.A(\count_cycle[25] ),
    .X(_18211_));
 sky130_fd_sc_hd__a41oi_2 _21652_ (.A1(_18210_),
    .A2(_18079_),
    .A3(_18211_),
    .A4(_18208_),
    .B1(_18159_),
    .Y(_18212_));
 sky130_fd_sc_hd__o21a_2 _21653_ (.A1(_18208_),
    .A2(_18194_),
    .B1(_18212_),
    .X(_03757_));
 sky130_fd_sc_hd__and3_2 _21654_ (.A(_18052_),
    .B(_18053_),
    .C(_18054_),
    .X(_18213_));
 sky130_fd_sc_hd__a31oi_2 _21655_ (.A1(_18079_),
    .A2(_18210_),
    .A3(_18211_),
    .B1(_18186_),
    .Y(_18214_));
 sky130_fd_sc_hd__o21a_2 _21656_ (.A1(_18211_),
    .A2(_18213_),
    .B1(_18214_),
    .X(_03756_));
 sky130_fd_sc_hd__buf_1 _21657_ (.A(_18052_),
    .X(_18215_));
 sky130_fd_sc_hd__a31oi_2 _21658_ (.A1(_18215_),
    .A2(_18053_),
    .A3(_18054_),
    .B1(_18186_),
    .Y(_18216_));
 sky130_fd_sc_hd__o21a_2 _21659_ (.A1(_18210_),
    .A2(_18079_),
    .B1(_18216_),
    .X(_03755_));
 sky130_fd_sc_hd__buf_1 _21660_ (.A(\count_cycle[22] ),
    .X(_18217_));
 sky130_fd_sc_hd__and3_2 _21661_ (.A(_18215_),
    .B(_18217_),
    .C(\count_cycle[23] ),
    .X(_18218_));
 sky130_fd_sc_hd__buf_1 _21662_ (.A(_18078_),
    .X(_18219_));
 sky130_fd_sc_hd__buf_1 _21663_ (.A(\count_cycle[20] ),
    .X(_18220_));
 sky130_fd_sc_hd__buf_1 _21664_ (.A(\count_cycle[21] ),
    .X(_18221_));
 sky130_fd_sc_hd__and4_2 _21665_ (.A(_18219_),
    .B(_18220_),
    .C(_18221_),
    .D(\count_cycle[22] ),
    .X(_18222_));
 sky130_fd_sc_hd__o21bai_2 _21666_ (.A1(\count_cycle[23] ),
    .A2(_18222_),
    .B1_N(_17657_),
    .Y(_18223_));
 sky130_fd_sc_hd__nor2_2 _21667_ (.A(_18218_),
    .B(_18223_),
    .Y(_03754_));
 sky130_fd_sc_hd__a41oi_2 _21668_ (.A1(_18220_),
    .A2(_18219_),
    .A3(_18221_),
    .A4(_18217_),
    .B1(_18159_),
    .Y(_18224_));
 sky130_fd_sc_hd__o21a_2 _21669_ (.A1(_18217_),
    .A2(_18215_),
    .B1(_18224_),
    .X(_03753_));
 sky130_fd_sc_hd__buf_1 _21670_ (.A(_17748_),
    .X(_18225_));
 sky130_fd_sc_hd__a31oi_2 _21671_ (.A1(_18051_),
    .A2(\count_cycle[19] ),
    .A3(_18220_),
    .B1(_18221_),
    .Y(_18226_));
 sky130_fd_sc_hd__nor3_2 _21672_ (.A(_18225_),
    .B(_18226_),
    .C(_18215_),
    .Y(_03752_));
 sky130_fd_sc_hd__inv_2 _21673_ (.A(_18220_),
    .Y(_01956_));
 sky130_vsdinv _21674_ (.A(_18219_),
    .Y(_18227_));
 sky130_fd_sc_hd__o41ai_2 _21675_ (.A1(_01938_),
    .A2(_01947_),
    .A3(_01956_),
    .A4(_18050_),
    .B1(_17718_),
    .Y(_18228_));
 sky130_fd_sc_hd__a21oi_2 _21676_ (.A1(_01956_),
    .A2(_18227_),
    .B1(_18228_),
    .Y(_03751_));
 sky130_fd_sc_hd__inv_2 _21677_ (.A(\count_cycle[12] ),
    .Y(_01872_));
 sky130_fd_sc_hd__nor3_2 _21678_ (.A(_01859_),
    .B(_01872_),
    .C(_18046_),
    .Y(_18229_));
 sky130_fd_sc_hd__buf_1 _21679_ (.A(\count_cycle[13] ),
    .X(_18230_));
 sky130_fd_sc_hd__and4_2 _21680_ (.A(_18229_),
    .B(_18230_),
    .C(\count_cycle[16] ),
    .D(_18048_),
    .X(_18231_));
 sky130_fd_sc_hd__buf_1 _21681_ (.A(\count_cycle[17] ),
    .X(_18232_));
 sky130_fd_sc_hd__a31oi_2 _21682_ (.A1(_18231_),
    .A2(_18232_),
    .A3(\count_cycle[18] ),
    .B1(\count_cycle[19] ),
    .Y(_18233_));
 sky130_fd_sc_hd__nor3_2 _21683_ (.A(_18225_),
    .B(_18233_),
    .C(_18219_),
    .Y(_03750_));
 sky130_fd_sc_hd__buf_1 _21684_ (.A(\count_cycle[16] ),
    .X(_18234_));
 sky130_fd_sc_hd__a31oi_2 _21685_ (.A1(_18049_),
    .A2(_18234_),
    .A3(_18232_),
    .B1(\count_cycle[18] ),
    .Y(_18235_));
 sky130_fd_sc_hd__nor3_2 _21686_ (.A(_18225_),
    .B(_18235_),
    .C(_18051_),
    .Y(_03749_));
 sky130_fd_sc_hd__a41o_2 _21687_ (.A1(_18229_),
    .A2(_18230_),
    .A3(_18234_),
    .A4(_18048_),
    .B1(_18232_),
    .X(_18236_));
 sky130_fd_sc_hd__and3_2 _21688_ (.A(_18050_),
    .B(_18236_),
    .C(_17998_),
    .X(_03748_));
 sky130_fd_sc_hd__buf_1 _21689_ (.A(_18230_),
    .X(_18237_));
 sky130_fd_sc_hd__a31oi_2 _21690_ (.A1(_18229_),
    .A2(_18237_),
    .A3(_18048_),
    .B1(_18234_),
    .Y(_18238_));
 sky130_fd_sc_hd__nor3_2 _21691_ (.A(_18225_),
    .B(_18238_),
    .C(_18231_),
    .Y(_03747_));
 sky130_fd_sc_hd__inv_2 _21692_ (.A(\count_cycle[14] ),
    .Y(_01898_));
 sky130_fd_sc_hd__buf_1 _21693_ (.A(\count_cycle[12] ),
    .X(_18239_));
 sky130_fd_sc_hd__nand3_2 _21694_ (.A(_18047_),
    .B(_18239_),
    .C(_18230_),
    .Y(_18240_));
 sky130_fd_sc_hd__nor2_2 _21695_ (.A(_01898_),
    .B(_18240_),
    .Y(_18241_));
 sky130_fd_sc_hd__o21a_2 _21696_ (.A1(\count_cycle[15] ),
    .A2(_18241_),
    .B1(_16838_),
    .X(_18242_));
 sky130_fd_sc_hd__nand3b_2 _21697_ (.A_N(_18240_),
    .B(\count_cycle[14] ),
    .C(\count_cycle[15] ),
    .Y(_18243_));
 sky130_fd_sc_hd__nand2_2 _21698_ (.A(_18242_),
    .B(_18243_),
    .Y(_18244_));
 sky130_vsdinv _21699_ (.A(_18244_),
    .Y(_03746_));
 sky130_fd_sc_hd__buf_1 _21700_ (.A(_17748_),
    .X(_18245_));
 sky130_fd_sc_hd__a31oi_2 _21701_ (.A1(_18047_),
    .A2(_18239_),
    .A3(_18237_),
    .B1(\count_cycle[14] ),
    .Y(_18246_));
 sky130_fd_sc_hd__nor3_2 _21702_ (.A(_18245_),
    .B(_18246_),
    .C(_18241_),
    .Y(_03745_));
 sky130_fd_sc_hd__inv_2 _21703_ (.A(\count_cycle[9] ),
    .Y(_01833_));
 sky130_fd_sc_hd__nor3_2 _21704_ (.A(_01820_),
    .B(_01833_),
    .C(_18044_),
    .Y(_18247_));
 sky130_fd_sc_hd__buf_1 _21705_ (.A(\count_cycle[10] ),
    .X(_18248_));
 sky130_fd_sc_hd__a41o_2 _21706_ (.A1(_18247_),
    .A2(_18248_),
    .A3(\count_cycle[11] ),
    .A4(_18239_),
    .B1(_18237_),
    .X(_18249_));
 sky130_fd_sc_hd__and3_2 _21707_ (.A(_18240_),
    .B(_18249_),
    .C(_17998_),
    .X(_03744_));
 sky130_fd_sc_hd__a31oi_2 _21708_ (.A1(_18247_),
    .A2(_18248_),
    .A3(\count_cycle[11] ),
    .B1(_18239_),
    .Y(_18250_));
 sky130_fd_sc_hd__nor3_2 _21709_ (.A(_18245_),
    .B(_18250_),
    .C(_18229_),
    .Y(_03743_));
 sky130_fd_sc_hd__a31oi_2 _21710_ (.A1(_18045_),
    .A2(\count_cycle[9] ),
    .A3(_18248_),
    .B1(\count_cycle[11] ),
    .Y(_18251_));
 sky130_fd_sc_hd__nor3_2 _21711_ (.A(_18245_),
    .B(_18251_),
    .C(_18047_),
    .Y(_03742_));
 sky130_fd_sc_hd__inv_2 _21712_ (.A(_18248_),
    .Y(_01846_));
 sky130_fd_sc_hd__o31ai_2 _21713_ (.A1(_01820_),
    .A2(_01833_),
    .A3(_18044_),
    .B1(_01846_),
    .Y(_18252_));
 sky130_fd_sc_hd__and3_2 _21714_ (.A(_18252_),
    .B(_18046_),
    .C(_17804_),
    .X(_03741_));
 sky130_fd_sc_hd__buf_1 _21715_ (.A(\count_cycle[6] ),
    .X(_18253_));
 sky130_fd_sc_hd__buf_1 _21716_ (.A(\count_cycle[7] ),
    .X(_18254_));
 sky130_fd_sc_hd__a41oi_2 _21717_ (.A1(_18253_),
    .A2(_18043_),
    .A3(_18254_),
    .A4(\count_cycle[8] ),
    .B1(\count_cycle[9] ),
    .Y(_18255_));
 sky130_fd_sc_hd__nor3_2 _21718_ (.A(_18245_),
    .B(_18255_),
    .C(_18247_),
    .Y(_03740_));
 sky130_fd_sc_hd__a31oi_2 _21719_ (.A1(_18043_),
    .A2(\count_cycle[6] ),
    .A3(_18254_),
    .B1(\count_cycle[8] ),
    .Y(_18256_));
 sky130_fd_sc_hd__nor3_2 _21720_ (.A(_17749_),
    .B(_18256_),
    .C(_18045_),
    .Y(_03739_));
 sky130_fd_sc_hd__buf_1 _21721_ (.A(\count_cycle[4] ),
    .X(_18257_));
 sky130_fd_sc_hd__a41o_2 _21722_ (.A1(_18042_),
    .A2(_18257_),
    .A3(\count_cycle[5] ),
    .A4(\count_cycle[6] ),
    .B1(_18254_),
    .X(_18258_));
 sky130_fd_sc_hd__and3_2 _21723_ (.A(_18044_),
    .B(_17804_),
    .C(_18258_),
    .X(_03738_));
 sky130_fd_sc_hd__buf_1 _21724_ (.A(\count_cycle[5] ),
    .X(_18259_));
 sky130_fd_sc_hd__a41oi_2 _21725_ (.A1(_18257_),
    .A2(_18042_),
    .A3(_18259_),
    .A4(_18253_),
    .B1(_17049_),
    .Y(_18260_));
 sky130_fd_sc_hd__o21a_2 _21726_ (.A1(_18253_),
    .A2(_18043_),
    .B1(_18260_),
    .X(_03737_));
 sky130_fd_sc_hd__inv_2 _21727_ (.A(_18257_),
    .Y(_01767_));
 sky130_fd_sc_hd__nor3_2 _21728_ (.A(_01754_),
    .B(_01767_),
    .C(_18041_),
    .Y(_18261_));
 sky130_fd_sc_hd__o21bai_2 _21729_ (.A1(_18259_),
    .A2(_18261_),
    .B1_N(_17683_),
    .Y(_18262_));
 sky130_fd_sc_hd__a21oi_2 _21730_ (.A1(_18259_),
    .A2(_18261_),
    .B1(_18262_),
    .Y(_03736_));
 sky130_fd_sc_hd__buf_1 _21731_ (.A(\count_cycle[0] ),
    .X(_18263_));
 sky130_fd_sc_hd__buf_1 _21732_ (.A(\count_cycle[2] ),
    .X(_18264_));
 sky130_fd_sc_hd__a41oi_2 _21733_ (.A1(_18263_),
    .A2(\count_cycle[1] ),
    .A3(_18264_),
    .A4(\count_cycle[3] ),
    .B1(_18257_),
    .Y(_18265_));
 sky130_fd_sc_hd__nor3_2 _21734_ (.A(_17749_),
    .B(_18261_),
    .C(_18265_),
    .Y(_03735_));
 sky130_fd_sc_hd__a31oi_2 _21735_ (.A1(_18263_),
    .A2(\count_cycle[1] ),
    .A3(_18264_),
    .B1(\count_cycle[3] ),
    .Y(_18266_));
 sky130_fd_sc_hd__nor3_2 _21736_ (.A(_17749_),
    .B(_18042_),
    .C(_18266_),
    .Y(_03734_));
 sky130_fd_sc_hd__buf_1 _21737_ (.A(\count_cycle[1] ),
    .X(_18267_));
 sky130_fd_sc_hd__a21oi_2 _21738_ (.A1(_18263_),
    .A2(_18267_),
    .B1(_18264_),
    .Y(_18268_));
 sky130_fd_sc_hd__nor3b_2 _21739_ (.A(_17782_),
    .B(_18268_),
    .C_N(_18041_),
    .Y(_03733_));
 sky130_fd_sc_hd__buf_1 _21740_ (.A(_18263_),
    .X(_18269_));
 sky130_fd_sc_hd__a21boi_2 _21741_ (.A1(_18269_),
    .A2(_18267_),
    .B1_N(_17325_),
    .Y(_18270_));
 sky130_fd_sc_hd__o21a_2 _21742_ (.A1(_18269_),
    .A2(_18267_),
    .B1(_18270_),
    .X(_03732_));
 sky130_vsdinv _21743_ (.A(_18269_),
    .Y(_02559_));
 sky130_fd_sc_hd__nor2b_2 _21744_ (.A(_18269_),
    .B_N(_16832_),
    .Y(_03731_));
 sky130_fd_sc_hd__and2_2 _21745_ (.A(_18040_),
    .B(\cpu_state[0] ),
    .X(_03730_));
 sky130_fd_sc_hd__buf_1 _21746_ (.A(_18038_),
    .X(_18271_));
 sky130_fd_sc_hd__and2_2 _21747_ (.A(_18271_),
    .B(\pcpi_mul.active[0] ),
    .X(_03729_));
 sky130_fd_sc_hd__buf_1 _21748_ (.A(\cpuregs_wrdata[31] ),
    .X(_18272_));
 sky130_fd_sc_hd__buf_1 _21749_ (.A(_18272_),
    .X(_18273_));
 sky130_fd_sc_hd__or2_2 _21750_ (.A(\latched_rd[0] ),
    .B(\latched_rd[1] ),
    .X(_18274_));
 sky130_fd_sc_hd__buf_1 _21751_ (.A(_18274_),
    .X(_18275_));
 sky130_fd_sc_hd__buf_1 _21752_ (.A(_18275_),
    .X(_18276_));
 sky130_vsdinv _21753_ (.A(\latched_rd[2] ),
    .Y(_18277_));
 sky130_vsdinv _21754_ (.A(\latched_rd[3] ),
    .Y(_18278_));
 sky130_fd_sc_hd__nand3b_2 _21755_ (.A_N(\latched_rd[4] ),
    .B(_18277_),
    .C(_18278_),
    .Y(_18279_));
 sky130_fd_sc_hd__buf_1 _21756_ (.A(_18279_),
    .X(_18280_));
 sky130_fd_sc_hd__buf_1 _21757_ (.A(_18280_),
    .X(_18281_));
 sky130_fd_sc_hd__buf_1 _21758_ (.A(_18281_),
    .X(_18282_));
 sky130_fd_sc_hd__buf_1 _21759_ (.A(\latched_rd[0] ),
    .X(_18283_));
 sky130_fd_sc_hd__buf_1 _21760_ (.A(\latched_rd[1] ),
    .X(_18284_));
 sky130_fd_sc_hd__and2b_2 _21761_ (.A_N(_18283_),
    .B(_18284_),
    .X(_18285_));
 sky130_fd_sc_hd__buf_1 _21762_ (.A(_18285_),
    .X(_18286_));
 sky130_fd_sc_hd__buf_1 _21763_ (.A(\latched_rd[4] ),
    .X(_18287_));
 sky130_fd_sc_hd__buf_1 _21764_ (.A(\latched_rd[3] ),
    .X(_18288_));
 sky130_fd_sc_hd__buf_1 _21765_ (.A(\latched_rd[2] ),
    .X(_18289_));
 sky130_fd_sc_hd__nor3b_2 _21766_ (.A(_18287_),
    .B(_18288_),
    .C_N(_18289_),
    .Y(_18290_));
 sky130_fd_sc_hd__and2_2 _21767_ (.A(resetn),
    .B(\cpu_state[1] ),
    .X(_18291_));
 sky130_fd_sc_hd__o41a_2 _21768_ (.A1(latched_branch),
    .A2(latched_store),
    .A3(\irq_state[1] ),
    .A4(\irq_state[0] ),
    .B1(_18291_),
    .X(_18292_));
 sky130_fd_sc_hd__buf_1 _21769_ (.A(_18292_),
    .X(_18293_));
 sky130_fd_sc_hd__buf_1 _21770_ (.A(_18293_),
    .X(_18294_));
 sky130_fd_sc_hd__o2111ai_2 _21771_ (.A1(_18276_),
    .A2(_18282_),
    .B1(_18286_),
    .C1(_18290_),
    .D1(_18294_),
    .Y(_18295_));
 sky130_fd_sc_hd__buf_1 _21772_ (.A(_18295_),
    .X(_18296_));
 sky130_fd_sc_hd__buf_1 _21773_ (.A(_18296_),
    .X(_18297_));
 sky130_fd_sc_hd__mux2_2 _21774_ (.A0(_18273_),
    .A1(\cpuregs[6][31] ),
    .S(_18297_),
    .X(_03727_));
 sky130_fd_sc_hd__buf_1 _21775_ (.A(\cpuregs_wrdata[30] ),
    .X(_18298_));
 sky130_fd_sc_hd__buf_1 _21776_ (.A(_18298_),
    .X(_18299_));
 sky130_fd_sc_hd__mux2_2 _21777_ (.A0(_18299_),
    .A1(\cpuregs[6][30] ),
    .S(_18297_),
    .X(_03726_));
 sky130_fd_sc_hd__buf_1 _21778_ (.A(\cpuregs_wrdata[29] ),
    .X(_18300_));
 sky130_fd_sc_hd__buf_1 _21779_ (.A(_18300_),
    .X(_18301_));
 sky130_fd_sc_hd__mux2_2 _21780_ (.A0(_18301_),
    .A1(\cpuregs[6][29] ),
    .S(_18297_),
    .X(_03725_));
 sky130_fd_sc_hd__buf_1 _21781_ (.A(\cpuregs_wrdata[28] ),
    .X(_18302_));
 sky130_fd_sc_hd__buf_1 _21782_ (.A(_18302_),
    .X(_18303_));
 sky130_fd_sc_hd__mux2_2 _21783_ (.A0(_18303_),
    .A1(\cpuregs[6][28] ),
    .S(_18297_),
    .X(_03724_));
 sky130_fd_sc_hd__buf_1 _21784_ (.A(\cpuregs_wrdata[27] ),
    .X(_18304_));
 sky130_fd_sc_hd__buf_1 _21785_ (.A(_18304_),
    .X(_18305_));
 sky130_fd_sc_hd__buf_1 _21786_ (.A(_18296_),
    .X(_18306_));
 sky130_fd_sc_hd__mux2_2 _21787_ (.A0(_18305_),
    .A1(\cpuregs[6][27] ),
    .S(_18306_),
    .X(_03723_));
 sky130_fd_sc_hd__buf_1 _21788_ (.A(\cpuregs_wrdata[26] ),
    .X(_18307_));
 sky130_fd_sc_hd__buf_1 _21789_ (.A(_18307_),
    .X(_18308_));
 sky130_fd_sc_hd__mux2_2 _21790_ (.A0(_18308_),
    .A1(\cpuregs[6][26] ),
    .S(_18306_),
    .X(_03722_));
 sky130_fd_sc_hd__buf_1 _21791_ (.A(\cpuregs_wrdata[25] ),
    .X(_18309_));
 sky130_fd_sc_hd__buf_1 _21792_ (.A(_18309_),
    .X(_18310_));
 sky130_fd_sc_hd__mux2_2 _21793_ (.A0(_18310_),
    .A1(\cpuregs[6][25] ),
    .S(_18306_),
    .X(_03721_));
 sky130_fd_sc_hd__buf_1 _21794_ (.A(\cpuregs_wrdata[24] ),
    .X(_18311_));
 sky130_fd_sc_hd__buf_1 _21795_ (.A(_18311_),
    .X(_18312_));
 sky130_fd_sc_hd__mux2_2 _21796_ (.A0(_18312_),
    .A1(\cpuregs[6][24] ),
    .S(_18306_),
    .X(_03720_));
 sky130_fd_sc_hd__buf_1 _21797_ (.A(\cpuregs_wrdata[23] ),
    .X(_18313_));
 sky130_fd_sc_hd__buf_1 _21798_ (.A(_18313_),
    .X(_18314_));
 sky130_fd_sc_hd__buf_1 _21799_ (.A(_18296_),
    .X(_18315_));
 sky130_fd_sc_hd__mux2_2 _21800_ (.A0(_18314_),
    .A1(\cpuregs[6][23] ),
    .S(_18315_),
    .X(_03719_));
 sky130_fd_sc_hd__buf_1 _21801_ (.A(\cpuregs_wrdata[22] ),
    .X(_18316_));
 sky130_fd_sc_hd__buf_1 _21802_ (.A(_18316_),
    .X(_18317_));
 sky130_fd_sc_hd__mux2_2 _21803_ (.A0(_18317_),
    .A1(\cpuregs[6][22] ),
    .S(_18315_),
    .X(_03718_));
 sky130_fd_sc_hd__buf_1 _21804_ (.A(\cpuregs_wrdata[21] ),
    .X(_18318_));
 sky130_fd_sc_hd__buf_1 _21805_ (.A(_18318_),
    .X(_18319_));
 sky130_fd_sc_hd__mux2_2 _21806_ (.A0(_18319_),
    .A1(\cpuregs[6][21] ),
    .S(_18315_),
    .X(_03717_));
 sky130_fd_sc_hd__buf_1 _21807_ (.A(\cpuregs_wrdata[20] ),
    .X(_18320_));
 sky130_fd_sc_hd__buf_1 _21808_ (.A(_18320_),
    .X(_18321_));
 sky130_fd_sc_hd__mux2_2 _21809_ (.A0(_18321_),
    .A1(\cpuregs[6][20] ),
    .S(_18315_),
    .X(_03716_));
 sky130_fd_sc_hd__buf_1 _21810_ (.A(\cpuregs_wrdata[19] ),
    .X(_18322_));
 sky130_fd_sc_hd__buf_1 _21811_ (.A(_18322_),
    .X(_18323_));
 sky130_fd_sc_hd__buf_1 _21812_ (.A(_18296_),
    .X(_18324_));
 sky130_fd_sc_hd__mux2_2 _21813_ (.A0(_18323_),
    .A1(\cpuregs[6][19] ),
    .S(_18324_),
    .X(_03715_));
 sky130_fd_sc_hd__buf_1 _21814_ (.A(\cpuregs_wrdata[18] ),
    .X(_18325_));
 sky130_fd_sc_hd__buf_1 _21815_ (.A(_18325_),
    .X(_18326_));
 sky130_fd_sc_hd__mux2_2 _21816_ (.A0(_18326_),
    .A1(\cpuregs[6][18] ),
    .S(_18324_),
    .X(_03714_));
 sky130_fd_sc_hd__buf_1 _21817_ (.A(\cpuregs_wrdata[17] ),
    .X(_18327_));
 sky130_fd_sc_hd__buf_1 _21818_ (.A(_18327_),
    .X(_18328_));
 sky130_fd_sc_hd__mux2_2 _21819_ (.A0(_18328_),
    .A1(\cpuregs[6][17] ),
    .S(_18324_),
    .X(_03713_));
 sky130_fd_sc_hd__buf_1 _21820_ (.A(\cpuregs_wrdata[16] ),
    .X(_18329_));
 sky130_fd_sc_hd__buf_1 _21821_ (.A(_18329_),
    .X(_18330_));
 sky130_fd_sc_hd__mux2_2 _21822_ (.A0(_18330_),
    .A1(\cpuregs[6][16] ),
    .S(_18324_),
    .X(_03712_));
 sky130_fd_sc_hd__buf_1 _21823_ (.A(\cpuregs_wrdata[15] ),
    .X(_18331_));
 sky130_fd_sc_hd__buf_1 _21824_ (.A(_18331_),
    .X(_18332_));
 sky130_fd_sc_hd__buf_1 _21825_ (.A(_18295_),
    .X(_18333_));
 sky130_fd_sc_hd__buf_1 _21826_ (.A(_18333_),
    .X(_18334_));
 sky130_fd_sc_hd__mux2_2 _21827_ (.A0(_18332_),
    .A1(\cpuregs[6][15] ),
    .S(_18334_),
    .X(_03711_));
 sky130_fd_sc_hd__buf_1 _21828_ (.A(\cpuregs_wrdata[14] ),
    .X(_18335_));
 sky130_fd_sc_hd__buf_1 _21829_ (.A(_18335_),
    .X(_18336_));
 sky130_fd_sc_hd__mux2_2 _21830_ (.A0(_18336_),
    .A1(\cpuregs[6][14] ),
    .S(_18334_),
    .X(_03710_));
 sky130_fd_sc_hd__buf_1 _21831_ (.A(\cpuregs_wrdata[13] ),
    .X(_18337_));
 sky130_fd_sc_hd__buf_1 _21832_ (.A(_18337_),
    .X(_18338_));
 sky130_fd_sc_hd__mux2_2 _21833_ (.A0(_18338_),
    .A1(\cpuregs[6][13] ),
    .S(_18334_),
    .X(_03709_));
 sky130_fd_sc_hd__buf_1 _21834_ (.A(\cpuregs_wrdata[12] ),
    .X(_18339_));
 sky130_fd_sc_hd__buf_1 _21835_ (.A(_18339_),
    .X(_18340_));
 sky130_fd_sc_hd__mux2_2 _21836_ (.A0(_18340_),
    .A1(\cpuregs[6][12] ),
    .S(_18334_),
    .X(_03708_));
 sky130_fd_sc_hd__buf_1 _21837_ (.A(\cpuregs_wrdata[11] ),
    .X(_18341_));
 sky130_fd_sc_hd__buf_1 _21838_ (.A(_18341_),
    .X(_18342_));
 sky130_fd_sc_hd__buf_1 _21839_ (.A(_18333_),
    .X(_18343_));
 sky130_fd_sc_hd__mux2_2 _21840_ (.A0(_18342_),
    .A1(\cpuregs[6][11] ),
    .S(_18343_),
    .X(_03707_));
 sky130_fd_sc_hd__buf_1 _21841_ (.A(\cpuregs_wrdata[10] ),
    .X(_18344_));
 sky130_fd_sc_hd__buf_1 _21842_ (.A(_18344_),
    .X(_18345_));
 sky130_fd_sc_hd__mux2_2 _21843_ (.A0(_18345_),
    .A1(\cpuregs[6][10] ),
    .S(_18343_),
    .X(_03706_));
 sky130_fd_sc_hd__buf_1 _21844_ (.A(\cpuregs_wrdata[9] ),
    .X(_18346_));
 sky130_fd_sc_hd__buf_1 _21845_ (.A(_18346_),
    .X(_18347_));
 sky130_fd_sc_hd__mux2_2 _21846_ (.A0(_18347_),
    .A1(\cpuregs[6][9] ),
    .S(_18343_),
    .X(_03705_));
 sky130_fd_sc_hd__buf_1 _21847_ (.A(\cpuregs_wrdata[8] ),
    .X(_18348_));
 sky130_fd_sc_hd__buf_1 _21848_ (.A(_18348_),
    .X(_18349_));
 sky130_fd_sc_hd__mux2_2 _21849_ (.A0(_18349_),
    .A1(\cpuregs[6][8] ),
    .S(_18343_),
    .X(_03704_));
 sky130_fd_sc_hd__buf_1 _21850_ (.A(\cpuregs_wrdata[7] ),
    .X(_18350_));
 sky130_fd_sc_hd__buf_1 _21851_ (.A(_18350_),
    .X(_18351_));
 sky130_fd_sc_hd__buf_1 _21852_ (.A(_18333_),
    .X(_18352_));
 sky130_fd_sc_hd__mux2_2 _21853_ (.A0(_18351_),
    .A1(\cpuregs[6][7] ),
    .S(_18352_),
    .X(_03703_));
 sky130_fd_sc_hd__buf_1 _21854_ (.A(\cpuregs_wrdata[6] ),
    .X(_18353_));
 sky130_fd_sc_hd__buf_1 _21855_ (.A(_18353_),
    .X(_18354_));
 sky130_fd_sc_hd__mux2_2 _21856_ (.A0(_18354_),
    .A1(\cpuregs[6][6] ),
    .S(_18352_),
    .X(_03702_));
 sky130_fd_sc_hd__buf_1 _21857_ (.A(\cpuregs_wrdata[5] ),
    .X(_18355_));
 sky130_fd_sc_hd__buf_1 _21858_ (.A(_18355_),
    .X(_18356_));
 sky130_fd_sc_hd__mux2_2 _21859_ (.A0(_18356_),
    .A1(\cpuregs[6][5] ),
    .S(_18352_),
    .X(_03701_));
 sky130_fd_sc_hd__buf_1 _21860_ (.A(\cpuregs_wrdata[4] ),
    .X(_18357_));
 sky130_fd_sc_hd__buf_1 _21861_ (.A(_18357_),
    .X(_18358_));
 sky130_fd_sc_hd__mux2_2 _21862_ (.A0(_18358_),
    .A1(\cpuregs[6][4] ),
    .S(_18352_),
    .X(_03700_));
 sky130_fd_sc_hd__buf_1 _21863_ (.A(\cpuregs_wrdata[3] ),
    .X(_18359_));
 sky130_fd_sc_hd__buf_1 _21864_ (.A(_18359_),
    .X(_18360_));
 sky130_fd_sc_hd__buf_1 _21865_ (.A(_18333_),
    .X(_18361_));
 sky130_fd_sc_hd__mux2_2 _21866_ (.A0(_18360_),
    .A1(\cpuregs[6][3] ),
    .S(_18361_),
    .X(_03699_));
 sky130_fd_sc_hd__buf_1 _21867_ (.A(\cpuregs_wrdata[2] ),
    .X(_18362_));
 sky130_fd_sc_hd__buf_1 _21868_ (.A(_18362_),
    .X(_18363_));
 sky130_fd_sc_hd__mux2_2 _21869_ (.A0(_18363_),
    .A1(\cpuregs[6][2] ),
    .S(_18361_),
    .X(_03698_));
 sky130_fd_sc_hd__buf_1 _21870_ (.A(\cpuregs_wrdata[1] ),
    .X(_18364_));
 sky130_fd_sc_hd__buf_1 _21871_ (.A(_18364_),
    .X(_18365_));
 sky130_fd_sc_hd__mux2_2 _21872_ (.A0(_18365_),
    .A1(\cpuregs[6][1] ),
    .S(_18361_),
    .X(_03697_));
 sky130_fd_sc_hd__buf_1 _21873_ (.A(\cpuregs_wrdata[0] ),
    .X(_18366_));
 sky130_fd_sc_hd__buf_1 _21874_ (.A(_18366_),
    .X(_18367_));
 sky130_fd_sc_hd__mux2_2 _21875_ (.A0(_18367_),
    .A1(\cpuregs[6][0] ),
    .S(_18361_),
    .X(_03696_));
 sky130_fd_sc_hd__nor3b_2 _21876_ (.A(_18287_),
    .B(_18289_),
    .C_N(_18288_),
    .Y(_18368_));
 sky130_fd_sc_hd__and2b_2 _21877_ (.A_N(_18284_),
    .B(_18283_),
    .X(_18369_));
 sky130_fd_sc_hd__buf_1 _21878_ (.A(_18369_),
    .X(_18370_));
 sky130_fd_sc_hd__o2111ai_2 _21879_ (.A1(_18276_),
    .A2(_18282_),
    .B1(_18368_),
    .C1(_18370_),
    .D1(_18294_),
    .Y(_18371_));
 sky130_fd_sc_hd__buf_1 _21880_ (.A(_18371_),
    .X(_18372_));
 sky130_fd_sc_hd__buf_1 _21881_ (.A(_18372_),
    .X(_18373_));
 sky130_fd_sc_hd__mux2_2 _21882_ (.A0(_18273_),
    .A1(\cpuregs[9][31] ),
    .S(_18373_),
    .X(_03695_));
 sky130_fd_sc_hd__mux2_2 _21883_ (.A0(_18299_),
    .A1(\cpuregs[9][30] ),
    .S(_18373_),
    .X(_03694_));
 sky130_fd_sc_hd__mux2_2 _21884_ (.A0(_18301_),
    .A1(\cpuregs[9][29] ),
    .S(_18373_),
    .X(_03693_));
 sky130_fd_sc_hd__mux2_2 _21885_ (.A0(_18303_),
    .A1(\cpuregs[9][28] ),
    .S(_18373_),
    .X(_03692_));
 sky130_fd_sc_hd__buf_1 _21886_ (.A(_18372_),
    .X(_18374_));
 sky130_fd_sc_hd__mux2_2 _21887_ (.A0(_18305_),
    .A1(\cpuregs[9][27] ),
    .S(_18374_),
    .X(_03691_));
 sky130_fd_sc_hd__mux2_2 _21888_ (.A0(_18308_),
    .A1(\cpuregs[9][26] ),
    .S(_18374_),
    .X(_03690_));
 sky130_fd_sc_hd__mux2_2 _21889_ (.A0(_18310_),
    .A1(\cpuregs[9][25] ),
    .S(_18374_),
    .X(_03689_));
 sky130_fd_sc_hd__mux2_2 _21890_ (.A0(_18312_),
    .A1(\cpuregs[9][24] ),
    .S(_18374_),
    .X(_03688_));
 sky130_fd_sc_hd__buf_1 _21891_ (.A(_18372_),
    .X(_18375_));
 sky130_fd_sc_hd__mux2_2 _21892_ (.A0(_18314_),
    .A1(\cpuregs[9][23] ),
    .S(_18375_),
    .X(_03687_));
 sky130_fd_sc_hd__mux2_2 _21893_ (.A0(_18317_),
    .A1(\cpuregs[9][22] ),
    .S(_18375_),
    .X(_03686_));
 sky130_fd_sc_hd__mux2_2 _21894_ (.A0(_18319_),
    .A1(\cpuregs[9][21] ),
    .S(_18375_),
    .X(_03685_));
 sky130_fd_sc_hd__mux2_2 _21895_ (.A0(_18321_),
    .A1(\cpuregs[9][20] ),
    .S(_18375_),
    .X(_03684_));
 sky130_fd_sc_hd__buf_1 _21896_ (.A(_18372_),
    .X(_18376_));
 sky130_fd_sc_hd__mux2_2 _21897_ (.A0(_18323_),
    .A1(\cpuregs[9][19] ),
    .S(_18376_),
    .X(_03683_));
 sky130_fd_sc_hd__mux2_2 _21898_ (.A0(_18326_),
    .A1(\cpuregs[9][18] ),
    .S(_18376_),
    .X(_03682_));
 sky130_fd_sc_hd__mux2_2 _21899_ (.A0(_18328_),
    .A1(\cpuregs[9][17] ),
    .S(_18376_),
    .X(_03681_));
 sky130_fd_sc_hd__mux2_2 _21900_ (.A0(_18330_),
    .A1(\cpuregs[9][16] ),
    .S(_18376_),
    .X(_03680_));
 sky130_fd_sc_hd__buf_1 _21901_ (.A(_18371_),
    .X(_18377_));
 sky130_fd_sc_hd__buf_1 _21902_ (.A(_18377_),
    .X(_18378_));
 sky130_fd_sc_hd__mux2_2 _21903_ (.A0(_18332_),
    .A1(\cpuregs[9][15] ),
    .S(_18378_),
    .X(_03679_));
 sky130_fd_sc_hd__mux2_2 _21904_ (.A0(_18336_),
    .A1(\cpuregs[9][14] ),
    .S(_18378_),
    .X(_03678_));
 sky130_fd_sc_hd__mux2_2 _21905_ (.A0(_18338_),
    .A1(\cpuregs[9][13] ),
    .S(_18378_),
    .X(_03677_));
 sky130_fd_sc_hd__mux2_2 _21906_ (.A0(_18340_),
    .A1(\cpuregs[9][12] ),
    .S(_18378_),
    .X(_03676_));
 sky130_fd_sc_hd__buf_1 _21907_ (.A(_18377_),
    .X(_18379_));
 sky130_fd_sc_hd__mux2_2 _21908_ (.A0(_18342_),
    .A1(\cpuregs[9][11] ),
    .S(_18379_),
    .X(_03675_));
 sky130_fd_sc_hd__mux2_2 _21909_ (.A0(_18345_),
    .A1(\cpuregs[9][10] ),
    .S(_18379_),
    .X(_03674_));
 sky130_fd_sc_hd__mux2_2 _21910_ (.A0(_18347_),
    .A1(\cpuregs[9][9] ),
    .S(_18379_),
    .X(_03673_));
 sky130_fd_sc_hd__mux2_2 _21911_ (.A0(_18349_),
    .A1(\cpuregs[9][8] ),
    .S(_18379_),
    .X(_03672_));
 sky130_fd_sc_hd__buf_1 _21912_ (.A(_18377_),
    .X(_18380_));
 sky130_fd_sc_hd__mux2_2 _21913_ (.A0(_18351_),
    .A1(\cpuregs[9][7] ),
    .S(_18380_),
    .X(_03671_));
 sky130_fd_sc_hd__mux2_2 _21914_ (.A0(_18354_),
    .A1(\cpuregs[9][6] ),
    .S(_18380_),
    .X(_03670_));
 sky130_fd_sc_hd__mux2_2 _21915_ (.A0(_18356_),
    .A1(\cpuregs[9][5] ),
    .S(_18380_),
    .X(_03669_));
 sky130_fd_sc_hd__mux2_2 _21916_ (.A0(_18358_),
    .A1(\cpuregs[9][4] ),
    .S(_18380_),
    .X(_03668_));
 sky130_fd_sc_hd__buf_1 _21917_ (.A(_18377_),
    .X(_18381_));
 sky130_fd_sc_hd__mux2_2 _21918_ (.A0(_18360_),
    .A1(\cpuregs[9][3] ),
    .S(_18381_),
    .X(_03667_));
 sky130_fd_sc_hd__mux2_2 _21919_ (.A0(_18363_),
    .A1(\cpuregs[9][2] ),
    .S(_18381_),
    .X(_03666_));
 sky130_fd_sc_hd__mux2_2 _21920_ (.A0(_18365_),
    .A1(\cpuregs[9][1] ),
    .S(_18381_),
    .X(_03665_));
 sky130_fd_sc_hd__mux2_2 _21921_ (.A0(_18367_),
    .A1(\cpuregs[9][0] ),
    .S(_18381_),
    .X(_03664_));
 sky130_fd_sc_hd__buf_1 _21922_ (.A(_17221_),
    .X(_18382_));
 sky130_fd_sc_hd__o21ai_2 _21923_ (.A1(_16828_),
    .A2(_17017_),
    .B1(_18382_),
    .Y(_18383_));
 sky130_fd_sc_hd__buf_1 _21924_ (.A(_18383_),
    .X(_18384_));
 sky130_fd_sc_hd__mux2_2 _21925_ (.A0(_02467_),
    .A1(_16978_),
    .S(_18384_),
    .X(_03663_));
 sky130_fd_sc_hd__buf_1 _21926_ (.A(pcpi_rs2[30]),
    .X(_18385_));
 sky130_fd_sc_hd__mux2_2 _21927_ (.A0(_02466_),
    .A1(_18385_),
    .S(_18384_),
    .X(_03662_));
 sky130_fd_sc_hd__buf_1 _21928_ (.A(pcpi_rs2[29]),
    .X(_18386_));
 sky130_fd_sc_hd__buf_1 _21929_ (.A(_18386_),
    .X(_18387_));
 sky130_fd_sc_hd__mux2_2 _21930_ (.A0(_02464_),
    .A1(_18387_),
    .S(_18384_),
    .X(_03661_));
 sky130_fd_sc_hd__buf_1 _21931_ (.A(pcpi_rs2[28]),
    .X(_18388_));
 sky130_fd_sc_hd__buf_1 _21932_ (.A(_18383_),
    .X(_18389_));
 sky130_fd_sc_hd__buf_1 _21933_ (.A(_18389_),
    .X(_18390_));
 sky130_fd_sc_hd__mux2_2 _21934_ (.A0(_02463_),
    .A1(_18388_),
    .S(_18390_),
    .X(_03660_));
 sky130_fd_sc_hd__buf_1 _21935_ (.A(pcpi_rs2[27]),
    .X(_18391_));
 sky130_fd_sc_hd__mux2_2 _21936_ (.A0(_02462_),
    .A1(_18391_),
    .S(_18390_),
    .X(_03659_));
 sky130_fd_sc_hd__buf_1 _21937_ (.A(pcpi_rs2[26]),
    .X(_18392_));
 sky130_fd_sc_hd__buf_1 _21938_ (.A(_18392_),
    .X(_18393_));
 sky130_fd_sc_hd__mux2_2 _21939_ (.A0(_02461_),
    .A1(_18393_),
    .S(_18390_),
    .X(_03658_));
 sky130_fd_sc_hd__buf_1 _21940_ (.A(pcpi_rs2[25]),
    .X(_18394_));
 sky130_fd_sc_hd__buf_1 _21941_ (.A(_18394_),
    .X(_18395_));
 sky130_fd_sc_hd__mux2_2 _21942_ (.A0(_02460_),
    .A1(_18395_),
    .S(_18390_),
    .X(_03657_));
 sky130_fd_sc_hd__buf_1 _21943_ (.A(pcpi_rs2[24]),
    .X(_18396_));
 sky130_fd_sc_hd__buf_1 _21944_ (.A(_18389_),
    .X(_18397_));
 sky130_fd_sc_hd__mux2_2 _21945_ (.A0(_02459_),
    .A1(_18396_),
    .S(_18397_),
    .X(_03656_));
 sky130_fd_sc_hd__buf_1 _21946_ (.A(pcpi_rs2[23]),
    .X(_18398_));
 sky130_fd_sc_hd__buf_1 _21947_ (.A(_18398_),
    .X(_18399_));
 sky130_fd_sc_hd__mux2_2 _21948_ (.A0(_02458_),
    .A1(_18399_),
    .S(_18397_),
    .X(_03655_));
 sky130_fd_sc_hd__buf_1 _21949_ (.A(pcpi_rs2[22]),
    .X(_18400_));
 sky130_fd_sc_hd__buf_1 _21950_ (.A(_18400_),
    .X(_18401_));
 sky130_fd_sc_hd__mux2_2 _21951_ (.A0(_02457_),
    .A1(_18401_),
    .S(_18397_),
    .X(_03654_));
 sky130_fd_sc_hd__buf_1 _21952_ (.A(pcpi_rs2[21]),
    .X(_18402_));
 sky130_fd_sc_hd__buf_1 _21953_ (.A(_18402_),
    .X(_18403_));
 sky130_fd_sc_hd__mux2_2 _21954_ (.A0(_02456_),
    .A1(_18403_),
    .S(_18397_),
    .X(_03653_));
 sky130_fd_sc_hd__buf_1 _21955_ (.A(pcpi_rs2[20]),
    .X(_18404_));
 sky130_fd_sc_hd__buf_1 _21956_ (.A(_18389_),
    .X(_18405_));
 sky130_fd_sc_hd__mux2_2 _21957_ (.A0(_02455_),
    .A1(_18404_),
    .S(_18405_),
    .X(_03652_));
 sky130_fd_sc_hd__buf_1 _21958_ (.A(pcpi_rs2[19]),
    .X(_18406_));
 sky130_fd_sc_hd__buf_1 _21959_ (.A(_18406_),
    .X(_18407_));
 sky130_fd_sc_hd__mux2_2 _21960_ (.A0(_02453_),
    .A1(_18407_),
    .S(_18405_),
    .X(_03651_));
 sky130_fd_sc_hd__buf_1 _21961_ (.A(pcpi_rs2[18]),
    .X(_18408_));
 sky130_fd_sc_hd__buf_1 _21962_ (.A(_18408_),
    .X(_18409_));
 sky130_fd_sc_hd__mux2_2 _21963_ (.A0(_02452_),
    .A1(_18409_),
    .S(_18405_),
    .X(_03650_));
 sky130_fd_sc_hd__buf_1 _21964_ (.A(pcpi_rs2[17]),
    .X(_18410_));
 sky130_fd_sc_hd__buf_1 _21965_ (.A(_18410_),
    .X(_18411_));
 sky130_fd_sc_hd__mux2_2 _21966_ (.A0(_02451_),
    .A1(_18411_),
    .S(_18405_),
    .X(_03649_));
 sky130_fd_sc_hd__buf_1 _21967_ (.A(pcpi_rs2[16]),
    .X(_18412_));
 sky130_fd_sc_hd__buf_1 _21968_ (.A(_18383_),
    .X(_18413_));
 sky130_fd_sc_hd__buf_1 _21969_ (.A(_18413_),
    .X(_18414_));
 sky130_fd_sc_hd__mux2_2 _21970_ (.A0(_02450_),
    .A1(_18412_),
    .S(_18414_),
    .X(_03648_));
 sky130_fd_sc_hd__buf_1 _21971_ (.A(pcpi_rs2[15]),
    .X(_18415_));
 sky130_fd_sc_hd__buf_1 _21972_ (.A(_18415_),
    .X(_18416_));
 sky130_fd_sc_hd__mux2_2 _21973_ (.A0(_02449_),
    .A1(_18416_),
    .S(_18414_),
    .X(_03647_));
 sky130_fd_sc_hd__buf_1 _21974_ (.A(pcpi_rs2[14]),
    .X(_18417_));
 sky130_fd_sc_hd__buf_1 _21975_ (.A(_18417_),
    .X(_18418_));
 sky130_fd_sc_hd__mux2_2 _21976_ (.A0(_02448_),
    .A1(_18418_),
    .S(_18414_),
    .X(_03646_));
 sky130_fd_sc_hd__buf_1 _21977_ (.A(pcpi_rs2[13]),
    .X(_18419_));
 sky130_fd_sc_hd__buf_1 _21978_ (.A(_18419_),
    .X(_18420_));
 sky130_fd_sc_hd__mux2_2 _21979_ (.A0(_02447_),
    .A1(_18420_),
    .S(_18414_),
    .X(_03645_));
 sky130_fd_sc_hd__buf_1 _21980_ (.A(pcpi_rs2[12]),
    .X(_18421_));
 sky130_fd_sc_hd__buf_1 _21981_ (.A(_18413_),
    .X(_18422_));
 sky130_fd_sc_hd__mux2_2 _21982_ (.A0(_02446_),
    .A1(_18421_),
    .S(_18422_),
    .X(_03644_));
 sky130_fd_sc_hd__buf_1 _21983_ (.A(pcpi_rs2[11]),
    .X(_18423_));
 sky130_fd_sc_hd__buf_1 _21984_ (.A(_18423_),
    .X(_18424_));
 sky130_fd_sc_hd__mux2_2 _21985_ (.A0(_02445_),
    .A1(_18424_),
    .S(_18422_),
    .X(_03643_));
 sky130_fd_sc_hd__buf_1 _21986_ (.A(pcpi_rs2[10]),
    .X(_18425_));
 sky130_fd_sc_hd__buf_1 _21987_ (.A(_18425_),
    .X(_18426_));
 sky130_fd_sc_hd__mux2_2 _21988_ (.A0(_02444_),
    .A1(_18426_),
    .S(_18422_),
    .X(_03642_));
 sky130_fd_sc_hd__buf_1 _21989_ (.A(pcpi_rs2[9]),
    .X(_18427_));
 sky130_fd_sc_hd__buf_1 _21990_ (.A(_18427_),
    .X(_18428_));
 sky130_fd_sc_hd__mux2_2 _21991_ (.A0(_02474_),
    .A1(_18428_),
    .S(_18422_),
    .X(_03641_));
 sky130_fd_sc_hd__buf_1 _21992_ (.A(pcpi_rs2[8]),
    .X(_18429_));
 sky130_fd_sc_hd__buf_1 _21993_ (.A(_18429_),
    .X(_18430_));
 sky130_fd_sc_hd__buf_1 _21994_ (.A(_18413_),
    .X(_18431_));
 sky130_fd_sc_hd__mux2_2 _21995_ (.A0(_02473_),
    .A1(_18430_),
    .S(_18431_),
    .X(_03640_));
 sky130_fd_sc_hd__buf_1 _21996_ (.A(mem_la_wdata[7]),
    .X(_18432_));
 sky130_fd_sc_hd__buf_1 _21997_ (.A(_18432_),
    .X(_18433_));
 sky130_fd_sc_hd__buf_1 _21998_ (.A(_18433_),
    .X(_18434_));
 sky130_fd_sc_hd__mux2_2 _21999_ (.A0(_02472_),
    .A1(_18434_),
    .S(_18431_),
    .X(_03639_));
 sky130_fd_sc_hd__buf_1 _22000_ (.A(mem_la_wdata[6]),
    .X(_18435_));
 sky130_fd_sc_hd__buf_1 _22001_ (.A(_18435_),
    .X(_18436_));
 sky130_fd_sc_hd__buf_1 _22002_ (.A(_18436_),
    .X(_18437_));
 sky130_fd_sc_hd__mux2_2 _22003_ (.A0(_02471_),
    .A1(_18437_),
    .S(_18431_),
    .X(_03638_));
 sky130_fd_sc_hd__buf_1 _22004_ (.A(mem_la_wdata[5]),
    .X(_18438_));
 sky130_fd_sc_hd__buf_1 _22005_ (.A(_18438_),
    .X(_18439_));
 sky130_fd_sc_hd__buf_1 _22006_ (.A(_18439_),
    .X(_18440_));
 sky130_fd_sc_hd__mux2_2 _22007_ (.A0(_02470_),
    .A1(_18440_),
    .S(_18431_),
    .X(_03637_));
 sky130_fd_sc_hd__buf_1 _22008_ (.A(mem_la_wdata[4]),
    .X(_18441_));
 sky130_fd_sc_hd__buf_1 _22009_ (.A(_18441_),
    .X(_18442_));
 sky130_fd_sc_hd__buf_1 _22010_ (.A(_18413_),
    .X(_18443_));
 sky130_fd_sc_hd__mux2_2 _22011_ (.A0(_02469_),
    .A1(_18442_),
    .S(_18443_),
    .X(_03636_));
 sky130_fd_sc_hd__buf_1 _22012_ (.A(mem_la_wdata[3]),
    .X(_18444_));
 sky130_fd_sc_hd__buf_1 _22013_ (.A(_18444_),
    .X(_18445_));
 sky130_fd_sc_hd__buf_1 _22014_ (.A(_18445_),
    .X(_18446_));
 sky130_fd_sc_hd__mux2_2 _22015_ (.A0(_02468_),
    .A1(_18446_),
    .S(_18443_),
    .X(_03635_));
 sky130_fd_sc_hd__buf_1 _22016_ (.A(mem_la_wdata[2]),
    .X(_18447_));
 sky130_fd_sc_hd__buf_1 _22017_ (.A(_18447_),
    .X(_18448_));
 sky130_fd_sc_hd__mux2_2 _22018_ (.A0(_02465_),
    .A1(_18448_),
    .S(_18443_),
    .X(_03634_));
 sky130_fd_sc_hd__buf_1 _22019_ (.A(mem_la_wdata[1]),
    .X(_18449_));
 sky130_fd_sc_hd__buf_1 _22020_ (.A(_18449_),
    .X(_18450_));
 sky130_fd_sc_hd__buf_1 _22021_ (.A(_18450_),
    .X(_18451_));
 sky130_fd_sc_hd__mux2_2 _22022_ (.A0(_02454_),
    .A1(_18451_),
    .S(_18443_),
    .X(_03633_));
 sky130_fd_sc_hd__buf_1 _22023_ (.A(mem_la_wdata[0]),
    .X(_18452_));
 sky130_fd_sc_hd__buf_1 _22024_ (.A(_18452_),
    .X(_18453_));
 sky130_fd_sc_hd__buf_1 _22025_ (.A(_18453_),
    .X(_18454_));
 sky130_fd_sc_hd__buf_1 _22026_ (.A(_18454_),
    .X(_18455_));
 sky130_fd_sc_hd__mux2_2 _22027_ (.A0(_02443_),
    .A1(_18455_),
    .S(_18389_),
    .X(_03632_));
 sky130_fd_sc_hd__buf_1 _22028_ (.A(\cpuregs_wrdata[31] ),
    .X(_18456_));
 sky130_fd_sc_hd__o21a_2 _22029_ (.A1(_18274_),
    .A2(_18279_),
    .B1(_18292_),
    .X(_18457_));
 sky130_fd_sc_hd__buf_1 _22030_ (.A(_18457_),
    .X(_18458_));
 sky130_fd_sc_hd__and3b_2 _22031_ (.A_N(_18276_),
    .B(_18458_),
    .C(_18290_),
    .X(_18459_));
 sky130_fd_sc_hd__buf_1 _22032_ (.A(_18459_),
    .X(_18460_));
 sky130_fd_sc_hd__buf_1 _22033_ (.A(_18460_),
    .X(_18461_));
 sky130_fd_sc_hd__mux2_2 _22034_ (.A0(\cpuregs[4][31] ),
    .A1(_18456_),
    .S(_18461_),
    .X(_03631_));
 sky130_fd_sc_hd__buf_1 _22035_ (.A(\cpuregs_wrdata[30] ),
    .X(_18462_));
 sky130_fd_sc_hd__mux2_2 _22036_ (.A0(\cpuregs[4][30] ),
    .A1(_18462_),
    .S(_18461_),
    .X(_03630_));
 sky130_fd_sc_hd__buf_1 _22037_ (.A(\cpuregs_wrdata[29] ),
    .X(_18463_));
 sky130_fd_sc_hd__mux2_2 _22038_ (.A0(\cpuregs[4][29] ),
    .A1(_18463_),
    .S(_18461_),
    .X(_03629_));
 sky130_fd_sc_hd__buf_1 _22039_ (.A(\cpuregs_wrdata[28] ),
    .X(_18464_));
 sky130_fd_sc_hd__mux2_2 _22040_ (.A0(\cpuregs[4][28] ),
    .A1(_18464_),
    .S(_18461_),
    .X(_03628_));
 sky130_fd_sc_hd__buf_1 _22041_ (.A(\cpuregs_wrdata[27] ),
    .X(_18465_));
 sky130_fd_sc_hd__buf_1 _22042_ (.A(_18460_),
    .X(_18466_));
 sky130_fd_sc_hd__mux2_2 _22043_ (.A0(\cpuregs[4][27] ),
    .A1(_18465_),
    .S(_18466_),
    .X(_03627_));
 sky130_fd_sc_hd__buf_1 _22044_ (.A(\cpuregs_wrdata[26] ),
    .X(_18467_));
 sky130_fd_sc_hd__mux2_2 _22045_ (.A0(\cpuregs[4][26] ),
    .A1(_18467_),
    .S(_18466_),
    .X(_03626_));
 sky130_fd_sc_hd__buf_1 _22046_ (.A(\cpuregs_wrdata[25] ),
    .X(_18468_));
 sky130_fd_sc_hd__mux2_2 _22047_ (.A0(\cpuregs[4][25] ),
    .A1(_18468_),
    .S(_18466_),
    .X(_03625_));
 sky130_fd_sc_hd__buf_1 _22048_ (.A(\cpuregs_wrdata[24] ),
    .X(_18469_));
 sky130_fd_sc_hd__mux2_2 _22049_ (.A0(\cpuregs[4][24] ),
    .A1(_18469_),
    .S(_18466_),
    .X(_03624_));
 sky130_fd_sc_hd__buf_1 _22050_ (.A(\cpuregs_wrdata[23] ),
    .X(_18470_));
 sky130_fd_sc_hd__buf_1 _22051_ (.A(_18460_),
    .X(_18471_));
 sky130_fd_sc_hd__mux2_2 _22052_ (.A0(\cpuregs[4][23] ),
    .A1(_18470_),
    .S(_18471_),
    .X(_03623_));
 sky130_fd_sc_hd__buf_1 _22053_ (.A(\cpuregs_wrdata[22] ),
    .X(_18472_));
 sky130_fd_sc_hd__mux2_2 _22054_ (.A0(\cpuregs[4][22] ),
    .A1(_18472_),
    .S(_18471_),
    .X(_03622_));
 sky130_fd_sc_hd__buf_1 _22055_ (.A(\cpuregs_wrdata[21] ),
    .X(_18473_));
 sky130_fd_sc_hd__mux2_2 _22056_ (.A0(\cpuregs[4][21] ),
    .A1(_18473_),
    .S(_18471_),
    .X(_03621_));
 sky130_fd_sc_hd__buf_1 _22057_ (.A(\cpuregs_wrdata[20] ),
    .X(_18474_));
 sky130_fd_sc_hd__mux2_2 _22058_ (.A0(\cpuregs[4][20] ),
    .A1(_18474_),
    .S(_18471_),
    .X(_03620_));
 sky130_fd_sc_hd__buf_1 _22059_ (.A(\cpuregs_wrdata[19] ),
    .X(_18475_));
 sky130_fd_sc_hd__buf_1 _22060_ (.A(_18460_),
    .X(_18476_));
 sky130_fd_sc_hd__mux2_2 _22061_ (.A0(\cpuregs[4][19] ),
    .A1(_18475_),
    .S(_18476_),
    .X(_03619_));
 sky130_fd_sc_hd__buf_1 _22062_ (.A(\cpuregs_wrdata[18] ),
    .X(_18477_));
 sky130_fd_sc_hd__mux2_2 _22063_ (.A0(\cpuregs[4][18] ),
    .A1(_18477_),
    .S(_18476_),
    .X(_03618_));
 sky130_fd_sc_hd__buf_1 _22064_ (.A(\cpuregs_wrdata[17] ),
    .X(_18478_));
 sky130_fd_sc_hd__mux2_2 _22065_ (.A0(\cpuregs[4][17] ),
    .A1(_18478_),
    .S(_18476_),
    .X(_03617_));
 sky130_fd_sc_hd__buf_1 _22066_ (.A(\cpuregs_wrdata[16] ),
    .X(_18479_));
 sky130_fd_sc_hd__mux2_2 _22067_ (.A0(\cpuregs[4][16] ),
    .A1(_18479_),
    .S(_18476_),
    .X(_03616_));
 sky130_fd_sc_hd__buf_1 _22068_ (.A(\cpuregs_wrdata[15] ),
    .X(_18480_));
 sky130_fd_sc_hd__buf_1 _22069_ (.A(_18459_),
    .X(_18481_));
 sky130_fd_sc_hd__buf_1 _22070_ (.A(_18481_),
    .X(_18482_));
 sky130_fd_sc_hd__mux2_2 _22071_ (.A0(\cpuregs[4][15] ),
    .A1(_18480_),
    .S(_18482_),
    .X(_03615_));
 sky130_fd_sc_hd__buf_1 _22072_ (.A(\cpuregs_wrdata[14] ),
    .X(_18483_));
 sky130_fd_sc_hd__mux2_2 _22073_ (.A0(\cpuregs[4][14] ),
    .A1(_18483_),
    .S(_18482_),
    .X(_03614_));
 sky130_fd_sc_hd__buf_1 _22074_ (.A(\cpuregs_wrdata[13] ),
    .X(_18484_));
 sky130_fd_sc_hd__mux2_2 _22075_ (.A0(\cpuregs[4][13] ),
    .A1(_18484_),
    .S(_18482_),
    .X(_03613_));
 sky130_fd_sc_hd__buf_1 _22076_ (.A(\cpuregs_wrdata[12] ),
    .X(_18485_));
 sky130_fd_sc_hd__mux2_2 _22077_ (.A0(\cpuregs[4][12] ),
    .A1(_18485_),
    .S(_18482_),
    .X(_03612_));
 sky130_fd_sc_hd__buf_1 _22078_ (.A(\cpuregs_wrdata[11] ),
    .X(_18486_));
 sky130_fd_sc_hd__buf_1 _22079_ (.A(_18481_),
    .X(_18487_));
 sky130_fd_sc_hd__mux2_2 _22080_ (.A0(\cpuregs[4][11] ),
    .A1(_18486_),
    .S(_18487_),
    .X(_03611_));
 sky130_fd_sc_hd__buf_1 _22081_ (.A(\cpuregs_wrdata[10] ),
    .X(_18488_));
 sky130_fd_sc_hd__mux2_2 _22082_ (.A0(\cpuregs[4][10] ),
    .A1(_18488_),
    .S(_18487_),
    .X(_03610_));
 sky130_fd_sc_hd__buf_1 _22083_ (.A(\cpuregs_wrdata[9] ),
    .X(_18489_));
 sky130_fd_sc_hd__mux2_2 _22084_ (.A0(\cpuregs[4][9] ),
    .A1(_18489_),
    .S(_18487_),
    .X(_03609_));
 sky130_fd_sc_hd__buf_1 _22085_ (.A(\cpuregs_wrdata[8] ),
    .X(_18490_));
 sky130_fd_sc_hd__mux2_2 _22086_ (.A0(\cpuregs[4][8] ),
    .A1(_18490_),
    .S(_18487_),
    .X(_03608_));
 sky130_fd_sc_hd__buf_1 _22087_ (.A(\cpuregs_wrdata[7] ),
    .X(_18491_));
 sky130_fd_sc_hd__buf_1 _22088_ (.A(_18481_),
    .X(_18492_));
 sky130_fd_sc_hd__mux2_2 _22089_ (.A0(\cpuregs[4][7] ),
    .A1(_18491_),
    .S(_18492_),
    .X(_03607_));
 sky130_fd_sc_hd__buf_1 _22090_ (.A(\cpuregs_wrdata[6] ),
    .X(_18493_));
 sky130_fd_sc_hd__mux2_2 _22091_ (.A0(\cpuregs[4][6] ),
    .A1(_18493_),
    .S(_18492_),
    .X(_03606_));
 sky130_fd_sc_hd__buf_1 _22092_ (.A(\cpuregs_wrdata[5] ),
    .X(_18494_));
 sky130_fd_sc_hd__mux2_2 _22093_ (.A0(\cpuregs[4][5] ),
    .A1(_18494_),
    .S(_18492_),
    .X(_03605_));
 sky130_fd_sc_hd__buf_1 _22094_ (.A(\cpuregs_wrdata[4] ),
    .X(_18495_));
 sky130_fd_sc_hd__mux2_2 _22095_ (.A0(\cpuregs[4][4] ),
    .A1(_18495_),
    .S(_18492_),
    .X(_03604_));
 sky130_fd_sc_hd__buf_1 _22096_ (.A(\cpuregs_wrdata[3] ),
    .X(_18496_));
 sky130_fd_sc_hd__buf_1 _22097_ (.A(_18481_),
    .X(_18497_));
 sky130_fd_sc_hd__mux2_2 _22098_ (.A0(\cpuregs[4][3] ),
    .A1(_18496_),
    .S(_18497_),
    .X(_03603_));
 sky130_fd_sc_hd__buf_1 _22099_ (.A(\cpuregs_wrdata[2] ),
    .X(_18498_));
 sky130_fd_sc_hd__mux2_2 _22100_ (.A0(\cpuregs[4][2] ),
    .A1(_18498_),
    .S(_18497_),
    .X(_03602_));
 sky130_fd_sc_hd__buf_1 _22101_ (.A(\cpuregs_wrdata[1] ),
    .X(_18499_));
 sky130_fd_sc_hd__mux2_2 _22102_ (.A0(\cpuregs[4][1] ),
    .A1(_18499_),
    .S(_18497_),
    .X(_03601_));
 sky130_fd_sc_hd__buf_1 _22103_ (.A(\cpuregs_wrdata[0] ),
    .X(_18500_));
 sky130_fd_sc_hd__mux2_2 _22104_ (.A0(\cpuregs[4][0] ),
    .A1(_18500_),
    .S(_18497_),
    .X(_03600_));
 sky130_fd_sc_hd__nor3b_2 _22105_ (.A(_18289_),
    .B(_18288_),
    .C_N(_18287_),
    .Y(_18501_));
 sky130_fd_sc_hd__and2_2 _22106_ (.A(_18283_),
    .B(_18284_),
    .X(_18502_));
 sky130_fd_sc_hd__buf_1 _22107_ (.A(_18502_),
    .X(_18503_));
 sky130_fd_sc_hd__o2111ai_2 _22108_ (.A1(_18276_),
    .A2(_18282_),
    .B1(_18501_),
    .C1(_18503_),
    .D1(_18294_),
    .Y(_18504_));
 sky130_fd_sc_hd__buf_1 _22109_ (.A(_18504_),
    .X(_18505_));
 sky130_fd_sc_hd__buf_1 _22110_ (.A(_18505_),
    .X(_18506_));
 sky130_fd_sc_hd__mux2_2 _22111_ (.A0(_18273_),
    .A1(\cpuregs[19][31] ),
    .S(_18506_),
    .X(_03599_));
 sky130_fd_sc_hd__mux2_2 _22112_ (.A0(_18299_),
    .A1(\cpuregs[19][30] ),
    .S(_18506_),
    .X(_03598_));
 sky130_fd_sc_hd__mux2_2 _22113_ (.A0(_18301_),
    .A1(\cpuregs[19][29] ),
    .S(_18506_),
    .X(_03597_));
 sky130_fd_sc_hd__mux2_2 _22114_ (.A0(_18303_),
    .A1(\cpuregs[19][28] ),
    .S(_18506_),
    .X(_03596_));
 sky130_fd_sc_hd__buf_1 _22115_ (.A(_18505_),
    .X(_18507_));
 sky130_fd_sc_hd__mux2_2 _22116_ (.A0(_18305_),
    .A1(\cpuregs[19][27] ),
    .S(_18507_),
    .X(_03595_));
 sky130_fd_sc_hd__mux2_2 _22117_ (.A0(_18308_),
    .A1(\cpuregs[19][26] ),
    .S(_18507_),
    .X(_03594_));
 sky130_fd_sc_hd__mux2_2 _22118_ (.A0(_18310_),
    .A1(\cpuregs[19][25] ),
    .S(_18507_),
    .X(_03593_));
 sky130_fd_sc_hd__mux2_2 _22119_ (.A0(_18312_),
    .A1(\cpuregs[19][24] ),
    .S(_18507_),
    .X(_03592_));
 sky130_fd_sc_hd__buf_1 _22120_ (.A(_18505_),
    .X(_18508_));
 sky130_fd_sc_hd__mux2_2 _22121_ (.A0(_18314_),
    .A1(\cpuregs[19][23] ),
    .S(_18508_),
    .X(_03591_));
 sky130_fd_sc_hd__mux2_2 _22122_ (.A0(_18317_),
    .A1(\cpuregs[19][22] ),
    .S(_18508_),
    .X(_03590_));
 sky130_fd_sc_hd__mux2_2 _22123_ (.A0(_18319_),
    .A1(\cpuregs[19][21] ),
    .S(_18508_),
    .X(_03589_));
 sky130_fd_sc_hd__mux2_2 _22124_ (.A0(_18321_),
    .A1(\cpuregs[19][20] ),
    .S(_18508_),
    .X(_03588_));
 sky130_fd_sc_hd__buf_1 _22125_ (.A(_18505_),
    .X(_18509_));
 sky130_fd_sc_hd__mux2_2 _22126_ (.A0(_18323_),
    .A1(\cpuregs[19][19] ),
    .S(_18509_),
    .X(_03587_));
 sky130_fd_sc_hd__mux2_2 _22127_ (.A0(_18326_),
    .A1(\cpuregs[19][18] ),
    .S(_18509_),
    .X(_03586_));
 sky130_fd_sc_hd__mux2_2 _22128_ (.A0(_18328_),
    .A1(\cpuregs[19][17] ),
    .S(_18509_),
    .X(_03585_));
 sky130_fd_sc_hd__mux2_2 _22129_ (.A0(_18330_),
    .A1(\cpuregs[19][16] ),
    .S(_18509_),
    .X(_03584_));
 sky130_fd_sc_hd__buf_1 _22130_ (.A(_18504_),
    .X(_18510_));
 sky130_fd_sc_hd__buf_1 _22131_ (.A(_18510_),
    .X(_18511_));
 sky130_fd_sc_hd__mux2_2 _22132_ (.A0(_18332_),
    .A1(\cpuregs[19][15] ),
    .S(_18511_),
    .X(_03583_));
 sky130_fd_sc_hd__mux2_2 _22133_ (.A0(_18336_),
    .A1(\cpuregs[19][14] ),
    .S(_18511_),
    .X(_03582_));
 sky130_fd_sc_hd__mux2_2 _22134_ (.A0(_18338_),
    .A1(\cpuregs[19][13] ),
    .S(_18511_),
    .X(_03581_));
 sky130_fd_sc_hd__mux2_2 _22135_ (.A0(_18340_),
    .A1(\cpuregs[19][12] ),
    .S(_18511_),
    .X(_03580_));
 sky130_fd_sc_hd__buf_1 _22136_ (.A(_18510_),
    .X(_18512_));
 sky130_fd_sc_hd__mux2_2 _22137_ (.A0(_18342_),
    .A1(\cpuregs[19][11] ),
    .S(_18512_),
    .X(_03579_));
 sky130_fd_sc_hd__mux2_2 _22138_ (.A0(_18345_),
    .A1(\cpuregs[19][10] ),
    .S(_18512_),
    .X(_03578_));
 sky130_fd_sc_hd__mux2_2 _22139_ (.A0(_18347_),
    .A1(\cpuregs[19][9] ),
    .S(_18512_),
    .X(_03577_));
 sky130_fd_sc_hd__mux2_2 _22140_ (.A0(_18349_),
    .A1(\cpuregs[19][8] ),
    .S(_18512_),
    .X(_03576_));
 sky130_fd_sc_hd__buf_1 _22141_ (.A(_18510_),
    .X(_18513_));
 sky130_fd_sc_hd__mux2_2 _22142_ (.A0(_18351_),
    .A1(\cpuregs[19][7] ),
    .S(_18513_),
    .X(_03575_));
 sky130_fd_sc_hd__mux2_2 _22143_ (.A0(_18354_),
    .A1(\cpuregs[19][6] ),
    .S(_18513_),
    .X(_03574_));
 sky130_fd_sc_hd__mux2_2 _22144_ (.A0(_18356_),
    .A1(\cpuregs[19][5] ),
    .S(_18513_),
    .X(_03573_));
 sky130_fd_sc_hd__mux2_2 _22145_ (.A0(_18358_),
    .A1(\cpuregs[19][4] ),
    .S(_18513_),
    .X(_03572_));
 sky130_fd_sc_hd__buf_1 _22146_ (.A(_18510_),
    .X(_18514_));
 sky130_fd_sc_hd__mux2_2 _22147_ (.A0(_18360_),
    .A1(\cpuregs[19][3] ),
    .S(_18514_),
    .X(_03571_));
 sky130_fd_sc_hd__mux2_2 _22148_ (.A0(_18363_),
    .A1(\cpuregs[19][2] ),
    .S(_18514_),
    .X(_03570_));
 sky130_fd_sc_hd__mux2_2 _22149_ (.A0(_18365_),
    .A1(\cpuregs[19][1] ),
    .S(_18514_),
    .X(_03569_));
 sky130_fd_sc_hd__mux2_2 _22150_ (.A0(_18367_),
    .A1(\cpuregs[19][0] ),
    .S(_18514_),
    .X(_03568_));
 sky130_fd_sc_hd__nand3_2 _22151_ (.A(_17222_),
    .B(_17217_),
    .C(_17220_),
    .Y(_18515_));
 sky130_fd_sc_hd__buf_1 _22152_ (.A(_18515_),
    .X(_18516_));
 sky130_fd_sc_hd__buf_1 _22153_ (.A(_18516_),
    .X(_18517_));
 sky130_fd_sc_hd__mux2_2 _22154_ (.A0(mem_la_wdata[31]),
    .A1(mem_wdata[31]),
    .S(_18517_),
    .X(_03567_));
 sky130_fd_sc_hd__mux2_2 _22155_ (.A0(mem_la_wdata[30]),
    .A1(mem_wdata[30]),
    .S(_18517_),
    .X(_03566_));
 sky130_fd_sc_hd__mux2_2 _22156_ (.A0(mem_la_wdata[29]),
    .A1(mem_wdata[29]),
    .S(_18517_),
    .X(_03565_));
 sky130_fd_sc_hd__mux2_2 _22157_ (.A0(mem_la_wdata[28]),
    .A1(mem_wdata[28]),
    .S(_18517_),
    .X(_03564_));
 sky130_fd_sc_hd__buf_1 _22158_ (.A(_18516_),
    .X(_18518_));
 sky130_fd_sc_hd__mux2_2 _22159_ (.A0(mem_la_wdata[27]),
    .A1(mem_wdata[27]),
    .S(_18518_),
    .X(_03563_));
 sky130_fd_sc_hd__mux2_2 _22160_ (.A0(mem_la_wdata[26]),
    .A1(mem_wdata[26]),
    .S(_18518_),
    .X(_03562_));
 sky130_fd_sc_hd__mux2_2 _22161_ (.A0(mem_la_wdata[25]),
    .A1(mem_wdata[25]),
    .S(_18518_),
    .X(_03561_));
 sky130_fd_sc_hd__mux2_2 _22162_ (.A0(mem_la_wdata[24]),
    .A1(mem_wdata[24]),
    .S(_18518_),
    .X(_03560_));
 sky130_fd_sc_hd__buf_1 _22163_ (.A(_18516_),
    .X(_18519_));
 sky130_fd_sc_hd__mux2_2 _22164_ (.A0(mem_la_wdata[23]),
    .A1(mem_wdata[23]),
    .S(_18519_),
    .X(_03559_));
 sky130_fd_sc_hd__mux2_2 _22165_ (.A0(mem_la_wdata[22]),
    .A1(mem_wdata[22]),
    .S(_18519_),
    .X(_03558_));
 sky130_fd_sc_hd__mux2_2 _22166_ (.A0(mem_la_wdata[21]),
    .A1(mem_wdata[21]),
    .S(_18519_),
    .X(_03557_));
 sky130_fd_sc_hd__mux2_2 _22167_ (.A0(mem_la_wdata[20]),
    .A1(mem_wdata[20]),
    .S(_18519_),
    .X(_03556_));
 sky130_fd_sc_hd__buf_1 _22168_ (.A(_18516_),
    .X(_18520_));
 sky130_fd_sc_hd__mux2_2 _22169_ (.A0(mem_la_wdata[19]),
    .A1(mem_wdata[19]),
    .S(_18520_),
    .X(_03555_));
 sky130_fd_sc_hd__mux2_2 _22170_ (.A0(mem_la_wdata[18]),
    .A1(mem_wdata[18]),
    .S(_18520_),
    .X(_03554_));
 sky130_fd_sc_hd__mux2_2 _22171_ (.A0(mem_la_wdata[17]),
    .A1(mem_wdata[17]),
    .S(_18520_),
    .X(_03553_));
 sky130_fd_sc_hd__mux2_2 _22172_ (.A0(mem_la_wdata[16]),
    .A1(mem_wdata[16]),
    .S(_18520_),
    .X(_03552_));
 sky130_fd_sc_hd__buf_1 _22173_ (.A(_18515_),
    .X(_18521_));
 sky130_fd_sc_hd__buf_1 _22174_ (.A(_18521_),
    .X(_18522_));
 sky130_fd_sc_hd__mux2_2 _22175_ (.A0(mem_la_wdata[15]),
    .A1(mem_wdata[15]),
    .S(_18522_),
    .X(_03551_));
 sky130_fd_sc_hd__mux2_2 _22176_ (.A0(mem_la_wdata[14]),
    .A1(mem_wdata[14]),
    .S(_18522_),
    .X(_03550_));
 sky130_fd_sc_hd__mux2_2 _22177_ (.A0(mem_la_wdata[13]),
    .A1(mem_wdata[13]),
    .S(_18522_),
    .X(_03549_));
 sky130_fd_sc_hd__mux2_2 _22178_ (.A0(mem_la_wdata[12]),
    .A1(mem_wdata[12]),
    .S(_18522_),
    .X(_03548_));
 sky130_fd_sc_hd__buf_1 _22179_ (.A(_18521_),
    .X(_18523_));
 sky130_fd_sc_hd__mux2_2 _22180_ (.A0(mem_la_wdata[11]),
    .A1(mem_wdata[11]),
    .S(_18523_),
    .X(_03547_));
 sky130_fd_sc_hd__mux2_2 _22181_ (.A0(mem_la_wdata[10]),
    .A1(mem_wdata[10]),
    .S(_18523_),
    .X(_03546_));
 sky130_fd_sc_hd__mux2_2 _22182_ (.A0(mem_la_wdata[9]),
    .A1(mem_wdata[9]),
    .S(_18523_),
    .X(_03545_));
 sky130_fd_sc_hd__mux2_2 _22183_ (.A0(mem_la_wdata[8]),
    .A1(mem_wdata[8]),
    .S(_18523_),
    .X(_03544_));
 sky130_fd_sc_hd__buf_1 _22184_ (.A(_18521_),
    .X(_18524_));
 sky130_fd_sc_hd__mux2_2 _22185_ (.A0(_18434_),
    .A1(mem_wdata[7]),
    .S(_18524_),
    .X(_03543_));
 sky130_fd_sc_hd__mux2_2 _22186_ (.A0(_18437_),
    .A1(mem_wdata[6]),
    .S(_18524_),
    .X(_03542_));
 sky130_fd_sc_hd__mux2_2 _22187_ (.A0(_18440_),
    .A1(mem_wdata[5]),
    .S(_18524_),
    .X(_03541_));
 sky130_fd_sc_hd__mux2_2 _22188_ (.A0(_18442_),
    .A1(mem_wdata[4]),
    .S(_18524_),
    .X(_03540_));
 sky130_fd_sc_hd__buf_1 _22189_ (.A(_18521_),
    .X(_18525_));
 sky130_fd_sc_hd__mux2_2 _22190_ (.A0(_18446_),
    .A1(mem_wdata[3]),
    .S(_18525_),
    .X(_03539_));
 sky130_fd_sc_hd__buf_1 _22191_ (.A(_18448_),
    .X(_18526_));
 sky130_fd_sc_hd__mux2_2 _22192_ (.A0(_18526_),
    .A1(mem_wdata[2]),
    .S(_18525_),
    .X(_03538_));
 sky130_fd_sc_hd__buf_1 _22193_ (.A(_18450_),
    .X(_18527_));
 sky130_fd_sc_hd__mux2_2 _22194_ (.A0(_18527_),
    .A1(mem_wdata[1]),
    .S(_18525_),
    .X(_03537_));
 sky130_fd_sc_hd__mux2_2 _22195_ (.A0(_18455_),
    .A1(mem_wdata[0]),
    .S(_18525_),
    .X(_03536_));
 sky130_fd_sc_hd__buf_1 _22196_ (.A(_18275_),
    .X(_18528_));
 sky130_fd_sc_hd__o2111ai_2 _22197_ (.A1(_18528_),
    .A2(_18282_),
    .B1(_18290_),
    .C1(_18503_),
    .D1(_18294_),
    .Y(_18529_));
 sky130_fd_sc_hd__buf_1 _22198_ (.A(_18529_),
    .X(_18530_));
 sky130_fd_sc_hd__buf_1 _22199_ (.A(_18530_),
    .X(_18531_));
 sky130_fd_sc_hd__mux2_2 _22200_ (.A0(_18273_),
    .A1(\cpuregs[7][31] ),
    .S(_18531_),
    .X(_03535_));
 sky130_fd_sc_hd__mux2_2 _22201_ (.A0(_18299_),
    .A1(\cpuregs[7][30] ),
    .S(_18531_),
    .X(_03534_));
 sky130_fd_sc_hd__mux2_2 _22202_ (.A0(_18301_),
    .A1(\cpuregs[7][29] ),
    .S(_18531_),
    .X(_03533_));
 sky130_fd_sc_hd__mux2_2 _22203_ (.A0(_18303_),
    .A1(\cpuregs[7][28] ),
    .S(_18531_),
    .X(_03532_));
 sky130_fd_sc_hd__buf_1 _22204_ (.A(_18530_),
    .X(_18532_));
 sky130_fd_sc_hd__mux2_2 _22205_ (.A0(_18305_),
    .A1(\cpuregs[7][27] ),
    .S(_18532_),
    .X(_03531_));
 sky130_fd_sc_hd__mux2_2 _22206_ (.A0(_18308_),
    .A1(\cpuregs[7][26] ),
    .S(_18532_),
    .X(_03530_));
 sky130_fd_sc_hd__mux2_2 _22207_ (.A0(_18310_),
    .A1(\cpuregs[7][25] ),
    .S(_18532_),
    .X(_03529_));
 sky130_fd_sc_hd__mux2_2 _22208_ (.A0(_18312_),
    .A1(\cpuregs[7][24] ),
    .S(_18532_),
    .X(_03528_));
 sky130_fd_sc_hd__buf_1 _22209_ (.A(_18530_),
    .X(_18533_));
 sky130_fd_sc_hd__mux2_2 _22210_ (.A0(_18314_),
    .A1(\cpuregs[7][23] ),
    .S(_18533_),
    .X(_03527_));
 sky130_fd_sc_hd__mux2_2 _22211_ (.A0(_18317_),
    .A1(\cpuregs[7][22] ),
    .S(_18533_),
    .X(_03526_));
 sky130_fd_sc_hd__mux2_2 _22212_ (.A0(_18319_),
    .A1(\cpuregs[7][21] ),
    .S(_18533_),
    .X(_03525_));
 sky130_fd_sc_hd__mux2_2 _22213_ (.A0(_18321_),
    .A1(\cpuregs[7][20] ),
    .S(_18533_),
    .X(_03524_));
 sky130_fd_sc_hd__buf_1 _22214_ (.A(_18530_),
    .X(_18534_));
 sky130_fd_sc_hd__mux2_2 _22215_ (.A0(_18323_),
    .A1(\cpuregs[7][19] ),
    .S(_18534_),
    .X(_03523_));
 sky130_fd_sc_hd__mux2_2 _22216_ (.A0(_18326_),
    .A1(\cpuregs[7][18] ),
    .S(_18534_),
    .X(_03522_));
 sky130_fd_sc_hd__mux2_2 _22217_ (.A0(_18328_),
    .A1(\cpuregs[7][17] ),
    .S(_18534_),
    .X(_03521_));
 sky130_fd_sc_hd__mux2_2 _22218_ (.A0(_18330_),
    .A1(\cpuregs[7][16] ),
    .S(_18534_),
    .X(_03520_));
 sky130_fd_sc_hd__buf_1 _22219_ (.A(_18529_),
    .X(_18535_));
 sky130_fd_sc_hd__buf_1 _22220_ (.A(_18535_),
    .X(_18536_));
 sky130_fd_sc_hd__mux2_2 _22221_ (.A0(_18332_),
    .A1(\cpuregs[7][15] ),
    .S(_18536_),
    .X(_03519_));
 sky130_fd_sc_hd__mux2_2 _22222_ (.A0(_18336_),
    .A1(\cpuregs[7][14] ),
    .S(_18536_),
    .X(_03518_));
 sky130_fd_sc_hd__mux2_2 _22223_ (.A0(_18338_),
    .A1(\cpuregs[7][13] ),
    .S(_18536_),
    .X(_03517_));
 sky130_fd_sc_hd__mux2_2 _22224_ (.A0(_18340_),
    .A1(\cpuregs[7][12] ),
    .S(_18536_),
    .X(_03516_));
 sky130_fd_sc_hd__buf_1 _22225_ (.A(_18535_),
    .X(_18537_));
 sky130_fd_sc_hd__mux2_2 _22226_ (.A0(_18342_),
    .A1(\cpuregs[7][11] ),
    .S(_18537_),
    .X(_03515_));
 sky130_fd_sc_hd__mux2_2 _22227_ (.A0(_18345_),
    .A1(\cpuregs[7][10] ),
    .S(_18537_),
    .X(_03514_));
 sky130_fd_sc_hd__mux2_2 _22228_ (.A0(_18347_),
    .A1(\cpuregs[7][9] ),
    .S(_18537_),
    .X(_03513_));
 sky130_fd_sc_hd__mux2_2 _22229_ (.A0(_18349_),
    .A1(\cpuregs[7][8] ),
    .S(_18537_),
    .X(_03512_));
 sky130_fd_sc_hd__buf_1 _22230_ (.A(_18535_),
    .X(_18538_));
 sky130_fd_sc_hd__mux2_2 _22231_ (.A0(_18351_),
    .A1(\cpuregs[7][7] ),
    .S(_18538_),
    .X(_03511_));
 sky130_fd_sc_hd__mux2_2 _22232_ (.A0(_18354_),
    .A1(\cpuregs[7][6] ),
    .S(_18538_),
    .X(_03510_));
 sky130_fd_sc_hd__mux2_2 _22233_ (.A0(_18356_),
    .A1(\cpuregs[7][5] ),
    .S(_18538_),
    .X(_03509_));
 sky130_fd_sc_hd__mux2_2 _22234_ (.A0(_18358_),
    .A1(\cpuregs[7][4] ),
    .S(_18538_),
    .X(_03508_));
 sky130_fd_sc_hd__buf_1 _22235_ (.A(_18535_),
    .X(_18539_));
 sky130_fd_sc_hd__mux2_2 _22236_ (.A0(_18360_),
    .A1(\cpuregs[7][3] ),
    .S(_18539_),
    .X(_03507_));
 sky130_fd_sc_hd__mux2_2 _22237_ (.A0(_18363_),
    .A1(\cpuregs[7][2] ),
    .S(_18539_),
    .X(_03506_));
 sky130_fd_sc_hd__mux2_2 _22238_ (.A0(_18365_),
    .A1(\cpuregs[7][1] ),
    .S(_18539_),
    .X(_03505_));
 sky130_fd_sc_hd__mux2_2 _22239_ (.A0(_18367_),
    .A1(\cpuregs[7][0] ),
    .S(_18539_),
    .X(_03504_));
 sky130_fd_sc_hd__buf_1 _22240_ (.A(_17020_),
    .X(_18540_));
 sky130_fd_sc_hd__buf_1 _22241_ (.A(_18540_),
    .X(_18541_));
 sky130_vsdinv _22242_ (.A(is_beq_bne_blt_bge_bltu_bgeu),
    .Y(_18542_));
 sky130_fd_sc_hd__nand3_2 _22243_ (.A(_18542_),
    .B(_00302_),
    .C(\cpu_state[4] ),
    .Y(_18543_));
 sky130_fd_sc_hd__nor3b_2 _22244_ (.A(_16841_),
    .B(_00331_),
    .C_N(_18543_),
    .Y(_18544_));
 sky130_fd_sc_hd__o21ai_2 _22245_ (.A1(instr_setq),
    .A2(_18541_),
    .B1(_18544_),
    .Y(_18545_));
 sky130_fd_sc_hd__mux2_2 _22246_ (.A0(_19779_),
    .A1(_18287_),
    .S(_18545_),
    .X(_03503_));
 sky130_fd_sc_hd__buf_1 _22247_ (.A(\cpuregs_wrdata[31] ),
    .X(_18546_));
 sky130_fd_sc_hd__buf_1 _22248_ (.A(_18280_),
    .X(_18547_));
 sky130_fd_sc_hd__nand3b_2 _22249_ (.A_N(\latched_rd[4] ),
    .B(_18289_),
    .C(_18288_),
    .Y(_18548_));
 sky130_vsdinv _22250_ (.A(_18548_),
    .Y(_18549_));
 sky130_fd_sc_hd__buf_1 _22251_ (.A(_18293_),
    .X(_18550_));
 sky130_fd_sc_hd__o2111ai_2 _22252_ (.A1(_18528_),
    .A2(_18547_),
    .B1(_18503_),
    .C1(_18549_),
    .D1(_18550_),
    .Y(_18551_));
 sky130_fd_sc_hd__buf_1 _22253_ (.A(_18551_),
    .X(_18552_));
 sky130_fd_sc_hd__buf_1 _22254_ (.A(_18552_),
    .X(_18553_));
 sky130_fd_sc_hd__mux2_2 _22255_ (.A0(_18546_),
    .A1(\cpuregs[15][31] ),
    .S(_18553_),
    .X(_03502_));
 sky130_fd_sc_hd__buf_1 _22256_ (.A(\cpuregs_wrdata[30] ),
    .X(_18554_));
 sky130_fd_sc_hd__mux2_2 _22257_ (.A0(_18554_),
    .A1(\cpuregs[15][30] ),
    .S(_18553_),
    .X(_03501_));
 sky130_fd_sc_hd__buf_1 _22258_ (.A(\cpuregs_wrdata[29] ),
    .X(_18555_));
 sky130_fd_sc_hd__mux2_2 _22259_ (.A0(_18555_),
    .A1(\cpuregs[15][29] ),
    .S(_18553_),
    .X(_03500_));
 sky130_fd_sc_hd__buf_1 _22260_ (.A(\cpuregs_wrdata[28] ),
    .X(_18556_));
 sky130_fd_sc_hd__mux2_2 _22261_ (.A0(_18556_),
    .A1(\cpuregs[15][28] ),
    .S(_18553_),
    .X(_03499_));
 sky130_fd_sc_hd__buf_1 _22262_ (.A(\cpuregs_wrdata[27] ),
    .X(_18557_));
 sky130_fd_sc_hd__buf_1 _22263_ (.A(_18552_),
    .X(_18558_));
 sky130_fd_sc_hd__mux2_2 _22264_ (.A0(_18557_),
    .A1(\cpuregs[15][27] ),
    .S(_18558_),
    .X(_03498_));
 sky130_fd_sc_hd__buf_1 _22265_ (.A(\cpuregs_wrdata[26] ),
    .X(_18559_));
 sky130_fd_sc_hd__mux2_2 _22266_ (.A0(_18559_),
    .A1(\cpuregs[15][26] ),
    .S(_18558_),
    .X(_03497_));
 sky130_fd_sc_hd__buf_1 _22267_ (.A(\cpuregs_wrdata[25] ),
    .X(_18560_));
 sky130_fd_sc_hd__mux2_2 _22268_ (.A0(_18560_),
    .A1(\cpuregs[15][25] ),
    .S(_18558_),
    .X(_03496_));
 sky130_fd_sc_hd__buf_1 _22269_ (.A(\cpuregs_wrdata[24] ),
    .X(_18561_));
 sky130_fd_sc_hd__mux2_2 _22270_ (.A0(_18561_),
    .A1(\cpuregs[15][24] ),
    .S(_18558_),
    .X(_03495_));
 sky130_fd_sc_hd__buf_1 _22271_ (.A(\cpuregs_wrdata[23] ),
    .X(_18562_));
 sky130_fd_sc_hd__buf_1 _22272_ (.A(_18552_),
    .X(_18563_));
 sky130_fd_sc_hd__mux2_2 _22273_ (.A0(_18562_),
    .A1(\cpuregs[15][23] ),
    .S(_18563_),
    .X(_03494_));
 sky130_fd_sc_hd__buf_1 _22274_ (.A(\cpuregs_wrdata[22] ),
    .X(_18564_));
 sky130_fd_sc_hd__mux2_2 _22275_ (.A0(_18564_),
    .A1(\cpuregs[15][22] ),
    .S(_18563_),
    .X(_03493_));
 sky130_fd_sc_hd__buf_1 _22276_ (.A(\cpuregs_wrdata[21] ),
    .X(_18565_));
 sky130_fd_sc_hd__mux2_2 _22277_ (.A0(_18565_),
    .A1(\cpuregs[15][21] ),
    .S(_18563_),
    .X(_03492_));
 sky130_fd_sc_hd__buf_1 _22278_ (.A(\cpuregs_wrdata[20] ),
    .X(_18566_));
 sky130_fd_sc_hd__mux2_2 _22279_ (.A0(_18566_),
    .A1(\cpuregs[15][20] ),
    .S(_18563_),
    .X(_03491_));
 sky130_fd_sc_hd__buf_1 _22280_ (.A(\cpuregs_wrdata[19] ),
    .X(_18567_));
 sky130_fd_sc_hd__buf_1 _22281_ (.A(_18552_),
    .X(_18568_));
 sky130_fd_sc_hd__mux2_2 _22282_ (.A0(_18567_),
    .A1(\cpuregs[15][19] ),
    .S(_18568_),
    .X(_03490_));
 sky130_fd_sc_hd__buf_1 _22283_ (.A(\cpuregs_wrdata[18] ),
    .X(_18569_));
 sky130_fd_sc_hd__mux2_2 _22284_ (.A0(_18569_),
    .A1(\cpuregs[15][18] ),
    .S(_18568_),
    .X(_03489_));
 sky130_fd_sc_hd__buf_1 _22285_ (.A(\cpuregs_wrdata[17] ),
    .X(_18570_));
 sky130_fd_sc_hd__mux2_2 _22286_ (.A0(_18570_),
    .A1(\cpuregs[15][17] ),
    .S(_18568_),
    .X(_03488_));
 sky130_fd_sc_hd__buf_1 _22287_ (.A(\cpuregs_wrdata[16] ),
    .X(_18571_));
 sky130_fd_sc_hd__mux2_2 _22288_ (.A0(_18571_),
    .A1(\cpuregs[15][16] ),
    .S(_18568_),
    .X(_03487_));
 sky130_fd_sc_hd__buf_1 _22289_ (.A(\cpuregs_wrdata[15] ),
    .X(_18572_));
 sky130_fd_sc_hd__buf_1 _22290_ (.A(_18551_),
    .X(_18573_));
 sky130_fd_sc_hd__buf_1 _22291_ (.A(_18573_),
    .X(_18574_));
 sky130_fd_sc_hd__mux2_2 _22292_ (.A0(_18572_),
    .A1(\cpuregs[15][15] ),
    .S(_18574_),
    .X(_03486_));
 sky130_fd_sc_hd__buf_1 _22293_ (.A(\cpuregs_wrdata[14] ),
    .X(_18575_));
 sky130_fd_sc_hd__mux2_2 _22294_ (.A0(_18575_),
    .A1(\cpuregs[15][14] ),
    .S(_18574_),
    .X(_03485_));
 sky130_fd_sc_hd__buf_1 _22295_ (.A(\cpuregs_wrdata[13] ),
    .X(_18576_));
 sky130_fd_sc_hd__mux2_2 _22296_ (.A0(_18576_),
    .A1(\cpuregs[15][13] ),
    .S(_18574_),
    .X(_03484_));
 sky130_fd_sc_hd__buf_1 _22297_ (.A(\cpuregs_wrdata[12] ),
    .X(_18577_));
 sky130_fd_sc_hd__mux2_2 _22298_ (.A0(_18577_),
    .A1(\cpuregs[15][12] ),
    .S(_18574_),
    .X(_03483_));
 sky130_fd_sc_hd__buf_1 _22299_ (.A(\cpuregs_wrdata[11] ),
    .X(_18578_));
 sky130_fd_sc_hd__buf_1 _22300_ (.A(_18573_),
    .X(_18579_));
 sky130_fd_sc_hd__mux2_2 _22301_ (.A0(_18578_),
    .A1(\cpuregs[15][11] ),
    .S(_18579_),
    .X(_03482_));
 sky130_fd_sc_hd__buf_1 _22302_ (.A(\cpuregs_wrdata[10] ),
    .X(_18580_));
 sky130_fd_sc_hd__mux2_2 _22303_ (.A0(_18580_),
    .A1(\cpuregs[15][10] ),
    .S(_18579_),
    .X(_03481_));
 sky130_fd_sc_hd__buf_1 _22304_ (.A(\cpuregs_wrdata[9] ),
    .X(_18581_));
 sky130_fd_sc_hd__mux2_2 _22305_ (.A0(_18581_),
    .A1(\cpuregs[15][9] ),
    .S(_18579_),
    .X(_03480_));
 sky130_fd_sc_hd__buf_1 _22306_ (.A(\cpuregs_wrdata[8] ),
    .X(_18582_));
 sky130_fd_sc_hd__mux2_2 _22307_ (.A0(_18582_),
    .A1(\cpuregs[15][8] ),
    .S(_18579_),
    .X(_03479_));
 sky130_fd_sc_hd__buf_1 _22308_ (.A(\cpuregs_wrdata[7] ),
    .X(_18583_));
 sky130_fd_sc_hd__buf_1 _22309_ (.A(_18573_),
    .X(_18584_));
 sky130_fd_sc_hd__mux2_2 _22310_ (.A0(_18583_),
    .A1(\cpuregs[15][7] ),
    .S(_18584_),
    .X(_03478_));
 sky130_fd_sc_hd__buf_1 _22311_ (.A(\cpuregs_wrdata[6] ),
    .X(_18585_));
 sky130_fd_sc_hd__mux2_2 _22312_ (.A0(_18585_),
    .A1(\cpuregs[15][6] ),
    .S(_18584_),
    .X(_03477_));
 sky130_fd_sc_hd__buf_1 _22313_ (.A(\cpuregs_wrdata[5] ),
    .X(_18586_));
 sky130_fd_sc_hd__mux2_2 _22314_ (.A0(_18586_),
    .A1(\cpuregs[15][5] ),
    .S(_18584_),
    .X(_03476_));
 sky130_fd_sc_hd__buf_1 _22315_ (.A(\cpuregs_wrdata[4] ),
    .X(_18587_));
 sky130_fd_sc_hd__mux2_2 _22316_ (.A0(_18587_),
    .A1(\cpuregs[15][4] ),
    .S(_18584_),
    .X(_03475_));
 sky130_fd_sc_hd__buf_1 _22317_ (.A(\cpuregs_wrdata[3] ),
    .X(_18588_));
 sky130_fd_sc_hd__buf_1 _22318_ (.A(_18573_),
    .X(_18589_));
 sky130_fd_sc_hd__mux2_2 _22319_ (.A0(_18588_),
    .A1(\cpuregs[15][3] ),
    .S(_18589_),
    .X(_03474_));
 sky130_fd_sc_hd__buf_1 _22320_ (.A(\cpuregs_wrdata[2] ),
    .X(_18590_));
 sky130_fd_sc_hd__mux2_2 _22321_ (.A0(_18590_),
    .A1(\cpuregs[15][2] ),
    .S(_18589_),
    .X(_03473_));
 sky130_fd_sc_hd__buf_1 _22322_ (.A(\cpuregs_wrdata[1] ),
    .X(_18591_));
 sky130_fd_sc_hd__mux2_2 _22323_ (.A0(_18591_),
    .A1(\cpuregs[15][1] ),
    .S(_18589_),
    .X(_03472_));
 sky130_fd_sc_hd__buf_1 _22324_ (.A(\cpuregs_wrdata[0] ),
    .X(_18592_));
 sky130_fd_sc_hd__mux2_2 _22325_ (.A0(_18592_),
    .A1(\cpuregs[15][0] ),
    .S(_18589_),
    .X(_03471_));
 sky130_fd_sc_hd__o2111ai_2 _22326_ (.A1(_18528_),
    .A2(_18547_),
    .B1(_18368_),
    .C1(_18503_),
    .D1(_18550_),
    .Y(_18593_));
 sky130_fd_sc_hd__buf_1 _22327_ (.A(_18593_),
    .X(_18594_));
 sky130_fd_sc_hd__buf_1 _22328_ (.A(_18594_),
    .X(_18595_));
 sky130_fd_sc_hd__mux2_2 _22329_ (.A0(_18546_),
    .A1(\cpuregs[11][31] ),
    .S(_18595_),
    .X(_03470_));
 sky130_fd_sc_hd__mux2_2 _22330_ (.A0(_18554_),
    .A1(\cpuregs[11][30] ),
    .S(_18595_),
    .X(_03469_));
 sky130_fd_sc_hd__mux2_2 _22331_ (.A0(_18555_),
    .A1(\cpuregs[11][29] ),
    .S(_18595_),
    .X(_03468_));
 sky130_fd_sc_hd__mux2_2 _22332_ (.A0(_18556_),
    .A1(\cpuregs[11][28] ),
    .S(_18595_),
    .X(_03467_));
 sky130_fd_sc_hd__buf_1 _22333_ (.A(_18594_),
    .X(_18596_));
 sky130_fd_sc_hd__mux2_2 _22334_ (.A0(_18557_),
    .A1(\cpuregs[11][27] ),
    .S(_18596_),
    .X(_03466_));
 sky130_fd_sc_hd__mux2_2 _22335_ (.A0(_18559_),
    .A1(\cpuregs[11][26] ),
    .S(_18596_),
    .X(_03465_));
 sky130_fd_sc_hd__mux2_2 _22336_ (.A0(_18560_),
    .A1(\cpuregs[11][25] ),
    .S(_18596_),
    .X(_03464_));
 sky130_fd_sc_hd__mux2_2 _22337_ (.A0(_18561_),
    .A1(\cpuregs[11][24] ),
    .S(_18596_),
    .X(_03463_));
 sky130_fd_sc_hd__buf_1 _22338_ (.A(_18594_),
    .X(_18597_));
 sky130_fd_sc_hd__mux2_2 _22339_ (.A0(_18562_),
    .A1(\cpuregs[11][23] ),
    .S(_18597_),
    .X(_03462_));
 sky130_fd_sc_hd__mux2_2 _22340_ (.A0(_18564_),
    .A1(\cpuregs[11][22] ),
    .S(_18597_),
    .X(_03461_));
 sky130_fd_sc_hd__mux2_2 _22341_ (.A0(_18565_),
    .A1(\cpuregs[11][21] ),
    .S(_18597_),
    .X(_03460_));
 sky130_fd_sc_hd__mux2_2 _22342_ (.A0(_18566_),
    .A1(\cpuregs[11][20] ),
    .S(_18597_),
    .X(_03459_));
 sky130_fd_sc_hd__buf_1 _22343_ (.A(_18594_),
    .X(_18598_));
 sky130_fd_sc_hd__mux2_2 _22344_ (.A0(_18567_),
    .A1(\cpuregs[11][19] ),
    .S(_18598_),
    .X(_03458_));
 sky130_fd_sc_hd__mux2_2 _22345_ (.A0(_18569_),
    .A1(\cpuregs[11][18] ),
    .S(_18598_),
    .X(_03457_));
 sky130_fd_sc_hd__mux2_2 _22346_ (.A0(_18570_),
    .A1(\cpuregs[11][17] ),
    .S(_18598_),
    .X(_03456_));
 sky130_fd_sc_hd__mux2_2 _22347_ (.A0(_18571_),
    .A1(\cpuregs[11][16] ),
    .S(_18598_),
    .X(_03455_));
 sky130_fd_sc_hd__buf_1 _22348_ (.A(_18593_),
    .X(_18599_));
 sky130_fd_sc_hd__buf_1 _22349_ (.A(_18599_),
    .X(_18600_));
 sky130_fd_sc_hd__mux2_2 _22350_ (.A0(_18572_),
    .A1(\cpuregs[11][15] ),
    .S(_18600_),
    .X(_03454_));
 sky130_fd_sc_hd__mux2_2 _22351_ (.A0(_18575_),
    .A1(\cpuregs[11][14] ),
    .S(_18600_),
    .X(_03453_));
 sky130_fd_sc_hd__mux2_2 _22352_ (.A0(_18576_),
    .A1(\cpuregs[11][13] ),
    .S(_18600_),
    .X(_03452_));
 sky130_fd_sc_hd__mux2_2 _22353_ (.A0(_18577_),
    .A1(\cpuregs[11][12] ),
    .S(_18600_),
    .X(_03451_));
 sky130_fd_sc_hd__buf_1 _22354_ (.A(_18599_),
    .X(_18601_));
 sky130_fd_sc_hd__mux2_2 _22355_ (.A0(_18578_),
    .A1(\cpuregs[11][11] ),
    .S(_18601_),
    .X(_03450_));
 sky130_fd_sc_hd__mux2_2 _22356_ (.A0(_18580_),
    .A1(\cpuregs[11][10] ),
    .S(_18601_),
    .X(_03449_));
 sky130_fd_sc_hd__mux2_2 _22357_ (.A0(_18581_),
    .A1(\cpuregs[11][9] ),
    .S(_18601_),
    .X(_03448_));
 sky130_fd_sc_hd__mux2_2 _22358_ (.A0(_18582_),
    .A1(\cpuregs[11][8] ),
    .S(_18601_),
    .X(_03447_));
 sky130_fd_sc_hd__buf_1 _22359_ (.A(_18599_),
    .X(_18602_));
 sky130_fd_sc_hd__mux2_2 _22360_ (.A0(_18583_),
    .A1(\cpuregs[11][7] ),
    .S(_18602_),
    .X(_03446_));
 sky130_fd_sc_hd__mux2_2 _22361_ (.A0(_18585_),
    .A1(\cpuregs[11][6] ),
    .S(_18602_),
    .X(_03445_));
 sky130_fd_sc_hd__mux2_2 _22362_ (.A0(_18586_),
    .A1(\cpuregs[11][5] ),
    .S(_18602_),
    .X(_03444_));
 sky130_fd_sc_hd__mux2_2 _22363_ (.A0(_18587_),
    .A1(\cpuregs[11][4] ),
    .S(_18602_),
    .X(_03443_));
 sky130_fd_sc_hd__buf_1 _22364_ (.A(_18599_),
    .X(_18603_));
 sky130_fd_sc_hd__mux2_2 _22365_ (.A0(_18588_),
    .A1(\cpuregs[11][3] ),
    .S(_18603_),
    .X(_03442_));
 sky130_fd_sc_hd__mux2_2 _22366_ (.A0(_18590_),
    .A1(\cpuregs[11][2] ),
    .S(_18603_),
    .X(_03441_));
 sky130_fd_sc_hd__mux2_2 _22367_ (.A0(_18591_),
    .A1(\cpuregs[11][1] ),
    .S(_18603_),
    .X(_03440_));
 sky130_fd_sc_hd__mux2_2 _22368_ (.A0(_18592_),
    .A1(\cpuregs[11][0] ),
    .S(_18603_),
    .X(_03439_));
 sky130_fd_sc_hd__and3b_2 _22369_ (.A_N(_18281_),
    .B(_18458_),
    .C(_18502_),
    .X(_18604_));
 sky130_fd_sc_hd__buf_1 _22370_ (.A(_18604_),
    .X(_18605_));
 sky130_fd_sc_hd__buf_1 _22371_ (.A(_18605_),
    .X(_18606_));
 sky130_fd_sc_hd__mux2_2 _22372_ (.A0(\cpuregs[3][31] ),
    .A1(_18272_),
    .S(_18606_),
    .X(_03438_));
 sky130_fd_sc_hd__mux2_2 _22373_ (.A0(\cpuregs[3][30] ),
    .A1(_18298_),
    .S(_18606_),
    .X(_03437_));
 sky130_fd_sc_hd__mux2_2 _22374_ (.A0(\cpuregs[3][29] ),
    .A1(_18300_),
    .S(_18606_),
    .X(_03436_));
 sky130_fd_sc_hd__mux2_2 _22375_ (.A0(\cpuregs[3][28] ),
    .A1(_18302_),
    .S(_18606_),
    .X(_03435_));
 sky130_fd_sc_hd__buf_1 _22376_ (.A(_18605_),
    .X(_18607_));
 sky130_fd_sc_hd__mux2_2 _22377_ (.A0(\cpuregs[3][27] ),
    .A1(_18304_),
    .S(_18607_),
    .X(_03434_));
 sky130_fd_sc_hd__mux2_2 _22378_ (.A0(\cpuregs[3][26] ),
    .A1(_18307_),
    .S(_18607_),
    .X(_03433_));
 sky130_fd_sc_hd__mux2_2 _22379_ (.A0(\cpuregs[3][25] ),
    .A1(_18309_),
    .S(_18607_),
    .X(_03432_));
 sky130_fd_sc_hd__mux2_2 _22380_ (.A0(\cpuregs[3][24] ),
    .A1(_18311_),
    .S(_18607_),
    .X(_03431_));
 sky130_fd_sc_hd__buf_1 _22381_ (.A(_18605_),
    .X(_18608_));
 sky130_fd_sc_hd__mux2_2 _22382_ (.A0(\cpuregs[3][23] ),
    .A1(_18313_),
    .S(_18608_),
    .X(_03430_));
 sky130_fd_sc_hd__mux2_2 _22383_ (.A0(\cpuregs[3][22] ),
    .A1(_18316_),
    .S(_18608_),
    .X(_03429_));
 sky130_fd_sc_hd__mux2_2 _22384_ (.A0(\cpuregs[3][21] ),
    .A1(_18318_),
    .S(_18608_),
    .X(_03428_));
 sky130_fd_sc_hd__mux2_2 _22385_ (.A0(\cpuregs[3][20] ),
    .A1(_18320_),
    .S(_18608_),
    .X(_03427_));
 sky130_fd_sc_hd__buf_1 _22386_ (.A(_18605_),
    .X(_18609_));
 sky130_fd_sc_hd__mux2_2 _22387_ (.A0(\cpuregs[3][19] ),
    .A1(_18322_),
    .S(_18609_),
    .X(_03426_));
 sky130_fd_sc_hd__mux2_2 _22388_ (.A0(\cpuregs[3][18] ),
    .A1(_18325_),
    .S(_18609_),
    .X(_03425_));
 sky130_fd_sc_hd__mux2_2 _22389_ (.A0(\cpuregs[3][17] ),
    .A1(_18327_),
    .S(_18609_),
    .X(_03424_));
 sky130_fd_sc_hd__mux2_2 _22390_ (.A0(\cpuregs[3][16] ),
    .A1(_18329_),
    .S(_18609_),
    .X(_03423_));
 sky130_fd_sc_hd__buf_1 _22391_ (.A(_18604_),
    .X(_18610_));
 sky130_fd_sc_hd__buf_1 _22392_ (.A(_18610_),
    .X(_18611_));
 sky130_fd_sc_hd__mux2_2 _22393_ (.A0(\cpuregs[3][15] ),
    .A1(_18331_),
    .S(_18611_),
    .X(_03422_));
 sky130_fd_sc_hd__mux2_2 _22394_ (.A0(\cpuregs[3][14] ),
    .A1(_18335_),
    .S(_18611_),
    .X(_03421_));
 sky130_fd_sc_hd__mux2_2 _22395_ (.A0(\cpuregs[3][13] ),
    .A1(_18337_),
    .S(_18611_),
    .X(_03420_));
 sky130_fd_sc_hd__mux2_2 _22396_ (.A0(\cpuregs[3][12] ),
    .A1(_18339_),
    .S(_18611_),
    .X(_03419_));
 sky130_fd_sc_hd__buf_1 _22397_ (.A(_18610_),
    .X(_18612_));
 sky130_fd_sc_hd__mux2_2 _22398_ (.A0(\cpuregs[3][11] ),
    .A1(_18341_),
    .S(_18612_),
    .X(_03418_));
 sky130_fd_sc_hd__mux2_2 _22399_ (.A0(\cpuregs[3][10] ),
    .A1(_18344_),
    .S(_18612_),
    .X(_03417_));
 sky130_fd_sc_hd__mux2_2 _22400_ (.A0(\cpuregs[3][9] ),
    .A1(_18346_),
    .S(_18612_),
    .X(_03416_));
 sky130_fd_sc_hd__mux2_2 _22401_ (.A0(\cpuregs[3][8] ),
    .A1(_18348_),
    .S(_18612_),
    .X(_03415_));
 sky130_fd_sc_hd__buf_1 _22402_ (.A(_18610_),
    .X(_18613_));
 sky130_fd_sc_hd__mux2_2 _22403_ (.A0(\cpuregs[3][7] ),
    .A1(_18350_),
    .S(_18613_),
    .X(_03414_));
 sky130_fd_sc_hd__mux2_2 _22404_ (.A0(\cpuregs[3][6] ),
    .A1(_18353_),
    .S(_18613_),
    .X(_03413_));
 sky130_fd_sc_hd__mux2_2 _22405_ (.A0(\cpuregs[3][5] ),
    .A1(_18355_),
    .S(_18613_),
    .X(_03412_));
 sky130_fd_sc_hd__mux2_2 _22406_ (.A0(\cpuregs[3][4] ),
    .A1(_18357_),
    .S(_18613_),
    .X(_03411_));
 sky130_fd_sc_hd__buf_1 _22407_ (.A(_18610_),
    .X(_18614_));
 sky130_fd_sc_hd__mux2_2 _22408_ (.A0(\cpuregs[3][3] ),
    .A1(_18359_),
    .S(_18614_),
    .X(_03410_));
 sky130_fd_sc_hd__mux2_2 _22409_ (.A0(\cpuregs[3][2] ),
    .A1(_18362_),
    .S(_18614_),
    .X(_03409_));
 sky130_fd_sc_hd__mux2_2 _22410_ (.A0(\cpuregs[3][1] ),
    .A1(_18364_),
    .S(_18614_),
    .X(_03408_));
 sky130_fd_sc_hd__mux2_2 _22411_ (.A0(\cpuregs[3][0] ),
    .A1(_18366_),
    .S(_18614_),
    .X(_03407_));
 sky130_fd_sc_hd__and3b_2 _22412_ (.A_N(_18281_),
    .B(_18457_),
    .C(_18369_),
    .X(_18615_));
 sky130_fd_sc_hd__buf_1 _22413_ (.A(_18615_),
    .X(_18616_));
 sky130_fd_sc_hd__buf_1 _22414_ (.A(_18616_),
    .X(_18617_));
 sky130_fd_sc_hd__mux2_2 _22415_ (.A0(\cpuregs[1][31] ),
    .A1(_18272_),
    .S(_18617_),
    .X(_03406_));
 sky130_fd_sc_hd__mux2_2 _22416_ (.A0(\cpuregs[1][30] ),
    .A1(_18298_),
    .S(_18617_),
    .X(_03405_));
 sky130_fd_sc_hd__mux2_2 _22417_ (.A0(\cpuregs[1][29] ),
    .A1(_18300_),
    .S(_18617_),
    .X(_03404_));
 sky130_fd_sc_hd__mux2_2 _22418_ (.A0(\cpuregs[1][28] ),
    .A1(_18302_),
    .S(_18617_),
    .X(_03403_));
 sky130_fd_sc_hd__buf_1 _22419_ (.A(_18616_),
    .X(_18618_));
 sky130_fd_sc_hd__mux2_2 _22420_ (.A0(\cpuregs[1][27] ),
    .A1(_18304_),
    .S(_18618_),
    .X(_03402_));
 sky130_fd_sc_hd__mux2_2 _22421_ (.A0(\cpuregs[1][26] ),
    .A1(_18307_),
    .S(_18618_),
    .X(_03401_));
 sky130_fd_sc_hd__mux2_2 _22422_ (.A0(\cpuregs[1][25] ),
    .A1(_18309_),
    .S(_18618_),
    .X(_03400_));
 sky130_fd_sc_hd__mux2_2 _22423_ (.A0(\cpuregs[1][24] ),
    .A1(_18311_),
    .S(_18618_),
    .X(_03399_));
 sky130_fd_sc_hd__buf_1 _22424_ (.A(_18616_),
    .X(_18619_));
 sky130_fd_sc_hd__mux2_2 _22425_ (.A0(\cpuregs[1][23] ),
    .A1(_18313_),
    .S(_18619_),
    .X(_03398_));
 sky130_fd_sc_hd__mux2_2 _22426_ (.A0(\cpuregs[1][22] ),
    .A1(_18316_),
    .S(_18619_),
    .X(_03397_));
 sky130_fd_sc_hd__mux2_2 _22427_ (.A0(\cpuregs[1][21] ),
    .A1(_18318_),
    .S(_18619_),
    .X(_03396_));
 sky130_fd_sc_hd__mux2_2 _22428_ (.A0(\cpuregs[1][20] ),
    .A1(_18320_),
    .S(_18619_),
    .X(_03395_));
 sky130_fd_sc_hd__buf_1 _22429_ (.A(_18616_),
    .X(_18620_));
 sky130_fd_sc_hd__mux2_2 _22430_ (.A0(\cpuregs[1][19] ),
    .A1(_18322_),
    .S(_18620_),
    .X(_03394_));
 sky130_fd_sc_hd__mux2_2 _22431_ (.A0(\cpuregs[1][18] ),
    .A1(_18325_),
    .S(_18620_),
    .X(_03393_));
 sky130_fd_sc_hd__mux2_2 _22432_ (.A0(\cpuregs[1][17] ),
    .A1(_18327_),
    .S(_18620_),
    .X(_03392_));
 sky130_fd_sc_hd__mux2_2 _22433_ (.A0(\cpuregs[1][16] ),
    .A1(_18329_),
    .S(_18620_),
    .X(_03391_));
 sky130_fd_sc_hd__buf_1 _22434_ (.A(_18615_),
    .X(_18621_));
 sky130_fd_sc_hd__buf_1 _22435_ (.A(_18621_),
    .X(_18622_));
 sky130_fd_sc_hd__mux2_2 _22436_ (.A0(\cpuregs[1][15] ),
    .A1(_18331_),
    .S(_18622_),
    .X(_03390_));
 sky130_fd_sc_hd__mux2_2 _22437_ (.A0(\cpuregs[1][14] ),
    .A1(_18335_),
    .S(_18622_),
    .X(_03389_));
 sky130_fd_sc_hd__mux2_2 _22438_ (.A0(\cpuregs[1][13] ),
    .A1(_18337_),
    .S(_18622_),
    .X(_03388_));
 sky130_fd_sc_hd__mux2_2 _22439_ (.A0(\cpuregs[1][12] ),
    .A1(_18339_),
    .S(_18622_),
    .X(_03387_));
 sky130_fd_sc_hd__buf_1 _22440_ (.A(_18621_),
    .X(_18623_));
 sky130_fd_sc_hd__mux2_2 _22441_ (.A0(\cpuregs[1][11] ),
    .A1(_18341_),
    .S(_18623_),
    .X(_03386_));
 sky130_fd_sc_hd__mux2_2 _22442_ (.A0(\cpuregs[1][10] ),
    .A1(_18344_),
    .S(_18623_),
    .X(_03385_));
 sky130_fd_sc_hd__mux2_2 _22443_ (.A0(\cpuregs[1][9] ),
    .A1(_18346_),
    .S(_18623_),
    .X(_03384_));
 sky130_fd_sc_hd__mux2_2 _22444_ (.A0(\cpuregs[1][8] ),
    .A1(_18348_),
    .S(_18623_),
    .X(_03383_));
 sky130_fd_sc_hd__buf_1 _22445_ (.A(_18621_),
    .X(_18624_));
 sky130_fd_sc_hd__mux2_2 _22446_ (.A0(\cpuregs[1][7] ),
    .A1(_18350_),
    .S(_18624_),
    .X(_03382_));
 sky130_fd_sc_hd__mux2_2 _22447_ (.A0(\cpuregs[1][6] ),
    .A1(_18353_),
    .S(_18624_),
    .X(_03381_));
 sky130_fd_sc_hd__mux2_2 _22448_ (.A0(\cpuregs[1][5] ),
    .A1(_18355_),
    .S(_18624_),
    .X(_03380_));
 sky130_fd_sc_hd__mux2_2 _22449_ (.A0(\cpuregs[1][4] ),
    .A1(_18357_),
    .S(_18624_),
    .X(_03379_));
 sky130_fd_sc_hd__buf_1 _22450_ (.A(_18621_),
    .X(_18625_));
 sky130_fd_sc_hd__mux2_2 _22451_ (.A0(\cpuregs[1][3] ),
    .A1(_18359_),
    .S(_18625_),
    .X(_03378_));
 sky130_fd_sc_hd__mux2_2 _22452_ (.A0(\cpuregs[1][2] ),
    .A1(_18362_),
    .S(_18625_),
    .X(_03377_));
 sky130_fd_sc_hd__mux2_2 _22453_ (.A0(\cpuregs[1][1] ),
    .A1(_18364_),
    .S(_18625_),
    .X(_03376_));
 sky130_fd_sc_hd__mux2_2 _22454_ (.A0(\cpuregs[1][0] ),
    .A1(_18366_),
    .S(_18625_),
    .X(_03375_));
 sky130_fd_sc_hd__buf_1 _22455_ (.A(_18275_),
    .X(_18626_));
 sky130_fd_sc_hd__nand3b_2 _22456_ (.A_N(_18626_),
    .B(_18458_),
    .C(_18549_),
    .Y(_18627_));
 sky130_fd_sc_hd__buf_1 _22457_ (.A(_18627_),
    .X(_18628_));
 sky130_fd_sc_hd__buf_1 _22458_ (.A(_18628_),
    .X(_18629_));
 sky130_fd_sc_hd__mux2_2 _22459_ (.A0(_18546_),
    .A1(\cpuregs[12][31] ),
    .S(_18629_),
    .X(_03374_));
 sky130_fd_sc_hd__mux2_2 _22460_ (.A0(_18554_),
    .A1(\cpuregs[12][30] ),
    .S(_18629_),
    .X(_03373_));
 sky130_fd_sc_hd__mux2_2 _22461_ (.A0(_18555_),
    .A1(\cpuregs[12][29] ),
    .S(_18629_),
    .X(_03372_));
 sky130_fd_sc_hd__mux2_2 _22462_ (.A0(_18556_),
    .A1(\cpuregs[12][28] ),
    .S(_18629_),
    .X(_03371_));
 sky130_fd_sc_hd__buf_1 _22463_ (.A(_18628_),
    .X(_18630_));
 sky130_fd_sc_hd__mux2_2 _22464_ (.A0(_18557_),
    .A1(\cpuregs[12][27] ),
    .S(_18630_),
    .X(_03370_));
 sky130_fd_sc_hd__mux2_2 _22465_ (.A0(_18559_),
    .A1(\cpuregs[12][26] ),
    .S(_18630_),
    .X(_03369_));
 sky130_fd_sc_hd__mux2_2 _22466_ (.A0(_18560_),
    .A1(\cpuregs[12][25] ),
    .S(_18630_),
    .X(_03368_));
 sky130_fd_sc_hd__mux2_2 _22467_ (.A0(_18561_),
    .A1(\cpuregs[12][24] ),
    .S(_18630_),
    .X(_03367_));
 sky130_fd_sc_hd__buf_1 _22468_ (.A(_18628_),
    .X(_18631_));
 sky130_fd_sc_hd__mux2_2 _22469_ (.A0(_18562_),
    .A1(\cpuregs[12][23] ),
    .S(_18631_),
    .X(_03366_));
 sky130_fd_sc_hd__mux2_2 _22470_ (.A0(_18564_),
    .A1(\cpuregs[12][22] ),
    .S(_18631_),
    .X(_03365_));
 sky130_fd_sc_hd__mux2_2 _22471_ (.A0(_18565_),
    .A1(\cpuregs[12][21] ),
    .S(_18631_),
    .X(_03364_));
 sky130_fd_sc_hd__mux2_2 _22472_ (.A0(_18566_),
    .A1(\cpuregs[12][20] ),
    .S(_18631_),
    .X(_03363_));
 sky130_fd_sc_hd__buf_1 _22473_ (.A(_18628_),
    .X(_18632_));
 sky130_fd_sc_hd__mux2_2 _22474_ (.A0(_18567_),
    .A1(\cpuregs[12][19] ),
    .S(_18632_),
    .X(_03362_));
 sky130_fd_sc_hd__mux2_2 _22475_ (.A0(_18569_),
    .A1(\cpuregs[12][18] ),
    .S(_18632_),
    .X(_03361_));
 sky130_fd_sc_hd__mux2_2 _22476_ (.A0(_18570_),
    .A1(\cpuregs[12][17] ),
    .S(_18632_),
    .X(_03360_));
 sky130_fd_sc_hd__mux2_2 _22477_ (.A0(_18571_),
    .A1(\cpuregs[12][16] ),
    .S(_18632_),
    .X(_03359_));
 sky130_fd_sc_hd__buf_1 _22478_ (.A(_18627_),
    .X(_18633_));
 sky130_fd_sc_hd__buf_1 _22479_ (.A(_18633_),
    .X(_18634_));
 sky130_fd_sc_hd__mux2_2 _22480_ (.A0(_18572_),
    .A1(\cpuregs[12][15] ),
    .S(_18634_),
    .X(_03358_));
 sky130_fd_sc_hd__mux2_2 _22481_ (.A0(_18575_),
    .A1(\cpuregs[12][14] ),
    .S(_18634_),
    .X(_03357_));
 sky130_fd_sc_hd__mux2_2 _22482_ (.A0(_18576_),
    .A1(\cpuregs[12][13] ),
    .S(_18634_),
    .X(_03356_));
 sky130_fd_sc_hd__mux2_2 _22483_ (.A0(_18577_),
    .A1(\cpuregs[12][12] ),
    .S(_18634_),
    .X(_03355_));
 sky130_fd_sc_hd__buf_1 _22484_ (.A(_18633_),
    .X(_18635_));
 sky130_fd_sc_hd__mux2_2 _22485_ (.A0(_18578_),
    .A1(\cpuregs[12][11] ),
    .S(_18635_),
    .X(_03354_));
 sky130_fd_sc_hd__mux2_2 _22486_ (.A0(_18580_),
    .A1(\cpuregs[12][10] ),
    .S(_18635_),
    .X(_03353_));
 sky130_fd_sc_hd__mux2_2 _22487_ (.A0(_18581_),
    .A1(\cpuregs[12][9] ),
    .S(_18635_),
    .X(_03352_));
 sky130_fd_sc_hd__mux2_2 _22488_ (.A0(_18582_),
    .A1(\cpuregs[12][8] ),
    .S(_18635_),
    .X(_03351_));
 sky130_fd_sc_hd__buf_1 _22489_ (.A(_18633_),
    .X(_18636_));
 sky130_fd_sc_hd__mux2_2 _22490_ (.A0(_18583_),
    .A1(\cpuregs[12][7] ),
    .S(_18636_),
    .X(_03350_));
 sky130_fd_sc_hd__mux2_2 _22491_ (.A0(_18585_),
    .A1(\cpuregs[12][6] ),
    .S(_18636_),
    .X(_03349_));
 sky130_fd_sc_hd__mux2_2 _22492_ (.A0(_18586_),
    .A1(\cpuregs[12][5] ),
    .S(_18636_),
    .X(_03348_));
 sky130_fd_sc_hd__mux2_2 _22493_ (.A0(_18587_),
    .A1(\cpuregs[12][4] ),
    .S(_18636_),
    .X(_03347_));
 sky130_fd_sc_hd__buf_1 _22494_ (.A(_18633_),
    .X(_18637_));
 sky130_fd_sc_hd__mux2_2 _22495_ (.A0(_18588_),
    .A1(\cpuregs[12][3] ),
    .S(_18637_),
    .X(_03346_));
 sky130_fd_sc_hd__mux2_2 _22496_ (.A0(_18590_),
    .A1(\cpuregs[12][2] ),
    .S(_18637_),
    .X(_03345_));
 sky130_fd_sc_hd__mux2_2 _22497_ (.A0(_18591_),
    .A1(\cpuregs[12][1] ),
    .S(_18637_),
    .X(_03344_));
 sky130_fd_sc_hd__mux2_2 _22498_ (.A0(_18592_),
    .A1(\cpuregs[12][0] ),
    .S(_18637_),
    .X(_03343_));
 sky130_fd_sc_hd__and3b_2 _22499_ (.A_N(_18626_),
    .B(_18293_),
    .C(_18280_),
    .X(_18638_));
 sky130_fd_sc_hd__nand3_2 _22500_ (.A(_18638_),
    .B(_18277_),
    .C(_18278_),
    .Y(_18639_));
 sky130_fd_sc_hd__buf_1 _22501_ (.A(_18639_),
    .X(_18640_));
 sky130_fd_sc_hd__buf_1 _22502_ (.A(_18640_),
    .X(_18641_));
 sky130_fd_sc_hd__mux2_2 _22503_ (.A0(_18546_),
    .A1(\cpuregs[16][31] ),
    .S(_18641_),
    .X(_03342_));
 sky130_fd_sc_hd__mux2_2 _22504_ (.A0(_18554_),
    .A1(\cpuregs[16][30] ),
    .S(_18641_),
    .X(_03341_));
 sky130_fd_sc_hd__mux2_2 _22505_ (.A0(_18555_),
    .A1(\cpuregs[16][29] ),
    .S(_18641_),
    .X(_03340_));
 sky130_fd_sc_hd__mux2_2 _22506_ (.A0(_18556_),
    .A1(\cpuregs[16][28] ),
    .S(_18641_),
    .X(_03339_));
 sky130_fd_sc_hd__buf_1 _22507_ (.A(_18640_),
    .X(_18642_));
 sky130_fd_sc_hd__mux2_2 _22508_ (.A0(_18557_),
    .A1(\cpuregs[16][27] ),
    .S(_18642_),
    .X(_03338_));
 sky130_fd_sc_hd__mux2_2 _22509_ (.A0(_18559_),
    .A1(\cpuregs[16][26] ),
    .S(_18642_),
    .X(_03337_));
 sky130_fd_sc_hd__mux2_2 _22510_ (.A0(_18560_),
    .A1(\cpuregs[16][25] ),
    .S(_18642_),
    .X(_03336_));
 sky130_fd_sc_hd__mux2_2 _22511_ (.A0(_18561_),
    .A1(\cpuregs[16][24] ),
    .S(_18642_),
    .X(_03335_));
 sky130_fd_sc_hd__buf_1 _22512_ (.A(_18640_),
    .X(_18643_));
 sky130_fd_sc_hd__mux2_2 _22513_ (.A0(_18562_),
    .A1(\cpuregs[16][23] ),
    .S(_18643_),
    .X(_03334_));
 sky130_fd_sc_hd__mux2_2 _22514_ (.A0(_18564_),
    .A1(\cpuregs[16][22] ),
    .S(_18643_),
    .X(_03333_));
 sky130_fd_sc_hd__mux2_2 _22515_ (.A0(_18565_),
    .A1(\cpuregs[16][21] ),
    .S(_18643_),
    .X(_03332_));
 sky130_fd_sc_hd__mux2_2 _22516_ (.A0(_18566_),
    .A1(\cpuregs[16][20] ),
    .S(_18643_),
    .X(_03331_));
 sky130_fd_sc_hd__buf_1 _22517_ (.A(_18640_),
    .X(_18644_));
 sky130_fd_sc_hd__mux2_2 _22518_ (.A0(_18567_),
    .A1(\cpuregs[16][19] ),
    .S(_18644_),
    .X(_03330_));
 sky130_fd_sc_hd__mux2_2 _22519_ (.A0(_18569_),
    .A1(\cpuregs[16][18] ),
    .S(_18644_),
    .X(_03329_));
 sky130_fd_sc_hd__mux2_2 _22520_ (.A0(_18570_),
    .A1(\cpuregs[16][17] ),
    .S(_18644_),
    .X(_03328_));
 sky130_fd_sc_hd__mux2_2 _22521_ (.A0(_18571_),
    .A1(\cpuregs[16][16] ),
    .S(_18644_),
    .X(_03327_));
 sky130_fd_sc_hd__buf_1 _22522_ (.A(_18639_),
    .X(_18645_));
 sky130_fd_sc_hd__buf_1 _22523_ (.A(_18645_),
    .X(_18646_));
 sky130_fd_sc_hd__mux2_2 _22524_ (.A0(_18572_),
    .A1(\cpuregs[16][15] ),
    .S(_18646_),
    .X(_03326_));
 sky130_fd_sc_hd__mux2_2 _22525_ (.A0(_18575_),
    .A1(\cpuregs[16][14] ),
    .S(_18646_),
    .X(_03325_));
 sky130_fd_sc_hd__mux2_2 _22526_ (.A0(_18576_),
    .A1(\cpuregs[16][13] ),
    .S(_18646_),
    .X(_03324_));
 sky130_fd_sc_hd__mux2_2 _22527_ (.A0(_18577_),
    .A1(\cpuregs[16][12] ),
    .S(_18646_),
    .X(_03323_));
 sky130_fd_sc_hd__buf_1 _22528_ (.A(_18645_),
    .X(_18647_));
 sky130_fd_sc_hd__mux2_2 _22529_ (.A0(_18578_),
    .A1(\cpuregs[16][11] ),
    .S(_18647_),
    .X(_03322_));
 sky130_fd_sc_hd__mux2_2 _22530_ (.A0(_18580_),
    .A1(\cpuregs[16][10] ),
    .S(_18647_),
    .X(_03321_));
 sky130_fd_sc_hd__mux2_2 _22531_ (.A0(_18581_),
    .A1(\cpuregs[16][9] ),
    .S(_18647_),
    .X(_03320_));
 sky130_fd_sc_hd__mux2_2 _22532_ (.A0(_18582_),
    .A1(\cpuregs[16][8] ),
    .S(_18647_),
    .X(_03319_));
 sky130_fd_sc_hd__buf_1 _22533_ (.A(_18645_),
    .X(_18648_));
 sky130_fd_sc_hd__mux2_2 _22534_ (.A0(_18583_),
    .A1(\cpuregs[16][7] ),
    .S(_18648_),
    .X(_03318_));
 sky130_fd_sc_hd__mux2_2 _22535_ (.A0(_18585_),
    .A1(\cpuregs[16][6] ),
    .S(_18648_),
    .X(_03317_));
 sky130_fd_sc_hd__mux2_2 _22536_ (.A0(_18586_),
    .A1(\cpuregs[16][5] ),
    .S(_18648_),
    .X(_03316_));
 sky130_fd_sc_hd__mux2_2 _22537_ (.A0(_18587_),
    .A1(\cpuregs[16][4] ),
    .S(_18648_),
    .X(_03315_));
 sky130_fd_sc_hd__buf_1 _22538_ (.A(_18645_),
    .X(_18649_));
 sky130_fd_sc_hd__mux2_2 _22539_ (.A0(_18588_),
    .A1(\cpuregs[16][3] ),
    .S(_18649_),
    .X(_03314_));
 sky130_fd_sc_hd__mux2_2 _22540_ (.A0(_18590_),
    .A1(\cpuregs[16][2] ),
    .S(_18649_),
    .X(_03313_));
 sky130_fd_sc_hd__mux2_2 _22541_ (.A0(_18591_),
    .A1(\cpuregs[16][1] ),
    .S(_18649_),
    .X(_03312_));
 sky130_fd_sc_hd__mux2_2 _22542_ (.A0(_18592_),
    .A1(\cpuregs[16][0] ),
    .S(_18649_),
    .X(_03311_));
 sky130_fd_sc_hd__buf_1 _22543_ (.A(\cpuregs_wrdata[31] ),
    .X(_18650_));
 sky130_fd_sc_hd__o2111ai_2 _22544_ (.A1(_18528_),
    .A2(_18547_),
    .B1(_18370_),
    .C1(_18501_),
    .D1(_18550_),
    .Y(_18651_));
 sky130_fd_sc_hd__buf_1 _22545_ (.A(_18651_),
    .X(_18652_));
 sky130_fd_sc_hd__buf_1 _22546_ (.A(_18652_),
    .X(_18653_));
 sky130_fd_sc_hd__mux2_2 _22547_ (.A0(_18650_),
    .A1(\cpuregs[17][31] ),
    .S(_18653_),
    .X(_03310_));
 sky130_fd_sc_hd__buf_1 _22548_ (.A(\cpuregs_wrdata[30] ),
    .X(_18654_));
 sky130_fd_sc_hd__mux2_2 _22549_ (.A0(_18654_),
    .A1(\cpuregs[17][30] ),
    .S(_18653_),
    .X(_03309_));
 sky130_fd_sc_hd__buf_1 _22550_ (.A(\cpuregs_wrdata[29] ),
    .X(_18655_));
 sky130_fd_sc_hd__mux2_2 _22551_ (.A0(_18655_),
    .A1(\cpuregs[17][29] ),
    .S(_18653_),
    .X(_03308_));
 sky130_fd_sc_hd__buf_1 _22552_ (.A(\cpuregs_wrdata[28] ),
    .X(_18656_));
 sky130_fd_sc_hd__mux2_2 _22553_ (.A0(_18656_),
    .A1(\cpuregs[17][28] ),
    .S(_18653_),
    .X(_03307_));
 sky130_fd_sc_hd__buf_1 _22554_ (.A(\cpuregs_wrdata[27] ),
    .X(_18657_));
 sky130_fd_sc_hd__buf_1 _22555_ (.A(_18652_),
    .X(_18658_));
 sky130_fd_sc_hd__mux2_2 _22556_ (.A0(_18657_),
    .A1(\cpuregs[17][27] ),
    .S(_18658_),
    .X(_03306_));
 sky130_fd_sc_hd__buf_1 _22557_ (.A(\cpuregs_wrdata[26] ),
    .X(_18659_));
 sky130_fd_sc_hd__mux2_2 _22558_ (.A0(_18659_),
    .A1(\cpuregs[17][26] ),
    .S(_18658_),
    .X(_03305_));
 sky130_fd_sc_hd__buf_1 _22559_ (.A(\cpuregs_wrdata[25] ),
    .X(_18660_));
 sky130_fd_sc_hd__mux2_2 _22560_ (.A0(_18660_),
    .A1(\cpuregs[17][25] ),
    .S(_18658_),
    .X(_03304_));
 sky130_fd_sc_hd__buf_1 _22561_ (.A(\cpuregs_wrdata[24] ),
    .X(_18661_));
 sky130_fd_sc_hd__mux2_2 _22562_ (.A0(_18661_),
    .A1(\cpuregs[17][24] ),
    .S(_18658_),
    .X(_03303_));
 sky130_fd_sc_hd__buf_1 _22563_ (.A(\cpuregs_wrdata[23] ),
    .X(_18662_));
 sky130_fd_sc_hd__buf_1 _22564_ (.A(_18652_),
    .X(_18663_));
 sky130_fd_sc_hd__mux2_2 _22565_ (.A0(_18662_),
    .A1(\cpuregs[17][23] ),
    .S(_18663_),
    .X(_03302_));
 sky130_fd_sc_hd__buf_1 _22566_ (.A(\cpuregs_wrdata[22] ),
    .X(_18664_));
 sky130_fd_sc_hd__mux2_2 _22567_ (.A0(_18664_),
    .A1(\cpuregs[17][22] ),
    .S(_18663_),
    .X(_03301_));
 sky130_fd_sc_hd__buf_1 _22568_ (.A(\cpuregs_wrdata[21] ),
    .X(_18665_));
 sky130_fd_sc_hd__mux2_2 _22569_ (.A0(_18665_),
    .A1(\cpuregs[17][21] ),
    .S(_18663_),
    .X(_03300_));
 sky130_fd_sc_hd__buf_1 _22570_ (.A(\cpuregs_wrdata[20] ),
    .X(_18666_));
 sky130_fd_sc_hd__mux2_2 _22571_ (.A0(_18666_),
    .A1(\cpuregs[17][20] ),
    .S(_18663_),
    .X(_03299_));
 sky130_fd_sc_hd__buf_1 _22572_ (.A(\cpuregs_wrdata[19] ),
    .X(_18667_));
 sky130_fd_sc_hd__buf_1 _22573_ (.A(_18652_),
    .X(_18668_));
 sky130_fd_sc_hd__mux2_2 _22574_ (.A0(_18667_),
    .A1(\cpuregs[17][19] ),
    .S(_18668_),
    .X(_03298_));
 sky130_fd_sc_hd__buf_1 _22575_ (.A(\cpuregs_wrdata[18] ),
    .X(_18669_));
 sky130_fd_sc_hd__mux2_2 _22576_ (.A0(_18669_),
    .A1(\cpuregs[17][18] ),
    .S(_18668_),
    .X(_03297_));
 sky130_fd_sc_hd__buf_1 _22577_ (.A(\cpuregs_wrdata[17] ),
    .X(_18670_));
 sky130_fd_sc_hd__mux2_2 _22578_ (.A0(_18670_),
    .A1(\cpuregs[17][17] ),
    .S(_18668_),
    .X(_03296_));
 sky130_fd_sc_hd__buf_1 _22579_ (.A(\cpuregs_wrdata[16] ),
    .X(_18671_));
 sky130_fd_sc_hd__mux2_2 _22580_ (.A0(_18671_),
    .A1(\cpuregs[17][16] ),
    .S(_18668_),
    .X(_03295_));
 sky130_fd_sc_hd__buf_1 _22581_ (.A(\cpuregs_wrdata[15] ),
    .X(_18672_));
 sky130_fd_sc_hd__buf_1 _22582_ (.A(_18651_),
    .X(_18673_));
 sky130_fd_sc_hd__buf_1 _22583_ (.A(_18673_),
    .X(_18674_));
 sky130_fd_sc_hd__mux2_2 _22584_ (.A0(_18672_),
    .A1(\cpuregs[17][15] ),
    .S(_18674_),
    .X(_03294_));
 sky130_fd_sc_hd__buf_1 _22585_ (.A(\cpuregs_wrdata[14] ),
    .X(_18675_));
 sky130_fd_sc_hd__mux2_2 _22586_ (.A0(_18675_),
    .A1(\cpuregs[17][14] ),
    .S(_18674_),
    .X(_03293_));
 sky130_fd_sc_hd__buf_1 _22587_ (.A(\cpuregs_wrdata[13] ),
    .X(_18676_));
 sky130_fd_sc_hd__mux2_2 _22588_ (.A0(_18676_),
    .A1(\cpuregs[17][13] ),
    .S(_18674_),
    .X(_03292_));
 sky130_fd_sc_hd__buf_1 _22589_ (.A(\cpuregs_wrdata[12] ),
    .X(_18677_));
 sky130_fd_sc_hd__mux2_2 _22590_ (.A0(_18677_),
    .A1(\cpuregs[17][12] ),
    .S(_18674_),
    .X(_03291_));
 sky130_fd_sc_hd__buf_1 _22591_ (.A(\cpuregs_wrdata[11] ),
    .X(_18678_));
 sky130_fd_sc_hd__buf_1 _22592_ (.A(_18673_),
    .X(_18679_));
 sky130_fd_sc_hd__mux2_2 _22593_ (.A0(_18678_),
    .A1(\cpuregs[17][11] ),
    .S(_18679_),
    .X(_03290_));
 sky130_fd_sc_hd__buf_1 _22594_ (.A(\cpuregs_wrdata[10] ),
    .X(_18680_));
 sky130_fd_sc_hd__mux2_2 _22595_ (.A0(_18680_),
    .A1(\cpuregs[17][10] ),
    .S(_18679_),
    .X(_03289_));
 sky130_fd_sc_hd__buf_1 _22596_ (.A(\cpuregs_wrdata[9] ),
    .X(_18681_));
 sky130_fd_sc_hd__mux2_2 _22597_ (.A0(_18681_),
    .A1(\cpuregs[17][9] ),
    .S(_18679_),
    .X(_03288_));
 sky130_fd_sc_hd__buf_1 _22598_ (.A(\cpuregs_wrdata[8] ),
    .X(_18682_));
 sky130_fd_sc_hd__mux2_2 _22599_ (.A0(_18682_),
    .A1(\cpuregs[17][8] ),
    .S(_18679_),
    .X(_03287_));
 sky130_fd_sc_hd__buf_1 _22600_ (.A(\cpuregs_wrdata[7] ),
    .X(_18683_));
 sky130_fd_sc_hd__buf_1 _22601_ (.A(_18673_),
    .X(_18684_));
 sky130_fd_sc_hd__mux2_2 _22602_ (.A0(_18683_),
    .A1(\cpuregs[17][7] ),
    .S(_18684_),
    .X(_03286_));
 sky130_fd_sc_hd__buf_1 _22603_ (.A(\cpuregs_wrdata[6] ),
    .X(_18685_));
 sky130_fd_sc_hd__mux2_2 _22604_ (.A0(_18685_),
    .A1(\cpuregs[17][6] ),
    .S(_18684_),
    .X(_03285_));
 sky130_fd_sc_hd__buf_1 _22605_ (.A(\cpuregs_wrdata[5] ),
    .X(_18686_));
 sky130_fd_sc_hd__mux2_2 _22606_ (.A0(_18686_),
    .A1(\cpuregs[17][5] ),
    .S(_18684_),
    .X(_03284_));
 sky130_fd_sc_hd__buf_1 _22607_ (.A(\cpuregs_wrdata[4] ),
    .X(_18687_));
 sky130_fd_sc_hd__mux2_2 _22608_ (.A0(_18687_),
    .A1(\cpuregs[17][4] ),
    .S(_18684_),
    .X(_03283_));
 sky130_fd_sc_hd__buf_1 _22609_ (.A(\cpuregs_wrdata[3] ),
    .X(_18688_));
 sky130_fd_sc_hd__buf_1 _22610_ (.A(_18673_),
    .X(_18689_));
 sky130_fd_sc_hd__mux2_2 _22611_ (.A0(_18688_),
    .A1(\cpuregs[17][3] ),
    .S(_18689_),
    .X(_03282_));
 sky130_fd_sc_hd__buf_1 _22612_ (.A(\cpuregs_wrdata[2] ),
    .X(_18690_));
 sky130_fd_sc_hd__mux2_2 _22613_ (.A0(_18690_),
    .A1(\cpuregs[17][2] ),
    .S(_18689_),
    .X(_03281_));
 sky130_fd_sc_hd__buf_1 _22614_ (.A(\cpuregs_wrdata[1] ),
    .X(_18691_));
 sky130_fd_sc_hd__mux2_2 _22615_ (.A0(_18691_),
    .A1(\cpuregs[17][1] ),
    .S(_18689_),
    .X(_03280_));
 sky130_fd_sc_hd__buf_1 _22616_ (.A(\cpuregs_wrdata[0] ),
    .X(_18692_));
 sky130_fd_sc_hd__mux2_2 _22617_ (.A0(_18692_),
    .A1(\cpuregs[17][0] ),
    .S(_18689_),
    .X(_03279_));
 sky130_fd_sc_hd__buf_1 _22618_ (.A(\pcpi_mul.rs2[31] ),
    .X(_18693_));
 sky130_fd_sc_hd__buf_1 _22619_ (.A(_18693_),
    .X(_18694_));
 sky130_fd_sc_hd__buf_1 _22620_ (.A(_18694_),
    .X(_18695_));
 sky130_fd_sc_hd__buf_1 _22621_ (.A(_18695_),
    .X(_18696_));
 sky130_fd_sc_hd__buf_1 _22622_ (.A(_18696_),
    .X(_18697_));
 sky130_fd_sc_hd__buf_1 _22623_ (.A(_18697_),
    .X(_18698_));
 sky130_vsdinv _22624_ (.A(_16955_),
    .Y(_18699_));
 sky130_fd_sc_hd__buf_1 _22625_ (.A(_18699_),
    .X(_18700_));
 sky130_fd_sc_hd__buf_1 _22626_ (.A(_18700_),
    .X(_18701_));
 sky130_fd_sc_hd__and2_2 _22627_ (.A(_16974_),
    .B(_16978_),
    .X(_18702_));
 sky130_fd_sc_hd__a21o_2 _22628_ (.A1(_18698_),
    .A2(_18701_),
    .B1(_18702_),
    .X(_03278_));
 sky130_fd_sc_hd__buf_1 _22629_ (.A(\pcpi_mul.rs2[30] ),
    .X(_18703_));
 sky130_fd_sc_hd__buf_1 _22630_ (.A(_18703_),
    .X(_18704_));
 sky130_fd_sc_hd__buf_1 _22631_ (.A(_18704_),
    .X(_18705_));
 sky130_fd_sc_hd__buf_1 _22632_ (.A(_18705_),
    .X(_18706_));
 sky130_fd_sc_hd__buf_1 _22633_ (.A(_18706_),
    .X(_18707_));
 sky130_vsdinv _22634_ (.A(_18707_),
    .Y(_18708_));
 sky130_fd_sc_hd__nand2_2 _22635_ (.A(_16966_),
    .B(_18385_),
    .Y(_18709_));
 sky130_fd_sc_hd__o21ai_2 _22636_ (.A1(_18708_),
    .A2(_03728_),
    .B1(_18709_),
    .Y(_03277_));
 sky130_fd_sc_hd__buf_1 _22637_ (.A(\pcpi_mul.rs2[29] ),
    .X(_18710_));
 sky130_fd_sc_hd__buf_1 _22638_ (.A(_18710_),
    .X(_18711_));
 sky130_fd_sc_hd__buf_1 _22639_ (.A(_18711_),
    .X(_18712_));
 sky130_fd_sc_hd__buf_1 _22640_ (.A(_18712_),
    .X(_18713_));
 sky130_fd_sc_hd__buf_1 _22641_ (.A(_18713_),
    .X(_18714_));
 sky130_fd_sc_hd__and2_2 _22642_ (.A(_16974_),
    .B(_18387_),
    .X(_18715_));
 sky130_fd_sc_hd__a21o_2 _22643_ (.A1(_18714_),
    .A2(_18701_),
    .B1(_18715_),
    .X(_03276_));
 sky130_fd_sc_hd__buf_1 _22644_ (.A(\pcpi_mul.rs2[28] ),
    .X(_18716_));
 sky130_fd_sc_hd__buf_1 _22645_ (.A(_18716_),
    .X(_18717_));
 sky130_fd_sc_hd__buf_1 _22646_ (.A(_18717_),
    .X(_18718_));
 sky130_fd_sc_hd__buf_1 _22647_ (.A(_18718_),
    .X(_18719_));
 sky130_fd_sc_hd__buf_1 _22648_ (.A(_18719_),
    .X(_18720_));
 sky130_fd_sc_hd__and2_2 _22649_ (.A(_16974_),
    .B(_18388_),
    .X(_18721_));
 sky130_fd_sc_hd__a21o_2 _22650_ (.A1(_18720_),
    .A2(_18701_),
    .B1(_18721_),
    .X(_03275_));
 sky130_fd_sc_hd__buf_1 _22651_ (.A(\pcpi_mul.rs2[27] ),
    .X(_18722_));
 sky130_fd_sc_hd__buf_1 _22652_ (.A(_18722_),
    .X(_18723_));
 sky130_vsdinv _22653_ (.A(_18723_),
    .Y(_18724_));
 sky130_fd_sc_hd__buf_1 _22654_ (.A(_18724_),
    .X(_18725_));
 sky130_fd_sc_hd__nand2_2 _22655_ (.A(_16966_),
    .B(_18391_),
    .Y(_18726_));
 sky130_fd_sc_hd__o21ai_2 _22656_ (.A1(_18725_),
    .A2(_03728_),
    .B1(_18726_),
    .Y(_03274_));
 sky130_fd_sc_hd__buf_1 _22657_ (.A(\pcpi_mul.rs2[26] ),
    .X(_18727_));
 sky130_fd_sc_hd__buf_1 _22658_ (.A(_18727_),
    .X(_18728_));
 sky130_fd_sc_hd__buf_1 _22659_ (.A(_18728_),
    .X(_18729_));
 sky130_fd_sc_hd__buf_1 _22660_ (.A(_18729_),
    .X(_18730_));
 sky130_fd_sc_hd__buf_1 _22661_ (.A(_16955_),
    .X(_18731_));
 sky130_fd_sc_hd__buf_1 _22662_ (.A(_18731_),
    .X(_18732_));
 sky130_fd_sc_hd__and2_2 _22663_ (.A(_18732_),
    .B(_18393_),
    .X(_18733_));
 sky130_fd_sc_hd__a21o_2 _22664_ (.A1(_18730_),
    .A2(_18701_),
    .B1(_18733_),
    .X(_03273_));
 sky130_fd_sc_hd__buf_1 _22665_ (.A(\pcpi_mul.rs2[25] ),
    .X(_18734_));
 sky130_fd_sc_hd__buf_1 _22666_ (.A(_18734_),
    .X(_18735_));
 sky130_fd_sc_hd__buf_1 _22667_ (.A(_18735_),
    .X(_18736_));
 sky130_fd_sc_hd__buf_1 _22668_ (.A(_18736_),
    .X(_18737_));
 sky130_fd_sc_hd__buf_1 _22669_ (.A(_18700_),
    .X(_18738_));
 sky130_fd_sc_hd__and2_2 _22670_ (.A(_18732_),
    .B(_18395_),
    .X(_18739_));
 sky130_fd_sc_hd__a21o_2 _22671_ (.A1(_18737_),
    .A2(_18738_),
    .B1(_18739_),
    .X(_03272_));
 sky130_vsdinv _22672_ (.A(\pcpi_mul.rs2[24] ),
    .Y(_18740_));
 sky130_fd_sc_hd__buf_1 _22673_ (.A(_18740_),
    .X(_18741_));
 sky130_fd_sc_hd__buf_1 _22674_ (.A(_18741_),
    .X(_18742_));
 sky130_fd_sc_hd__buf_1 _22675_ (.A(_18742_),
    .X(_18743_));
 sky130_fd_sc_hd__buf_1 _22676_ (.A(_16975_),
    .X(_18744_));
 sky130_fd_sc_hd__buf_1 _22677_ (.A(_16965_),
    .X(_18745_));
 sky130_fd_sc_hd__nand2_2 _22678_ (.A(_18745_),
    .B(_18396_),
    .Y(_18746_));
 sky130_fd_sc_hd__o21ai_2 _22679_ (.A1(_18743_),
    .A2(_18744_),
    .B1(_18746_),
    .Y(_03271_));
 sky130_fd_sc_hd__buf_1 _22680_ (.A(\pcpi_mul.rs2[23] ),
    .X(_18747_));
 sky130_fd_sc_hd__buf_1 _22681_ (.A(_18747_),
    .X(_18748_));
 sky130_fd_sc_hd__buf_1 _22682_ (.A(_18748_),
    .X(_18749_));
 sky130_fd_sc_hd__buf_1 _22683_ (.A(_18749_),
    .X(_18750_));
 sky130_fd_sc_hd__and2_2 _22684_ (.A(_18732_),
    .B(_18399_),
    .X(_18751_));
 sky130_fd_sc_hd__a21o_2 _22685_ (.A1(_18750_),
    .A2(_18738_),
    .B1(_18751_),
    .X(_03270_));
 sky130_fd_sc_hd__buf_1 _22686_ (.A(\pcpi_mul.rs2[22] ),
    .X(_18752_));
 sky130_fd_sc_hd__buf_1 _22687_ (.A(_18752_),
    .X(_18753_));
 sky130_fd_sc_hd__buf_1 _22688_ (.A(_18753_),
    .X(_18754_));
 sky130_fd_sc_hd__buf_1 _22689_ (.A(_18754_),
    .X(_18755_));
 sky130_fd_sc_hd__buf_1 _22690_ (.A(_18755_),
    .X(_18756_));
 sky130_fd_sc_hd__and2_2 _22691_ (.A(_18732_),
    .B(_18401_),
    .X(_18757_));
 sky130_fd_sc_hd__a21o_2 _22692_ (.A1(_18756_),
    .A2(_18738_),
    .B1(_18757_),
    .X(_03269_));
 sky130_fd_sc_hd__buf_1 _22693_ (.A(\pcpi_mul.rs2[21] ),
    .X(_18758_));
 sky130_vsdinv _22694_ (.A(_18758_),
    .Y(_18759_));
 sky130_fd_sc_hd__buf_1 _22695_ (.A(_18759_),
    .X(_18760_));
 sky130_fd_sc_hd__buf_1 _22696_ (.A(_18760_),
    .X(_18761_));
 sky130_fd_sc_hd__nand2_2 _22697_ (.A(_18745_),
    .B(_18403_),
    .Y(_18762_));
 sky130_fd_sc_hd__o21ai_2 _22698_ (.A1(_18761_),
    .A2(_18744_),
    .B1(_18762_),
    .Y(_03268_));
 sky130_fd_sc_hd__buf_1 _22699_ (.A(\pcpi_mul.rs2[20] ),
    .X(_18763_));
 sky130_fd_sc_hd__buf_1 _22700_ (.A(_18763_),
    .X(_18764_));
 sky130_fd_sc_hd__buf_1 _22701_ (.A(_18764_),
    .X(_18765_));
 sky130_fd_sc_hd__buf_1 _22702_ (.A(_18765_),
    .X(_18766_));
 sky130_fd_sc_hd__buf_1 _22703_ (.A(_18731_),
    .X(_18767_));
 sky130_fd_sc_hd__and2_2 _22704_ (.A(_18767_),
    .B(_18404_),
    .X(_18768_));
 sky130_fd_sc_hd__a21o_2 _22705_ (.A1(_18766_),
    .A2(_18738_),
    .B1(_18768_),
    .X(_03267_));
 sky130_fd_sc_hd__buf_1 _22706_ (.A(\pcpi_mul.rs2[19] ),
    .X(_18769_));
 sky130_fd_sc_hd__buf_1 _22707_ (.A(_18769_),
    .X(_18770_));
 sky130_fd_sc_hd__buf_1 _22708_ (.A(_18770_),
    .X(_18771_));
 sky130_fd_sc_hd__buf_1 _22709_ (.A(_18771_),
    .X(_18772_));
 sky130_fd_sc_hd__buf_1 _22710_ (.A(_18700_),
    .X(_18773_));
 sky130_fd_sc_hd__and2_2 _22711_ (.A(_18767_),
    .B(_18407_),
    .X(_18774_));
 sky130_fd_sc_hd__a21o_2 _22712_ (.A1(_18772_),
    .A2(_18773_),
    .B1(_18774_),
    .X(_03266_));
 sky130_fd_sc_hd__buf_1 _22713_ (.A(\pcpi_mul.rs2[18] ),
    .X(_18775_));
 sky130_vsdinv _22714_ (.A(_18775_),
    .Y(_18776_));
 sky130_fd_sc_hd__buf_1 _22715_ (.A(_18776_),
    .X(_18777_));
 sky130_fd_sc_hd__nand2_2 _22716_ (.A(_18745_),
    .B(_18409_),
    .Y(_18778_));
 sky130_fd_sc_hd__o21ai_2 _22717_ (.A1(_18777_),
    .A2(_18744_),
    .B1(_18778_),
    .Y(_03265_));
 sky130_fd_sc_hd__buf_1 _22718_ (.A(\pcpi_mul.rs2[17] ),
    .X(_18779_));
 sky130_fd_sc_hd__buf_1 _22719_ (.A(_18779_),
    .X(_18780_));
 sky130_fd_sc_hd__buf_1 _22720_ (.A(_18780_),
    .X(_18781_));
 sky130_vsdinv _22721_ (.A(_18781_),
    .Y(_18782_));
 sky130_fd_sc_hd__nand2_2 _22722_ (.A(_18745_),
    .B(_18411_),
    .Y(_18783_));
 sky130_fd_sc_hd__o21ai_2 _22723_ (.A1(_18782_),
    .A2(_18744_),
    .B1(_18783_),
    .Y(_03264_));
 sky130_fd_sc_hd__buf_1 _22724_ (.A(\pcpi_mul.rs2[16] ),
    .X(_18784_));
 sky130_fd_sc_hd__buf_1 _22725_ (.A(_18784_),
    .X(_18785_));
 sky130_fd_sc_hd__buf_1 _22726_ (.A(_18785_),
    .X(_18786_));
 sky130_fd_sc_hd__buf_1 _22727_ (.A(_18786_),
    .X(_18787_));
 sky130_fd_sc_hd__and2_2 _22728_ (.A(_18767_),
    .B(_18412_),
    .X(_18788_));
 sky130_fd_sc_hd__a21o_2 _22729_ (.A1(_18787_),
    .A2(_18773_),
    .B1(_18788_),
    .X(_03263_));
 sky130_fd_sc_hd__buf_1 _22730_ (.A(\pcpi_mul.rs2[15] ),
    .X(_18789_));
 sky130_fd_sc_hd__buf_1 _22731_ (.A(_18789_),
    .X(_18790_));
 sky130_vsdinv _22732_ (.A(_18790_),
    .Y(_18791_));
 sky130_fd_sc_hd__buf_1 _22733_ (.A(_18791_),
    .X(_18792_));
 sky130_fd_sc_hd__buf_1 _22734_ (.A(_18792_),
    .X(_18793_));
 sky130_fd_sc_hd__buf_1 _22735_ (.A(_16975_),
    .X(_18794_));
 sky130_fd_sc_hd__buf_1 _22736_ (.A(_16965_),
    .X(_18795_));
 sky130_fd_sc_hd__nand2_2 _22737_ (.A(_18795_),
    .B(_18416_),
    .Y(_18796_));
 sky130_fd_sc_hd__o21ai_2 _22738_ (.A1(_18793_),
    .A2(_18794_),
    .B1(_18796_),
    .Y(_03262_));
 sky130_fd_sc_hd__buf_1 _22739_ (.A(\pcpi_mul.rs2[14] ),
    .X(_18797_));
 sky130_fd_sc_hd__buf_1 _22740_ (.A(_18797_),
    .X(_18798_));
 sky130_fd_sc_hd__buf_1 _22741_ (.A(_18798_),
    .X(_18799_));
 sky130_fd_sc_hd__and2_2 _22742_ (.A(_18767_),
    .B(_18418_),
    .X(_18800_));
 sky130_fd_sc_hd__a21o_2 _22743_ (.A1(_18799_),
    .A2(_18773_),
    .B1(_18800_),
    .X(_03261_));
 sky130_fd_sc_hd__buf_1 _22744_ (.A(\pcpi_mul.rs2[13] ),
    .X(_18801_));
 sky130_fd_sc_hd__buf_1 _22745_ (.A(_18801_),
    .X(_18802_));
 sky130_fd_sc_hd__buf_1 _22746_ (.A(_18802_),
    .X(_18803_));
 sky130_fd_sc_hd__buf_1 _22747_ (.A(_18803_),
    .X(_18804_));
 sky130_fd_sc_hd__buf_1 _22748_ (.A(_18731_),
    .X(_18805_));
 sky130_fd_sc_hd__and2_2 _22749_ (.A(_18805_),
    .B(_18420_),
    .X(_18806_));
 sky130_fd_sc_hd__a21o_2 _22750_ (.A1(_18804_),
    .A2(_18773_),
    .B1(_18806_),
    .X(_03260_));
 sky130_fd_sc_hd__buf_1 _22751_ (.A(\pcpi_mul.rs2[12] ),
    .X(_18807_));
 sky130_fd_sc_hd__buf_1 _22752_ (.A(_18807_),
    .X(_18808_));
 sky130_vsdinv _22753_ (.A(_18808_),
    .Y(_18809_));
 sky130_fd_sc_hd__buf_1 _22754_ (.A(_18809_),
    .X(_18810_));
 sky130_fd_sc_hd__buf_1 _22755_ (.A(_18810_),
    .X(_18811_));
 sky130_fd_sc_hd__nand2_2 _22756_ (.A(_18795_),
    .B(_18421_),
    .Y(_18812_));
 sky130_fd_sc_hd__o21ai_2 _22757_ (.A1(_18811_),
    .A2(_18794_),
    .B1(_18812_),
    .Y(_03259_));
 sky130_fd_sc_hd__buf_1 _22758_ (.A(\pcpi_mul.rs2[11] ),
    .X(_18813_));
 sky130_fd_sc_hd__buf_1 _22759_ (.A(_18813_),
    .X(_18814_));
 sky130_fd_sc_hd__buf_1 _22760_ (.A(_18814_),
    .X(_18815_));
 sky130_fd_sc_hd__buf_1 _22761_ (.A(_18699_),
    .X(_18816_));
 sky130_fd_sc_hd__and2_2 _22762_ (.A(_18805_),
    .B(_18424_),
    .X(_18817_));
 sky130_fd_sc_hd__a21o_2 _22763_ (.A1(_18815_),
    .A2(_18816_),
    .B1(_18817_),
    .X(_03258_));
 sky130_fd_sc_hd__buf_1 _22764_ (.A(\pcpi_mul.rs2[10] ),
    .X(_18818_));
 sky130_fd_sc_hd__buf_1 _22765_ (.A(_18818_),
    .X(_18819_));
 sky130_fd_sc_hd__buf_1 _22766_ (.A(_18819_),
    .X(_18820_));
 sky130_fd_sc_hd__and2_2 _22767_ (.A(_18805_),
    .B(_18426_),
    .X(_18821_));
 sky130_fd_sc_hd__a21o_2 _22768_ (.A1(_18820_),
    .A2(_18816_),
    .B1(_18821_),
    .X(_03257_));
 sky130_fd_sc_hd__buf_1 _22769_ (.A(\pcpi_mul.rs2[9] ),
    .X(_18822_));
 sky130_vsdinv _22770_ (.A(_18822_),
    .Y(_18823_));
 sky130_fd_sc_hd__buf_1 _22771_ (.A(_18823_),
    .X(_18824_));
 sky130_fd_sc_hd__buf_1 _22772_ (.A(_18824_),
    .X(_18825_));
 sky130_fd_sc_hd__nand2_2 _22773_ (.A(_18795_),
    .B(_18428_),
    .Y(_18826_));
 sky130_fd_sc_hd__o21ai_2 _22774_ (.A1(_18825_),
    .A2(_18794_),
    .B1(_18826_),
    .Y(_03256_));
 sky130_fd_sc_hd__buf_1 _22775_ (.A(\pcpi_mul.rs2[8] ),
    .X(_18827_));
 sky130_fd_sc_hd__buf_1 _22776_ (.A(_18827_),
    .X(_18828_));
 sky130_fd_sc_hd__buf_1 _22777_ (.A(_18828_),
    .X(_18829_));
 sky130_fd_sc_hd__buf_1 _22778_ (.A(_18829_),
    .X(_18830_));
 sky130_fd_sc_hd__and2_2 _22779_ (.A(_18805_),
    .B(_18430_),
    .X(_18831_));
 sky130_fd_sc_hd__a21o_2 _22780_ (.A1(_18830_),
    .A2(_18816_),
    .B1(_18831_),
    .X(_03255_));
 sky130_fd_sc_hd__buf_1 _22781_ (.A(\pcpi_mul.rs2[7] ),
    .X(_18832_));
 sky130_fd_sc_hd__buf_1 _22782_ (.A(_18832_),
    .X(_18833_));
 sky130_fd_sc_hd__buf_1 _22783_ (.A(_18833_),
    .X(_18834_));
 sky130_fd_sc_hd__buf_1 _22784_ (.A(_18834_),
    .X(_18835_));
 sky130_fd_sc_hd__buf_1 _22785_ (.A(_18731_),
    .X(_18836_));
 sky130_fd_sc_hd__and2_2 _22786_ (.A(_18836_),
    .B(_18433_),
    .X(_18837_));
 sky130_fd_sc_hd__a21o_2 _22787_ (.A1(_18835_),
    .A2(_18816_),
    .B1(_18837_),
    .X(_03254_));
 sky130_fd_sc_hd__buf_1 _22788_ (.A(\pcpi_mul.rs2[6] ),
    .X(_18838_));
 sky130_vsdinv _22789_ (.A(_18838_),
    .Y(_18839_));
 sky130_fd_sc_hd__buf_1 _22790_ (.A(_18839_),
    .X(_18840_));
 sky130_fd_sc_hd__buf_1 _22791_ (.A(_18840_),
    .X(_18841_));
 sky130_fd_sc_hd__nand2_2 _22792_ (.A(_18795_),
    .B(_18436_),
    .Y(_18842_));
 sky130_fd_sc_hd__o21ai_2 _22793_ (.A1(_18841_),
    .A2(_18794_),
    .B1(_18842_),
    .Y(_03253_));
 sky130_fd_sc_hd__buf_1 _22794_ (.A(\pcpi_mul.rs2[5] ),
    .X(_18843_));
 sky130_fd_sc_hd__buf_1 _22795_ (.A(_18843_),
    .X(_18844_));
 sky130_fd_sc_hd__buf_1 _22796_ (.A(_18844_),
    .X(_18845_));
 sky130_fd_sc_hd__buf_1 _22797_ (.A(_18699_),
    .X(_18846_));
 sky130_fd_sc_hd__and2_2 _22798_ (.A(_18836_),
    .B(_18439_),
    .X(_18847_));
 sky130_fd_sc_hd__a21o_2 _22799_ (.A1(_18845_),
    .A2(_18846_),
    .B1(_18847_),
    .X(_03252_));
 sky130_fd_sc_hd__buf_1 _22800_ (.A(\pcpi_mul.rs2[4] ),
    .X(_18848_));
 sky130_fd_sc_hd__buf_1 _22801_ (.A(_18848_),
    .X(_18849_));
 sky130_fd_sc_hd__buf_1 _22802_ (.A(_18849_),
    .X(_18850_));
 sky130_fd_sc_hd__buf_1 _22803_ (.A(_18850_),
    .X(_18851_));
 sky130_fd_sc_hd__buf_1 _22804_ (.A(_18441_),
    .X(_18852_));
 sky130_fd_sc_hd__and2_2 _22805_ (.A(_18836_),
    .B(_18852_),
    .X(_18853_));
 sky130_fd_sc_hd__a21o_2 _22806_ (.A1(_18851_),
    .A2(_18846_),
    .B1(_18853_),
    .X(_03251_));
 sky130_fd_sc_hd__buf_1 _22807_ (.A(\pcpi_mul.rs2[3] ),
    .X(_18854_));
 sky130_vsdinv _22808_ (.A(_18854_),
    .Y(_18855_));
 sky130_fd_sc_hd__buf_1 _22809_ (.A(_18855_),
    .X(_18856_));
 sky130_fd_sc_hd__buf_1 _22810_ (.A(_18856_),
    .X(_18857_));
 sky130_fd_sc_hd__buf_1 _22811_ (.A(_18857_),
    .X(_18858_));
 sky130_fd_sc_hd__buf_1 _22812_ (.A(_18858_),
    .X(_18859_));
 sky130_fd_sc_hd__buf_1 _22813_ (.A(_16956_),
    .X(_18860_));
 sky130_fd_sc_hd__buf_1 _22814_ (.A(_18860_),
    .X(_18861_));
 sky130_fd_sc_hd__buf_1 _22815_ (.A(_16964_),
    .X(_18862_));
 sky130_fd_sc_hd__buf_1 _22816_ (.A(_18862_),
    .X(_18863_));
 sky130_fd_sc_hd__nand2_2 _22817_ (.A(_18863_),
    .B(_18446_),
    .Y(_18864_));
 sky130_fd_sc_hd__o21ai_2 _22818_ (.A1(_18859_),
    .A2(_18861_),
    .B1(_18864_),
    .Y(_03250_));
 sky130_fd_sc_hd__buf_1 _22819_ (.A(\pcpi_mul.rs2[2] ),
    .X(_18865_));
 sky130_fd_sc_hd__buf_1 _22820_ (.A(_18865_),
    .X(_18866_));
 sky130_fd_sc_hd__buf_1 _22821_ (.A(_18866_),
    .X(_18867_));
 sky130_fd_sc_hd__buf_1 _22822_ (.A(_18867_),
    .X(_18868_));
 sky130_fd_sc_hd__buf_1 _22823_ (.A(_18868_),
    .X(_18869_));
 sky130_fd_sc_hd__and2_2 _22824_ (.A(_18836_),
    .B(_18448_),
    .X(_18870_));
 sky130_fd_sc_hd__a21o_2 _22825_ (.A1(_18869_),
    .A2(_18846_),
    .B1(_18870_),
    .X(_03249_));
 sky130_fd_sc_hd__buf_1 _22826_ (.A(\pcpi_mul.rs2[1] ),
    .X(_18871_));
 sky130_fd_sc_hd__buf_1 _22827_ (.A(_18871_),
    .X(_18872_));
 sky130_fd_sc_hd__buf_1 _22828_ (.A(_18872_),
    .X(_18873_));
 sky130_fd_sc_hd__buf_1 _22829_ (.A(_18873_),
    .X(_18874_));
 sky130_fd_sc_hd__buf_1 _22830_ (.A(_18874_),
    .X(_18875_));
 sky130_fd_sc_hd__and2_2 _22831_ (.A(_16965_),
    .B(_18451_),
    .X(_18876_));
 sky130_fd_sc_hd__a21o_2 _22832_ (.A1(_18875_),
    .A2(_18846_),
    .B1(_18876_),
    .X(_03248_));
 sky130_fd_sc_hd__buf_1 _22833_ (.A(\pcpi_mul.rs2[0] ),
    .X(_18877_));
 sky130_fd_sc_hd__buf_1 _22834_ (.A(_18877_),
    .X(_18878_));
 sky130_vsdinv _22835_ (.A(_18878_),
    .Y(_18879_));
 sky130_fd_sc_hd__buf_1 _22836_ (.A(_18879_),
    .X(_18880_));
 sky130_fd_sc_hd__buf_1 _22837_ (.A(_18880_),
    .X(_18881_));
 sky130_fd_sc_hd__nand2_2 _22838_ (.A(_18863_),
    .B(_18454_),
    .Y(_18882_));
 sky130_fd_sc_hd__o21ai_2 _22839_ (.A1(_18881_),
    .A2(_18861_),
    .B1(_18882_),
    .Y(_03247_));
 sky130_fd_sc_hd__mux2_2 _22840_ (.A0(mem_wstrb[3]),
    .A1(_02541_),
    .S(_16856_),
    .X(_03246_));
 sky130_fd_sc_hd__mux2_2 _22841_ (.A0(mem_wstrb[2]),
    .A1(_02540_),
    .S(_16856_),
    .X(_03245_));
 sky130_fd_sc_hd__mux2_2 _22842_ (.A0(mem_wstrb[1]),
    .A1(_02539_),
    .S(_16855_),
    .X(_03244_));
 sky130_fd_sc_hd__mux2_2 _22843_ (.A0(mem_wstrb[0]),
    .A1(_02538_),
    .S(_16855_),
    .X(_03243_));
 sky130_fd_sc_hd__and2_2 _22844_ (.A(_17230_),
    .B(_17229_),
    .X(_18883_));
 sky130_fd_sc_hd__and2b_2 _22845_ (.A_N(_00330_),
    .B(_16859_),
    .X(_18884_));
 sky130_fd_sc_hd__nor3b_2 _22846_ (.A(_17228_),
    .B(_16866_),
    .C_N(_18884_),
    .Y(_18885_));
 sky130_fd_sc_hd__buf_1 _22847_ (.A(_16872_),
    .X(_18886_));
 sky130_fd_sc_hd__o2bb2ai_2 _22848_ (.A1_N(_18883_),
    .A2_N(_18885_),
    .B1(_17279_),
    .B2(_18886_),
    .Y(_03242_));
 sky130_vsdinv _22849_ (.A(_17332_),
    .Y(_18887_));
 sky130_fd_sc_hd__and2b_2 _22850_ (.A_N(_17230_),
    .B(_17229_),
    .X(_18888_));
 sky130_fd_sc_hd__nand2_2 _22851_ (.A(_18885_),
    .B(_18888_),
    .Y(_18889_));
 sky130_fd_sc_hd__o21ai_2 _22852_ (.A1(_18887_),
    .A2(_19783_),
    .B1(_18889_),
    .Y(_03241_));
 sky130_fd_sc_hd__buf_1 _22853_ (.A(_18275_),
    .X(_18890_));
 sky130_fd_sc_hd__o2111ai_2 _22854_ (.A1(_18890_),
    .A2(_18547_),
    .B1(_18370_),
    .C1(_18549_),
    .D1(_18550_),
    .Y(_18891_));
 sky130_fd_sc_hd__buf_1 _22855_ (.A(_18891_),
    .X(_18892_));
 sky130_fd_sc_hd__buf_1 _22856_ (.A(_18892_),
    .X(_18893_));
 sky130_fd_sc_hd__mux2_2 _22857_ (.A0(_18650_),
    .A1(\cpuregs[13][31] ),
    .S(_18893_),
    .X(_03240_));
 sky130_fd_sc_hd__mux2_2 _22858_ (.A0(_18654_),
    .A1(\cpuregs[13][30] ),
    .S(_18893_),
    .X(_03239_));
 sky130_fd_sc_hd__mux2_2 _22859_ (.A0(_18655_),
    .A1(\cpuregs[13][29] ),
    .S(_18893_),
    .X(_03238_));
 sky130_fd_sc_hd__mux2_2 _22860_ (.A0(_18656_),
    .A1(\cpuregs[13][28] ),
    .S(_18893_),
    .X(_03237_));
 sky130_fd_sc_hd__buf_1 _22861_ (.A(_18892_),
    .X(_18894_));
 sky130_fd_sc_hd__mux2_2 _22862_ (.A0(_18657_),
    .A1(\cpuregs[13][27] ),
    .S(_18894_),
    .X(_03236_));
 sky130_fd_sc_hd__mux2_2 _22863_ (.A0(_18659_),
    .A1(\cpuregs[13][26] ),
    .S(_18894_),
    .X(_03235_));
 sky130_fd_sc_hd__mux2_2 _22864_ (.A0(_18660_),
    .A1(\cpuregs[13][25] ),
    .S(_18894_),
    .X(_03234_));
 sky130_fd_sc_hd__mux2_2 _22865_ (.A0(_18661_),
    .A1(\cpuregs[13][24] ),
    .S(_18894_),
    .X(_03233_));
 sky130_fd_sc_hd__buf_1 _22866_ (.A(_18892_),
    .X(_18895_));
 sky130_fd_sc_hd__mux2_2 _22867_ (.A0(_18662_),
    .A1(\cpuregs[13][23] ),
    .S(_18895_),
    .X(_03232_));
 sky130_fd_sc_hd__mux2_2 _22868_ (.A0(_18664_),
    .A1(\cpuregs[13][22] ),
    .S(_18895_),
    .X(_03231_));
 sky130_fd_sc_hd__mux2_2 _22869_ (.A0(_18665_),
    .A1(\cpuregs[13][21] ),
    .S(_18895_),
    .X(_03230_));
 sky130_fd_sc_hd__mux2_2 _22870_ (.A0(_18666_),
    .A1(\cpuregs[13][20] ),
    .S(_18895_),
    .X(_03229_));
 sky130_fd_sc_hd__buf_1 _22871_ (.A(_18892_),
    .X(_18896_));
 sky130_fd_sc_hd__mux2_2 _22872_ (.A0(_18667_),
    .A1(\cpuregs[13][19] ),
    .S(_18896_),
    .X(_03228_));
 sky130_fd_sc_hd__mux2_2 _22873_ (.A0(_18669_),
    .A1(\cpuregs[13][18] ),
    .S(_18896_),
    .X(_03227_));
 sky130_fd_sc_hd__mux2_2 _22874_ (.A0(_18670_),
    .A1(\cpuregs[13][17] ),
    .S(_18896_),
    .X(_03226_));
 sky130_fd_sc_hd__mux2_2 _22875_ (.A0(_18671_),
    .A1(\cpuregs[13][16] ),
    .S(_18896_),
    .X(_03225_));
 sky130_fd_sc_hd__buf_1 _22876_ (.A(_18891_),
    .X(_18897_));
 sky130_fd_sc_hd__buf_1 _22877_ (.A(_18897_),
    .X(_18898_));
 sky130_fd_sc_hd__mux2_2 _22878_ (.A0(_18672_),
    .A1(\cpuregs[13][15] ),
    .S(_18898_),
    .X(_03224_));
 sky130_fd_sc_hd__mux2_2 _22879_ (.A0(_18675_),
    .A1(\cpuregs[13][14] ),
    .S(_18898_),
    .X(_03223_));
 sky130_fd_sc_hd__mux2_2 _22880_ (.A0(_18676_),
    .A1(\cpuregs[13][13] ),
    .S(_18898_),
    .X(_03222_));
 sky130_fd_sc_hd__mux2_2 _22881_ (.A0(_18677_),
    .A1(\cpuregs[13][12] ),
    .S(_18898_),
    .X(_03221_));
 sky130_fd_sc_hd__buf_1 _22882_ (.A(_18897_),
    .X(_18899_));
 sky130_fd_sc_hd__mux2_2 _22883_ (.A0(_18678_),
    .A1(\cpuregs[13][11] ),
    .S(_18899_),
    .X(_03220_));
 sky130_fd_sc_hd__mux2_2 _22884_ (.A0(_18680_),
    .A1(\cpuregs[13][10] ),
    .S(_18899_),
    .X(_03219_));
 sky130_fd_sc_hd__mux2_2 _22885_ (.A0(_18681_),
    .A1(\cpuregs[13][9] ),
    .S(_18899_),
    .X(_03218_));
 sky130_fd_sc_hd__mux2_2 _22886_ (.A0(_18682_),
    .A1(\cpuregs[13][8] ),
    .S(_18899_),
    .X(_03217_));
 sky130_fd_sc_hd__buf_1 _22887_ (.A(_18897_),
    .X(_18900_));
 sky130_fd_sc_hd__mux2_2 _22888_ (.A0(_18683_),
    .A1(\cpuregs[13][7] ),
    .S(_18900_),
    .X(_03216_));
 sky130_fd_sc_hd__mux2_2 _22889_ (.A0(_18685_),
    .A1(\cpuregs[13][6] ),
    .S(_18900_),
    .X(_03215_));
 sky130_fd_sc_hd__mux2_2 _22890_ (.A0(_18686_),
    .A1(\cpuregs[13][5] ),
    .S(_18900_),
    .X(_03214_));
 sky130_fd_sc_hd__mux2_2 _22891_ (.A0(_18687_),
    .A1(\cpuregs[13][4] ),
    .S(_18900_),
    .X(_03213_));
 sky130_fd_sc_hd__buf_1 _22892_ (.A(_18897_),
    .X(_18901_));
 sky130_fd_sc_hd__mux2_2 _22893_ (.A0(_18688_),
    .A1(\cpuregs[13][3] ),
    .S(_18901_),
    .X(_03212_));
 sky130_fd_sc_hd__mux2_2 _22894_ (.A0(_18690_),
    .A1(\cpuregs[13][2] ),
    .S(_18901_),
    .X(_03211_));
 sky130_fd_sc_hd__mux2_2 _22895_ (.A0(_18691_),
    .A1(\cpuregs[13][1] ),
    .S(_18901_),
    .X(_03210_));
 sky130_fd_sc_hd__mux2_2 _22896_ (.A0(_18692_),
    .A1(\cpuregs[13][0] ),
    .S(_18901_),
    .X(_03209_));
 sky130_fd_sc_hd__and2b_2 _22897_ (.A_N(_17229_),
    .B(_17230_),
    .X(_18902_));
 sky130_fd_sc_hd__o2bb2ai_2 _22898_ (.A1_N(_18902_),
    .A2_N(_18885_),
    .B1(_17062_),
    .B2(_16863_),
    .Y(_03208_));
 sky130_fd_sc_hd__buf_1 _22899_ (.A(_17331_),
    .X(_18903_));
 sky130_fd_sc_hd__nor3b_2 _22900_ (.A(_17086_),
    .B(_17265_),
    .C_N(_17361_),
    .Y(_18904_));
 sky130_vsdinv _22901_ (.A(_17310_),
    .Y(_18905_));
 sky130_vsdinv _22902_ (.A(_17307_),
    .Y(_18906_));
 sky130_fd_sc_hd__a31o_2 _22903_ (.A1(_18905_),
    .A2(_18906_),
    .A3(_00335_),
    .B1(_18887_),
    .X(_18907_));
 sky130_fd_sc_hd__a2bb2oi_2 _22904_ (.A1_N(is_jalr_addi_slti_sltiu_xori_ori_andi),
    .A2_N(_18903_),
    .B1(_18904_),
    .B2(_18907_),
    .Y(_03207_));
 sky130_fd_sc_hd__buf_1 _22905_ (.A(is_slli_srli_srai),
    .X(_18908_));
 sky130_fd_sc_hd__buf_1 _22906_ (.A(_18908_),
    .X(_18909_));
 sky130_fd_sc_hd__buf_1 _22907_ (.A(_17341_),
    .X(_18910_));
 sky130_fd_sc_hd__buf_1 _22908_ (.A(_18910_),
    .X(_18911_));
 sky130_fd_sc_hd__buf_1 _22909_ (.A(_17243_),
    .X(_18912_));
 sky130_fd_sc_hd__buf_1 _22910_ (.A(_17305_),
    .X(_18913_));
 sky130_fd_sc_hd__or3b_2 _22911_ (.A(_18912_),
    .B(_17338_),
    .C_N(_18913_),
    .X(_18914_));
 sky130_fd_sc_hd__buf_1 _22912_ (.A(\mem_rdata_q[30] ),
    .X(_18915_));
 sky130_vsdinv _22913_ (.A(_17241_),
    .Y(_00334_));
 sky130_fd_sc_hd__buf_1 _22914_ (.A(\mem_rdata_q[31] ),
    .X(_18916_));
 sky130_fd_sc_hd__buf_1 _22915_ (.A(_18916_),
    .X(_18917_));
 sky130_fd_sc_hd__a2111o_2 _22916_ (.A1(_18915_),
    .A2(_00334_),
    .B1(_18917_),
    .C1(_17282_),
    .D1(_17254_),
    .X(_18918_));
 sky130_fd_sc_hd__o2bb2ai_2 _22917_ (.A1_N(_18909_),
    .A2_N(_18911_),
    .B1(_18914_),
    .B2(_18918_),
    .Y(_03206_));
 sky130_fd_sc_hd__o2bb2ai_2 _22918_ (.A1_N(_16867_),
    .A2_N(_18885_),
    .B1(_17059_),
    .B2(_16863_),
    .Y(_03205_));
 sky130_fd_sc_hd__buf_1 _22919_ (.A(\decoded_imm_uj[20] ),
    .X(_18919_));
 sky130_fd_sc_hd__buf_1 _22920_ (.A(_18919_),
    .X(_18920_));
 sky130_fd_sc_hd__buf_1 _22921_ (.A(_18920_),
    .X(_18921_));
 sky130_fd_sc_hd__buf_1 _22922_ (.A(_18921_),
    .X(_18922_));
 sky130_fd_sc_hd__buf_1 _22923_ (.A(_18922_),
    .X(_18923_));
 sky130_fd_sc_hd__buf_1 _22924_ (.A(_18923_),
    .X(_18924_));
 sky130_fd_sc_hd__buf_1 _22925_ (.A(_16862_),
    .X(_18925_));
 sky130_fd_sc_hd__mux2_2 _22926_ (.A0(_18924_),
    .A1(\mem_rdata_latched[31] ),
    .S(_18925_),
    .X(_03204_));
 sky130_fd_sc_hd__mux2_2 _22927_ (.A0(\decoded_imm_uj[19] ),
    .A1(\mem_rdata_latched[19] ),
    .S(_18925_),
    .X(_03203_));
 sky130_fd_sc_hd__buf_1 _22928_ (.A(\decoded_imm_uj[18] ),
    .X(_18926_));
 sky130_fd_sc_hd__buf_1 _22929_ (.A(_17237_),
    .X(_00337_));
 sky130_fd_sc_hd__a21o_2 _22930_ (.A1(_18926_),
    .A2(_00337_),
    .B1(_17235_),
    .X(_03202_));
 sky130_fd_sc_hd__a21o_2 _22931_ (.A1(\decoded_imm_uj[17] ),
    .A2(_00337_),
    .B1(_17238_),
    .X(_03201_));
 sky130_fd_sc_hd__a21o_2 _22932_ (.A1(\decoded_imm_uj[16] ),
    .A2(_00337_),
    .B1(_17239_),
    .X(_03200_));
 sky130_fd_sc_hd__a21o_2 _22933_ (.A1(\decoded_imm_uj[15] ),
    .A2(_17234_),
    .B1(_17240_),
    .X(_03199_));
 sky130_fd_sc_hd__mux2_2 _22934_ (.A0(\decoded_imm_uj[14] ),
    .A1(\mem_rdata_latched[14] ),
    .S(_18925_),
    .X(_03198_));
 sky130_fd_sc_hd__mux2_2 _22935_ (.A0(\decoded_imm_uj[13] ),
    .A1(\mem_rdata_latched[13] ),
    .S(_18925_),
    .X(_03197_));
 sky130_fd_sc_hd__buf_1 _22936_ (.A(_16859_),
    .X(_18927_));
 sky130_fd_sc_hd__buf_1 _22937_ (.A(_18927_),
    .X(_18928_));
 sky130_fd_sc_hd__mux2_2 _22938_ (.A0(\decoded_imm_uj[12] ),
    .A1(\mem_rdata_latched[12] ),
    .S(_18928_),
    .X(_03196_));
 sky130_fd_sc_hd__mux2_2 _22939_ (.A0(\decoded_imm_uj[11] ),
    .A1(\mem_rdata_latched[20] ),
    .S(_18928_),
    .X(_03195_));
 sky130_fd_sc_hd__buf_1 _22940_ (.A(\decoded_imm_uj[10] ),
    .X(_18929_));
 sky130_fd_sc_hd__mux2_2 _22941_ (.A0(_18929_),
    .A1(\mem_rdata_latched[30] ),
    .S(_18928_),
    .X(_03194_));
 sky130_fd_sc_hd__mux2_2 _22942_ (.A0(\decoded_imm_uj[9] ),
    .A1(\mem_rdata_latched[29] ),
    .S(_18928_),
    .X(_03193_));
 sky130_fd_sc_hd__buf_1 _22943_ (.A(\decoded_imm_uj[8] ),
    .X(_18930_));
 sky130_fd_sc_hd__buf_1 _22944_ (.A(_18927_),
    .X(_18931_));
 sky130_fd_sc_hd__mux2_2 _22945_ (.A0(_18930_),
    .A1(\mem_rdata_latched[28] ),
    .S(_18931_),
    .X(_03192_));
 sky130_fd_sc_hd__mux2_2 _22946_ (.A0(\decoded_imm_uj[7] ),
    .A1(\mem_rdata_latched[27] ),
    .S(_18931_),
    .X(_03191_));
 sky130_fd_sc_hd__mux2_2 _22947_ (.A0(\decoded_imm_uj[6] ),
    .A1(\mem_rdata_latched[26] ),
    .S(_18931_),
    .X(_03190_));
 sky130_fd_sc_hd__mux2_2 _22948_ (.A0(\decoded_imm_uj[5] ),
    .A1(\mem_rdata_latched[25] ),
    .S(_18931_),
    .X(_03189_));
 sky130_fd_sc_hd__buf_1 _22949_ (.A(\decoded_imm_uj[4] ),
    .X(_18932_));
 sky130_fd_sc_hd__buf_1 _22950_ (.A(_18927_),
    .X(_18933_));
 sky130_fd_sc_hd__mux2_2 _22951_ (.A0(_18932_),
    .A1(\mem_rdata_latched[24] ),
    .S(_18933_),
    .X(_03188_));
 sky130_fd_sc_hd__buf_1 _22952_ (.A(\decoded_imm_uj[3] ),
    .X(_18934_));
 sky130_fd_sc_hd__mux2_2 _22953_ (.A0(_18934_),
    .A1(\mem_rdata_latched[23] ),
    .S(_18933_),
    .X(_03187_));
 sky130_fd_sc_hd__mux2_2 _22954_ (.A0(\decoded_imm_uj[2] ),
    .A1(\mem_rdata_latched[22] ),
    .S(_18933_),
    .X(_03186_));
 sky130_fd_sc_hd__buf_1 _22955_ (.A(\decoded_imm_uj[1] ),
    .X(_18935_));
 sky130_fd_sc_hd__mux2_2 _22956_ (.A0(_18935_),
    .A1(\mem_rdata_latched[21] ),
    .S(_18933_),
    .X(_03185_));
 sky130_fd_sc_hd__buf_1 _22957_ (.A(is_sb_sh_sw),
    .X(_18936_));
 sky130_fd_sc_hd__buf_1 _22958_ (.A(\mem_rdata_q[7] ),
    .X(_18937_));
 sky130_vsdinv _22959_ (.A(\mem_rdata_q[20] ),
    .Y(_18938_));
 sky130_fd_sc_hd__nor3_2 _22960_ (.A(is_alu_reg_imm),
    .B(is_lb_lh_lw_lbu_lhu),
    .C(instr_jalr),
    .Y(_18939_));
 sky130_fd_sc_hd__o2bb2ai_2 _22961_ (.A1_N(_18936_),
    .A2_N(_18937_),
    .B1(_18938_),
    .B2(_18939_),
    .Y(_18940_));
 sky130_fd_sc_hd__buf_1 _22962_ (.A(\decoded_imm[0] ),
    .X(_18941_));
 sky130_fd_sc_hd__mux2_2 _22963_ (.A0(_18940_),
    .A1(_18941_),
    .S(_18910_),
    .X(_03184_));
 sky130_fd_sc_hd__buf_1 _22964_ (.A(_18927_),
    .X(_18942_));
 sky130_fd_sc_hd__mux2_2 _22965_ (.A0(\decoded_rd[4] ),
    .A1(\mem_rdata_latched[11] ),
    .S(_18942_),
    .X(_03183_));
 sky130_fd_sc_hd__mux2_2 _22966_ (.A0(\decoded_rd[3] ),
    .A1(\mem_rdata_latched[10] ),
    .S(_18942_),
    .X(_03182_));
 sky130_fd_sc_hd__mux2_2 _22967_ (.A0(\decoded_rd[2] ),
    .A1(\mem_rdata_latched[9] ),
    .S(_18942_),
    .X(_03181_));
 sky130_fd_sc_hd__mux2_2 _22968_ (.A0(\decoded_rd[1] ),
    .A1(\mem_rdata_latched[8] ),
    .S(_18942_),
    .X(_03180_));
 sky130_fd_sc_hd__mux2_2 _22969_ (.A0(\decoded_rd[0] ),
    .A1(\mem_rdata_latched[7] ),
    .S(_16872_),
    .X(_03179_));
 sky130_fd_sc_hd__nor3b_2 _22970_ (.A(\mem_rdata_q[4] ),
    .B(\mem_rdata_q[2] ),
    .C_N(\mem_rdata_q[3] ),
    .Y(_18943_));
 sky130_fd_sc_hd__nor2_2 _22971_ (.A(\mem_rdata_q[6] ),
    .B(\mem_rdata_q[5] ),
    .Y(_18944_));
 sky130_fd_sc_hd__and4_2 _22972_ (.A(_18943_),
    .B(\mem_rdata_q[1] ),
    .C(\mem_rdata_q[0] ),
    .D(_18944_),
    .X(_18945_));
 sky130_fd_sc_hd__buf_1 _22973_ (.A(\mem_rdata_q[25] ),
    .X(_18946_));
 sky130_vsdinv _22974_ (.A(_18946_),
    .Y(_18947_));
 sky130_fd_sc_hd__nor3b_2 _22975_ (.A(_18947_),
    .B(_17251_),
    .C_N(_17252_),
    .Y(_18948_));
 sky130_fd_sc_hd__buf_1 _22976_ (.A(\mem_rdata_q[27] ),
    .X(_18949_));
 sky130_fd_sc_hd__nand3b_2 _22977_ (.A_N(_17264_),
    .B(_18949_),
    .C(_17361_),
    .Y(_18950_));
 sky130_vsdinv _22978_ (.A(_18950_),
    .Y(_18951_));
 sky130_fd_sc_hd__buf_1 _22979_ (.A(_17022_),
    .X(_18952_));
 sky130_fd_sc_hd__buf_1 _22980_ (.A(_18952_),
    .X(_18953_));
 sky130_fd_sc_hd__buf_1 _22981_ (.A(_17258_),
    .X(_18954_));
 sky130_fd_sc_hd__buf_1 _22982_ (.A(_18954_),
    .X(_18955_));
 sky130_fd_sc_hd__a32o_2 _22983_ (.A1(_18945_),
    .A2(_18948_),
    .A3(_18951_),
    .B1(_18953_),
    .B2(_18955_),
    .X(_03178_));
 sky130_fd_sc_hd__buf_1 _22984_ (.A(_16879_),
    .X(_18956_));
 sky130_fd_sc_hd__nor2_2 _22985_ (.A(_16869_),
    .B(_16874_),
    .Y(_18957_));
 sky130_fd_sc_hd__nand3_2 _22986_ (.A(_18957_),
    .B(\mem_rdata_latched[27] ),
    .C(_16876_),
    .Y(_18958_));
 sky130_fd_sc_hd__o21ai_2 _22987_ (.A1(_18956_),
    .A2(_19783_),
    .B1(_18958_),
    .Y(_03177_));
 sky130_fd_sc_hd__buf_1 _22988_ (.A(\mem_rdata_q[28] ),
    .X(_18959_));
 sky130_fd_sc_hd__buf_1 _22989_ (.A(\mem_rdata_q[26] ),
    .X(_18960_));
 sky130_fd_sc_hd__nand3b_2 _22990_ (.A_N(_17283_),
    .B(_18960_),
    .C(_17337_),
    .Y(_18961_));
 sky130_fd_sc_hd__nor3_2 _22991_ (.A(_18959_),
    .B(_18949_),
    .C(_18961_),
    .Y(_18962_));
 sky130_fd_sc_hd__nor3b_2 _22992_ (.A(_18947_),
    .B(_17251_),
    .C_N(_18962_),
    .Y(_18963_));
 sky130_fd_sc_hd__o2bb2ai_2 _22993_ (.A1_N(_18945_),
    .A2_N(_18963_),
    .B1(_17006_),
    .B2(_18027_),
    .Y(_03176_));
 sky130_fd_sc_hd__o21ai_2 _22994_ (.A1(_17007_),
    .A2(_18886_),
    .B1(_16873_),
    .Y(_03175_));
 sky130_fd_sc_hd__nor3b_2 _22995_ (.A(\mem_rdata_q[27] ),
    .B(_17263_),
    .C_N(_17284_),
    .Y(_18964_));
 sky130_fd_sc_hd__a32o_2 _22996_ (.A1(_18945_),
    .A2(_18948_),
    .A3(_18964_),
    .B1(instr_setq),
    .B2(_18955_),
    .X(_03174_));
 sky130_fd_sc_hd__buf_1 _22997_ (.A(_17341_),
    .X(_18965_));
 sky130_fd_sc_hd__a22o_2 _22998_ (.A1(instr_getq),
    .A2(_18965_),
    .B1(_18945_),
    .B2(_17297_),
    .X(_03173_));
 sky130_fd_sc_hd__nor3_2 _22999_ (.A(\mem_rdata_q[17] ),
    .B(\mem_rdata_q[16] ),
    .C(\mem_rdata_q[15] ),
    .Y(_18966_));
 sky130_fd_sc_hd__or3b_2 _23000_ (.A(\mem_rdata_q[19] ),
    .B(\mem_rdata_q[18] ),
    .C_N(_18966_),
    .X(_18967_));
 sky130_fd_sc_hd__and4_2 _23001_ (.A(\mem_rdata_q[6] ),
    .B(\mem_rdata_q[5] ),
    .C(\mem_rdata_q[1] ),
    .D(\mem_rdata_q[0] ),
    .X(_18968_));
 sky130_fd_sc_hd__nor3b_2 _23002_ (.A(\mem_rdata_q[3] ),
    .B(\mem_rdata_q[2] ),
    .C_N(\mem_rdata_q[4] ),
    .Y(_18969_));
 sky130_fd_sc_hd__and2_2 _23003_ (.A(_18968_),
    .B(_18969_),
    .X(_18970_));
 sky130_fd_sc_hd__nand3b_2 _23004_ (.A_N(_18967_),
    .B(_17288_),
    .C(_18970_),
    .Y(_18971_));
 sky130_fd_sc_hd__buf_1 _23005_ (.A(_17258_),
    .X(_18972_));
 sky130_fd_sc_hd__or4_2 _23006_ (.A(\mem_rdata_q[11] ),
    .B(\mem_rdata_q[10] ),
    .C(\mem_rdata_q[8] ),
    .D(\mem_rdata_q[7] ),
    .X(_18973_));
 sky130_fd_sc_hd__or4_2 _23007_ (.A(\mem_rdata_q[24] ),
    .B(\mem_rdata_q[23] ),
    .C(\mem_rdata_q[22] ),
    .D(\mem_rdata_q[21] ),
    .X(_18974_));
 sky130_fd_sc_hd__or2_2 _23008_ (.A(_18973_),
    .B(_18974_),
    .X(_18975_));
 sky130_fd_sc_hd__or4_2 _23009_ (.A(\mem_rdata_q[9] ),
    .B(_18972_),
    .C(_17322_),
    .D(_18975_),
    .X(_18976_));
 sky130_fd_sc_hd__o2bb2ai_2 _23010_ (.A1_N(instr_ecall_ebreak),
    .A2_N(_18911_),
    .B1(_18971_),
    .B2(_18976_),
    .Y(_03172_));
 sky130_vsdinv _23011_ (.A(\mem_rdata_q[27] ),
    .Y(_18977_));
 sky130_fd_sc_hd__or4_2 _23012_ (.A(\mem_rdata_q[29] ),
    .B(\mem_rdata_q[28] ),
    .C(_17247_),
    .D(_17249_),
    .X(_18978_));
 sky130_fd_sc_hd__buf_1 _23013_ (.A(\mem_rdata_q[24] ),
    .X(_18979_));
 sky130_vsdinv _23014_ (.A(_18979_),
    .Y(_18980_));
 sky130_fd_sc_hd__nand3b_2 _23015_ (.A_N(_18978_),
    .B(_18947_),
    .C(_18980_),
    .Y(_18981_));
 sky130_fd_sc_hd__nor3_2 _23016_ (.A(_18977_),
    .B(_18960_),
    .C(_18981_),
    .Y(_18982_));
 sky130_fd_sc_hd__nor2_2 _23017_ (.A(_18905_),
    .B(_18967_),
    .Y(_18983_));
 sky130_fd_sc_hd__nor3b_2 _23018_ (.A(\mem_rdata_q[20] ),
    .B(_17283_),
    .C_N(_17284_),
    .Y(_18984_));
 sky130_fd_sc_hd__nor3b_2 _23019_ (.A(\mem_rdata_q[23] ),
    .B(\mem_rdata_q[22] ),
    .C_N(\mem_rdata_q[21] ),
    .Y(_18985_));
 sky130_fd_sc_hd__and4_2 _23020_ (.A(_18968_),
    .B(_18969_),
    .C(_18984_),
    .D(_18985_),
    .X(_18986_));
 sky130_fd_sc_hd__buf_1 _23021_ (.A(instr_rdinstrh),
    .X(_18987_));
 sky130_fd_sc_hd__buf_1 _23022_ (.A(_18987_),
    .X(_18988_));
 sky130_fd_sc_hd__buf_1 _23023_ (.A(_18954_),
    .X(_18989_));
 sky130_fd_sc_hd__a32o_2 _23024_ (.A1(_18982_),
    .A2(_18983_),
    .A3(_18986_),
    .B1(_18988_),
    .B2(_18989_),
    .X(_03171_));
 sky130_fd_sc_hd__buf_1 _23025_ (.A(instr_rdinstr),
    .X(_18990_));
 sky130_fd_sc_hd__buf_1 _23026_ (.A(_18990_),
    .X(_18991_));
 sky130_vsdinv _23027_ (.A(_18983_),
    .Y(_18992_));
 sky130_vsdinv _23028_ (.A(\mem_rdata_q[26] ),
    .Y(_18993_));
 sky130_fd_sc_hd__and4_2 _23029_ (.A(_18964_),
    .B(_18985_),
    .C(_18993_),
    .D(_18938_),
    .X(_18994_));
 sky130_fd_sc_hd__nand3b_2 _23030_ (.A_N(_18981_),
    .B(_18970_),
    .C(_18994_),
    .Y(_18995_));
 sky130_fd_sc_hd__o2bb2ai_2 _23031_ (.A1_N(_18991_),
    .A2_N(_18911_),
    .B1(_18992_),
    .B2(_18995_),
    .Y(_03170_));
 sky130_fd_sc_hd__buf_1 _23032_ (.A(instr_rdcycleh),
    .X(_18996_));
 sky130_fd_sc_hd__buf_1 _23033_ (.A(_18996_),
    .X(_18997_));
 sky130_vsdinv _23034_ (.A(_18970_),
    .Y(_18998_));
 sky130_fd_sc_hd__or4_2 _23035_ (.A(\mem_rdata_q[23] ),
    .B(\mem_rdata_q[22] ),
    .C(\mem_rdata_q[21] ),
    .D(_17257_),
    .X(_18999_));
 sky130_fd_sc_hd__nor2_2 _23036_ (.A(_18998_),
    .B(_18999_),
    .Y(_19000_));
 sky130_fd_sc_hd__nand2_2 _23037_ (.A(_18982_),
    .B(_19000_),
    .Y(_19001_));
 sky130_fd_sc_hd__o2bb2ai_2 _23038_ (.A1_N(_18997_),
    .A2_N(_18911_),
    .B1(_18992_),
    .B2(_19001_),
    .Y(_03169_));
 sky130_fd_sc_hd__buf_1 _23039_ (.A(_18910_),
    .X(_19002_));
 sky130_fd_sc_hd__nand3_2 _23040_ (.A(_17253_),
    .B(_18993_),
    .C(_18980_),
    .Y(_19003_));
 sky130_fd_sc_hd__nor3_2 _23041_ (.A(_19003_),
    .B(_18978_),
    .C(_18998_),
    .Y(_19004_));
 sky130_fd_sc_hd__or2b_2 _23042_ (.A(_18999_),
    .B_N(_19004_),
    .X(_19005_));
 sky130_fd_sc_hd__o2bb2ai_2 _23043_ (.A1_N(instr_rdcycle),
    .A2_N(_19002_),
    .B1(_18992_),
    .B2(_19005_),
    .Y(_03168_));
 sky130_fd_sc_hd__nor2_2 _23044_ (.A(_18887_),
    .B(_17280_),
    .Y(_19006_));
 sky130_fd_sc_hd__a32o_2 _23045_ (.A1(_17278_),
    .A2(_17285_),
    .A3(_19006_),
    .B1(instr_srai),
    .B2(_18989_),
    .X(_03167_));
 sky130_fd_sc_hd__buf_1 _23046_ (.A(_17330_),
    .X(_19007_));
 sky130_fd_sc_hd__nand3_2 _23047_ (.A(_17288_),
    .B(_19007_),
    .C(_19006_),
    .Y(_19008_));
 sky130_fd_sc_hd__o21ai_2 _23048_ (.A1(_16992_),
    .A2(_18903_),
    .B1(_19008_),
    .Y(_03166_));
 sky130_fd_sc_hd__buf_1 _23049_ (.A(instr_slli),
    .X(_19009_));
 sky130_fd_sc_hd__a32o_2 _23050_ (.A1(_17297_),
    .A2(_17344_),
    .A3(_17367_),
    .B1(_19009_),
    .B2(_18989_),
    .X(_03165_));
 sky130_fd_sc_hd__nand3b_2 _23051_ (.A_N(_17264_),
    .B(_18936_),
    .C(_17810_),
    .Y(_19010_));
 sky130_fd_sc_hd__o2bb2ai_2 _23052_ (.A1_N(instr_sw),
    .A2_N(_19002_),
    .B1(_19010_),
    .B2(_18905_),
    .Y(_03164_));
 sky130_vsdinv _23053_ (.A(instr_sh),
    .Y(_19011_));
 sky130_fd_sc_hd__nand3_2 _23054_ (.A(_17367_),
    .B(_18936_),
    .C(_19007_),
    .Y(_19012_));
 sky130_fd_sc_hd__o21ai_2 _23055_ (.A1(_19011_),
    .A2(_18903_),
    .B1(_19012_),
    .Y(_03163_));
 sky130_vsdinv _23056_ (.A(instr_sb),
    .Y(_19013_));
 sky130_fd_sc_hd__buf_1 _23057_ (.A(_18026_),
    .X(_19014_));
 sky130_fd_sc_hd__o22ai_2 _23058_ (.A1(_19013_),
    .A2(_19014_),
    .B1(_19010_),
    .B2(_17357_),
    .Y(_03162_));
 sky130_fd_sc_hd__nand3b_2 _23059_ (.A_N(_17283_),
    .B(is_lb_lh_lw_lbu_lhu),
    .C(_17337_),
    .Y(_19015_));
 sky130_fd_sc_hd__o2bb2ai_2 _23060_ (.A1_N(instr_lhu),
    .A2_N(_19002_),
    .B1(_17280_),
    .B2(_19015_),
    .Y(_03161_));
 sky130_vsdinv _23061_ (.A(_19015_),
    .Y(_19016_));
 sky130_fd_sc_hd__a22o_2 _23062_ (.A1(_19016_),
    .A2(_17299_),
    .B1(instr_lbu),
    .B2(_18965_),
    .X(_03160_));
 sky130_fd_sc_hd__o2bb2ai_2 _23063_ (.A1_N(instr_lw),
    .A2_N(_19002_),
    .B1(_19015_),
    .B2(_18905_),
    .Y(_03159_));
 sky130_fd_sc_hd__o2bb2ai_2 _23064_ (.A1_N(_17367_),
    .A2_N(_19016_),
    .B1(_16826_),
    .B2(_18027_),
    .Y(_03158_));
 sky130_fd_sc_hd__o22ai_2 _23065_ (.A1(_16820_),
    .A2(_19014_),
    .B1(_19015_),
    .B2(_17357_),
    .Y(_03157_));
 sky130_fd_sc_hd__inv_2 _23066_ (.A(_17086_),
    .Y(_02063_));
 sky130_fd_sc_hd__nand3_2 _23067_ (.A(_00325_),
    .B(_00324_),
    .C(_00326_),
    .Y(_19017_));
 sky130_fd_sc_hd__nor2_2 _23068_ (.A(_17228_),
    .B(_19017_),
    .Y(_19018_));
 sky130_fd_sc_hd__nor3_2 _23069_ (.A(\mem_rdata_latched[14] ),
    .B(\mem_rdata_latched[13] ),
    .C(\mem_rdata_latched[12] ),
    .Y(_19019_));
 sky130_fd_sc_hd__and3b_2 _23070_ (.A_N(_17231_),
    .B(_19018_),
    .C(_19019_),
    .X(_19020_));
 sky130_fd_sc_hd__nand2_2 _23071_ (.A(_16876_),
    .B(_19020_),
    .Y(_19021_));
 sky130_fd_sc_hd__o21ai_2 _23072_ (.A1(_02063_),
    .A2(_18886_),
    .B1(_19021_),
    .Y(_03156_));
 sky130_fd_sc_hd__buf_1 _23073_ (.A(_16989_),
    .X(_00323_));
 sky130_fd_sc_hd__nor3b_2 _23074_ (.A(_19017_),
    .B(_17231_),
    .C_N(_17228_),
    .Y(_19022_));
 sky130_fd_sc_hd__nand2_2 _23075_ (.A(_16876_),
    .B(_19022_),
    .Y(_19023_));
 sky130_fd_sc_hd__o21ai_2 _23076_ (.A1(_00323_),
    .A2(_18886_),
    .B1(_19023_),
    .Y(_03155_));
 sky130_fd_sc_hd__a32o_2 _23077_ (.A1(_18884_),
    .A2(_18888_),
    .A3(_19018_),
    .B1(instr_auipc),
    .B2(_17234_),
    .X(_03154_));
 sky130_fd_sc_hd__buf_1 _23078_ (.A(instr_lui),
    .X(_19024_));
 sky130_fd_sc_hd__a32o_2 _23079_ (.A1(_18884_),
    .A2(_18883_),
    .A3(_19018_),
    .B1(_19024_),
    .B2(_17234_),
    .X(_03153_));
 sky130_fd_sc_hd__mux2_2 _23080_ (.A0(pcpi_insn[31]),
    .A1(_18917_),
    .S(_19007_),
    .X(_03152_));
 sky130_fd_sc_hd__mux2_2 _23081_ (.A0(pcpi_insn[30]),
    .A1(_18915_),
    .S(_19007_),
    .X(_03151_));
 sky130_fd_sc_hd__buf_1 _23082_ (.A(_18026_),
    .X(_19025_));
 sky130_fd_sc_hd__o21ba_2 _23083_ (.A1(pcpi_insn[29]),
    .A2(_19025_),
    .B1_N(_17285_),
    .X(_03150_));
 sky130_fd_sc_hd__buf_1 _23084_ (.A(_17256_),
    .X(_19026_));
 sky130_fd_sc_hd__buf_1 _23085_ (.A(_19026_),
    .X(_19027_));
 sky130_fd_sc_hd__mux2_2 _23086_ (.A0(pcpi_insn[28]),
    .A1(_18959_),
    .S(_19027_),
    .X(_03149_));
 sky130_fd_sc_hd__o21ba_2 _23087_ (.A1(pcpi_insn[27]),
    .A2(_19014_),
    .B1_N(_18964_),
    .X(_03148_));
 sky130_fd_sc_hd__a21bo_2 _23088_ (.A1(_18955_),
    .A2(pcpi_insn[26]),
    .B1_N(_18961_),
    .X(_03147_));
 sky130_fd_sc_hd__mux2_2 _23089_ (.A0(pcpi_insn[25]),
    .A1(_18946_),
    .S(_19027_),
    .X(_03146_));
 sky130_fd_sc_hd__mux2_2 _23090_ (.A0(pcpi_insn[24]),
    .A1(_18979_),
    .S(_19027_),
    .X(_03145_));
 sky130_fd_sc_hd__buf_1 _23091_ (.A(\mem_rdata_q[23] ),
    .X(_19028_));
 sky130_fd_sc_hd__mux2_2 _23092_ (.A0(pcpi_insn[23]),
    .A1(_19028_),
    .S(_19027_),
    .X(_03144_));
 sky130_fd_sc_hd__buf_1 _23093_ (.A(\mem_rdata_q[22] ),
    .X(_19029_));
 sky130_fd_sc_hd__buf_1 _23094_ (.A(_17289_),
    .X(_19030_));
 sky130_fd_sc_hd__buf_1 _23095_ (.A(_19030_),
    .X(_19031_));
 sky130_fd_sc_hd__mux2_2 _23096_ (.A0(pcpi_insn[22]),
    .A1(_19029_),
    .S(_19031_),
    .X(_03143_));
 sky130_fd_sc_hd__buf_1 _23097_ (.A(\mem_rdata_q[21] ),
    .X(_19032_));
 sky130_fd_sc_hd__mux2_2 _23098_ (.A0(pcpi_insn[21]),
    .A1(_19032_),
    .S(_19031_),
    .X(_03142_));
 sky130_fd_sc_hd__o21ba_2 _23099_ (.A1(pcpi_insn[20]),
    .A2(_19014_),
    .B1_N(_18984_),
    .X(_03141_));
 sky130_fd_sc_hd__mux2_2 _23100_ (.A0(pcpi_insn[19]),
    .A1(\mem_rdata_q[19] ),
    .S(_19031_),
    .X(_03140_));
 sky130_fd_sc_hd__mux2_2 _23101_ (.A0(pcpi_insn[18]),
    .A1(\mem_rdata_q[18] ),
    .S(_19031_),
    .X(_03139_));
 sky130_fd_sc_hd__buf_1 _23102_ (.A(_19030_),
    .X(_19033_));
 sky130_fd_sc_hd__mux2_2 _23103_ (.A0(pcpi_insn[17]),
    .A1(\mem_rdata_q[17] ),
    .S(_19033_),
    .X(_03138_));
 sky130_fd_sc_hd__mux2_2 _23104_ (.A0(pcpi_insn[16]),
    .A1(\mem_rdata_q[16] ),
    .S(_19033_),
    .X(_03137_));
 sky130_fd_sc_hd__mux2_2 _23105_ (.A0(pcpi_insn[15]),
    .A1(\mem_rdata_q[15] ),
    .S(_19033_),
    .X(_03136_));
 sky130_fd_sc_hd__mux2_2 _23106_ (.A0(pcpi_insn[14]),
    .A1(_17242_),
    .S(_19033_),
    .X(_03135_));
 sky130_fd_sc_hd__buf_1 _23107_ (.A(_19030_),
    .X(_19034_));
 sky130_fd_sc_hd__mux2_2 _23108_ (.A0(_16938_),
    .A1(_18912_),
    .S(_19034_),
    .X(_03134_));
 sky130_fd_sc_hd__mux2_2 _23109_ (.A0(pcpi_insn[12]),
    .A1(_18913_),
    .S(_19034_),
    .X(_03133_));
 sky130_fd_sc_hd__mux2_2 _23110_ (.A0(pcpi_insn[11]),
    .A1(\mem_rdata_q[11] ),
    .S(_19034_),
    .X(_03132_));
 sky130_fd_sc_hd__mux2_2 _23111_ (.A0(pcpi_insn[10]),
    .A1(\mem_rdata_q[10] ),
    .S(_19034_),
    .X(_03131_));
 sky130_fd_sc_hd__buf_1 _23112_ (.A(_19030_),
    .X(_19035_));
 sky130_fd_sc_hd__mux2_2 _23113_ (.A0(pcpi_insn[9]),
    .A1(\mem_rdata_q[9] ),
    .S(_19035_),
    .X(_03130_));
 sky130_fd_sc_hd__mux2_2 _23114_ (.A0(pcpi_insn[8]),
    .A1(\mem_rdata_q[8] ),
    .S(_19035_),
    .X(_03129_));
 sky130_fd_sc_hd__mux2_2 _23115_ (.A0(pcpi_insn[7]),
    .A1(_18937_),
    .S(_19035_),
    .X(_03128_));
 sky130_fd_sc_hd__mux2_2 _23116_ (.A0(pcpi_insn[6]),
    .A1(\mem_rdata_q[6] ),
    .S(_19035_),
    .X(_03127_));
 sky130_fd_sc_hd__buf_1 _23117_ (.A(_17330_),
    .X(_19036_));
 sky130_fd_sc_hd__mux2_2 _23118_ (.A0(pcpi_insn[5]),
    .A1(\mem_rdata_q[5] ),
    .S(_19036_),
    .X(_03126_));
 sky130_fd_sc_hd__mux2_2 _23119_ (.A0(pcpi_insn[4]),
    .A1(\mem_rdata_q[4] ),
    .S(_19036_),
    .X(_03125_));
 sky130_fd_sc_hd__mux2_2 _23120_ (.A0(pcpi_insn[3]),
    .A1(\mem_rdata_q[3] ),
    .S(_19036_),
    .X(_03124_));
 sky130_fd_sc_hd__mux2_2 _23121_ (.A0(pcpi_insn[2]),
    .A1(\mem_rdata_q[2] ),
    .S(_19036_),
    .X(_03123_));
 sky130_fd_sc_hd__mux2_2 _23122_ (.A0(pcpi_insn[1]),
    .A1(\mem_rdata_q[1] ),
    .S(_17345_),
    .X(_03122_));
 sky130_fd_sc_hd__mux2_2 _23123_ (.A0(pcpi_insn[0]),
    .A1(\mem_rdata_q[0] ),
    .S(_17345_),
    .X(_03121_));
 sky130_fd_sc_hd__nor2_2 _23124_ (.A(\cpu_state[2] ),
    .B(\cpu_state[6] ),
    .Y(_19037_));
 sky130_fd_sc_hd__a2111o_2 _23125_ (.A1(_19037_),
    .A2(_18029_),
    .B1(_16930_),
    .C1(_00318_),
    .D1(_00320_),
    .X(_19038_));
 sky130_fd_sc_hd__buf_1 _23126_ (.A(_19038_),
    .X(_19039_));
 sky130_fd_sc_hd__buf_1 _23127_ (.A(_19039_),
    .X(_19040_));
 sky130_fd_sc_hd__mux2_2 _23128_ (.A0(_02499_),
    .A1(_16958_),
    .S(_19040_),
    .X(_03120_));
 sky130_fd_sc_hd__buf_1 _23129_ (.A(pcpi_rs1[30]),
    .X(_19041_));
 sky130_fd_sc_hd__buf_1 _23130_ (.A(_19041_),
    .X(_19042_));
 sky130_fd_sc_hd__mux2_2 _23131_ (.A0(_02498_),
    .A1(_19042_),
    .S(_19040_),
    .X(_03119_));
 sky130_fd_sc_hd__buf_1 _23132_ (.A(pcpi_rs1[29]),
    .X(_19043_));
 sky130_fd_sc_hd__buf_1 _23133_ (.A(_19043_),
    .X(_19044_));
 sky130_fd_sc_hd__mux2_2 _23134_ (.A0(_02496_),
    .A1(_19044_),
    .S(_19040_),
    .X(_03118_));
 sky130_fd_sc_hd__buf_1 _23135_ (.A(pcpi_rs1[28]),
    .X(_19045_));
 sky130_fd_sc_hd__buf_1 _23136_ (.A(_19045_),
    .X(_19046_));
 sky130_fd_sc_hd__mux2_2 _23137_ (.A0(_02495_),
    .A1(_19046_),
    .S(_19040_),
    .X(_03117_));
 sky130_fd_sc_hd__buf_1 _23138_ (.A(pcpi_rs1[27]),
    .X(_19047_));
 sky130_fd_sc_hd__buf_1 _23139_ (.A(_19047_),
    .X(_19048_));
 sky130_fd_sc_hd__buf_1 _23140_ (.A(_19039_),
    .X(_19049_));
 sky130_fd_sc_hd__mux2_2 _23141_ (.A0(_02494_),
    .A1(_19048_),
    .S(_19049_),
    .X(_03116_));
 sky130_fd_sc_hd__buf_1 _23142_ (.A(pcpi_rs1[26]),
    .X(_19050_));
 sky130_fd_sc_hd__buf_1 _23143_ (.A(_19050_),
    .X(_19051_));
 sky130_fd_sc_hd__mux2_2 _23144_ (.A0(_02493_),
    .A1(_19051_),
    .S(_19049_),
    .X(_03115_));
 sky130_fd_sc_hd__buf_1 _23145_ (.A(pcpi_rs1[25]),
    .X(_19052_));
 sky130_fd_sc_hd__buf_1 _23146_ (.A(_19052_),
    .X(_19053_));
 sky130_fd_sc_hd__mux2_2 _23147_ (.A0(_02492_),
    .A1(_19053_),
    .S(_19049_),
    .X(_03114_));
 sky130_fd_sc_hd__buf_1 _23148_ (.A(pcpi_rs1[24]),
    .X(_19054_));
 sky130_fd_sc_hd__buf_1 _23149_ (.A(_19054_),
    .X(_19055_));
 sky130_fd_sc_hd__mux2_2 _23150_ (.A0(_02491_),
    .A1(_19055_),
    .S(_19049_),
    .X(_03113_));
 sky130_fd_sc_hd__buf_1 _23151_ (.A(pcpi_rs1[23]),
    .X(_19056_));
 sky130_fd_sc_hd__buf_1 _23152_ (.A(_19056_),
    .X(_19057_));
 sky130_fd_sc_hd__buf_1 _23153_ (.A(_19039_),
    .X(_19058_));
 sky130_fd_sc_hd__mux2_2 _23154_ (.A0(_02490_),
    .A1(_19057_),
    .S(_19058_),
    .X(_03112_));
 sky130_fd_sc_hd__buf_1 _23155_ (.A(pcpi_rs1[22]),
    .X(_19059_));
 sky130_fd_sc_hd__buf_1 _23156_ (.A(_19059_),
    .X(_19060_));
 sky130_fd_sc_hd__mux2_2 _23157_ (.A0(_02489_),
    .A1(_19060_),
    .S(_19058_),
    .X(_03111_));
 sky130_fd_sc_hd__buf_1 _23158_ (.A(pcpi_rs1[21]),
    .X(_19061_));
 sky130_fd_sc_hd__buf_1 _23159_ (.A(_19061_),
    .X(_19062_));
 sky130_fd_sc_hd__mux2_2 _23160_ (.A0(_02488_),
    .A1(_19062_),
    .S(_19058_),
    .X(_03110_));
 sky130_fd_sc_hd__buf_1 _23161_ (.A(pcpi_rs1[20]),
    .X(_19063_));
 sky130_fd_sc_hd__buf_1 _23162_ (.A(_19063_),
    .X(_19064_));
 sky130_fd_sc_hd__mux2_2 _23163_ (.A0(_02487_),
    .A1(_19064_),
    .S(_19058_),
    .X(_03109_));
 sky130_fd_sc_hd__buf_1 _23164_ (.A(pcpi_rs1[19]),
    .X(_19065_));
 sky130_fd_sc_hd__buf_1 _23165_ (.A(_19065_),
    .X(_19066_));
 sky130_fd_sc_hd__buf_1 _23166_ (.A(_19039_),
    .X(_19067_));
 sky130_fd_sc_hd__mux2_2 _23167_ (.A0(_02485_),
    .A1(_19066_),
    .S(_19067_),
    .X(_03108_));
 sky130_fd_sc_hd__buf_1 _23168_ (.A(pcpi_rs1[18]),
    .X(_19068_));
 sky130_fd_sc_hd__buf_1 _23169_ (.A(_19068_),
    .X(_19069_));
 sky130_fd_sc_hd__mux2_2 _23170_ (.A0(_02484_),
    .A1(_19069_),
    .S(_19067_),
    .X(_03107_));
 sky130_fd_sc_hd__buf_1 _23171_ (.A(pcpi_rs1[17]),
    .X(_19070_));
 sky130_fd_sc_hd__buf_1 _23172_ (.A(_19070_),
    .X(_19071_));
 sky130_fd_sc_hd__buf_1 _23173_ (.A(_19071_),
    .X(_19072_));
 sky130_fd_sc_hd__mux2_2 _23174_ (.A0(_02483_),
    .A1(_19072_),
    .S(_19067_),
    .X(_03106_));
 sky130_fd_sc_hd__buf_1 _23175_ (.A(pcpi_rs1[16]),
    .X(_19073_));
 sky130_fd_sc_hd__buf_1 _23176_ (.A(_19073_),
    .X(_19074_));
 sky130_fd_sc_hd__buf_1 _23177_ (.A(_19074_),
    .X(_19075_));
 sky130_fd_sc_hd__mux2_2 _23178_ (.A0(_02482_),
    .A1(_19075_),
    .S(_19067_),
    .X(_03105_));
 sky130_fd_sc_hd__buf_1 _23179_ (.A(pcpi_rs1[15]),
    .X(_19076_));
 sky130_fd_sc_hd__buf_1 _23180_ (.A(_19076_),
    .X(_19077_));
 sky130_fd_sc_hd__buf_1 _23181_ (.A(_19038_),
    .X(_19078_));
 sky130_fd_sc_hd__buf_1 _23182_ (.A(_19078_),
    .X(_19079_));
 sky130_fd_sc_hd__mux2_2 _23183_ (.A0(_02481_),
    .A1(_19077_),
    .S(_19079_),
    .X(_03104_));
 sky130_fd_sc_hd__buf_1 _23184_ (.A(pcpi_rs1[14]),
    .X(_19080_));
 sky130_fd_sc_hd__buf_1 _23185_ (.A(_19080_),
    .X(_19081_));
 sky130_fd_sc_hd__mux2_2 _23186_ (.A0(_02480_),
    .A1(_19081_),
    .S(_19079_),
    .X(_03103_));
 sky130_fd_sc_hd__buf_1 _23187_ (.A(pcpi_rs1[13]),
    .X(_19082_));
 sky130_fd_sc_hd__buf_1 _23188_ (.A(_19082_),
    .X(_19083_));
 sky130_fd_sc_hd__mux2_2 _23189_ (.A0(_02479_),
    .A1(_19083_),
    .S(_19079_),
    .X(_03102_));
 sky130_fd_sc_hd__buf_1 _23190_ (.A(pcpi_rs1[12]),
    .X(_19084_));
 sky130_fd_sc_hd__buf_1 _23191_ (.A(_19084_),
    .X(_19085_));
 sky130_fd_sc_hd__mux2_2 _23192_ (.A0(_02478_),
    .A1(_19085_),
    .S(_19079_),
    .X(_03101_));
 sky130_fd_sc_hd__buf_1 _23193_ (.A(pcpi_rs1[11]),
    .X(_19086_));
 sky130_fd_sc_hd__buf_1 _23194_ (.A(_19086_),
    .X(_19087_));
 sky130_fd_sc_hd__buf_1 _23195_ (.A(_19078_),
    .X(_19088_));
 sky130_fd_sc_hd__mux2_2 _23196_ (.A0(_02477_),
    .A1(_19087_),
    .S(_19088_),
    .X(_03100_));
 sky130_fd_sc_hd__buf_1 _23197_ (.A(pcpi_rs1[10]),
    .X(_19089_));
 sky130_fd_sc_hd__buf_1 _23198_ (.A(_19089_),
    .X(_19090_));
 sky130_fd_sc_hd__mux2_2 _23199_ (.A0(_02476_),
    .A1(_19090_),
    .S(_19088_),
    .X(_03099_));
 sky130_fd_sc_hd__buf_1 _23200_ (.A(pcpi_rs1[9]),
    .X(_19091_));
 sky130_fd_sc_hd__buf_1 _23201_ (.A(_19091_),
    .X(_19092_));
 sky130_fd_sc_hd__buf_1 _23202_ (.A(_19092_),
    .X(_19093_));
 sky130_fd_sc_hd__mux2_2 _23203_ (.A0(_02506_),
    .A1(_19093_),
    .S(_19088_),
    .X(_03098_));
 sky130_fd_sc_hd__buf_1 _23204_ (.A(pcpi_rs1[8]),
    .X(_19094_));
 sky130_fd_sc_hd__buf_1 _23205_ (.A(_19094_),
    .X(_19095_));
 sky130_fd_sc_hd__buf_1 _23206_ (.A(_19095_),
    .X(_19096_));
 sky130_fd_sc_hd__mux2_2 _23207_ (.A0(_02505_),
    .A1(_19096_),
    .S(_19088_),
    .X(_03097_));
 sky130_fd_sc_hd__buf_1 _23208_ (.A(pcpi_rs1[7]),
    .X(_19097_));
 sky130_fd_sc_hd__buf_1 _23209_ (.A(_19097_),
    .X(_19098_));
 sky130_fd_sc_hd__buf_1 _23210_ (.A(_19098_),
    .X(_19099_));
 sky130_fd_sc_hd__buf_1 _23211_ (.A(_19078_),
    .X(_19100_));
 sky130_fd_sc_hd__mux2_2 _23212_ (.A0(_02504_),
    .A1(_19099_),
    .S(_19100_),
    .X(_03096_));
 sky130_fd_sc_hd__buf_1 _23213_ (.A(pcpi_rs1[6]),
    .X(_19101_));
 sky130_fd_sc_hd__buf_1 _23214_ (.A(_19101_),
    .X(_19102_));
 sky130_fd_sc_hd__buf_1 _23215_ (.A(_19102_),
    .X(_19103_));
 sky130_fd_sc_hd__mux2_2 _23216_ (.A0(_02503_),
    .A1(_19103_),
    .S(_19100_),
    .X(_03095_));
 sky130_fd_sc_hd__buf_1 _23217_ (.A(pcpi_rs1[5]),
    .X(_19104_));
 sky130_fd_sc_hd__buf_1 _23218_ (.A(_19104_),
    .X(_19105_));
 sky130_fd_sc_hd__mux2_2 _23219_ (.A0(_02502_),
    .A1(_19105_),
    .S(_19100_),
    .X(_03094_));
 sky130_fd_sc_hd__buf_1 _23220_ (.A(pcpi_rs1[4]),
    .X(_19106_));
 sky130_fd_sc_hd__buf_1 _23221_ (.A(_19106_),
    .X(_19107_));
 sky130_fd_sc_hd__buf_1 _23222_ (.A(_19107_),
    .X(_19108_));
 sky130_fd_sc_hd__mux2_2 _23223_ (.A0(_02501_),
    .A1(_19108_),
    .S(_19100_),
    .X(_03093_));
 sky130_fd_sc_hd__buf_1 _23224_ (.A(pcpi_rs1[3]),
    .X(_19109_));
 sky130_fd_sc_hd__buf_1 _23225_ (.A(_19109_),
    .X(_19110_));
 sky130_fd_sc_hd__buf_1 _23226_ (.A(_19078_),
    .X(_19111_));
 sky130_fd_sc_hd__mux2_2 _23227_ (.A0(_02500_),
    .A1(_19110_),
    .S(_19111_),
    .X(_03092_));
 sky130_fd_sc_hd__buf_1 _23228_ (.A(pcpi_rs1[2]),
    .X(_19112_));
 sky130_fd_sc_hd__buf_1 _23229_ (.A(_19112_),
    .X(_19113_));
 sky130_fd_sc_hd__mux2_2 _23230_ (.A0(_02497_),
    .A1(_19113_),
    .S(_19111_),
    .X(_03091_));
 sky130_fd_sc_hd__buf_1 _23231_ (.A(pcpi_rs1[1]),
    .X(_19114_));
 sky130_fd_sc_hd__buf_1 _23232_ (.A(_19114_),
    .X(_19115_));
 sky130_fd_sc_hd__buf_1 _23233_ (.A(_19115_),
    .X(_19116_));
 sky130_fd_sc_hd__buf_1 _23234_ (.A(_19116_),
    .X(_19117_));
 sky130_fd_sc_hd__buf_1 _23235_ (.A(_19117_),
    .X(_19118_));
 sky130_fd_sc_hd__mux2_2 _23236_ (.A0(_02486_),
    .A1(_19118_),
    .S(_19111_),
    .X(_03090_));
 sky130_fd_sc_hd__buf_1 _23237_ (.A(pcpi_rs1[0]),
    .X(_19119_));
 sky130_fd_sc_hd__buf_1 _23238_ (.A(_19119_),
    .X(_19120_));
 sky130_fd_sc_hd__buf_1 _23239_ (.A(_19120_),
    .X(_19121_));
 sky130_fd_sc_hd__buf_1 _23240_ (.A(_19121_),
    .X(_19122_));
 sky130_fd_sc_hd__buf_1 _23241_ (.A(_19122_),
    .X(_19123_));
 sky130_fd_sc_hd__buf_1 _23242_ (.A(_19123_),
    .X(_19124_));
 sky130_fd_sc_hd__mux2_2 _23243_ (.A0(_02475_),
    .A1(_19124_),
    .S(_19111_),
    .X(_03089_));
 sky130_fd_sc_hd__mux2_2 _23244_ (.A0(mem_la_addr[31]),
    .A1(mem_addr[31]),
    .S(_17225_),
    .X(_03088_));
 sky130_fd_sc_hd__mux2_2 _23245_ (.A0(mem_la_addr[30]),
    .A1(mem_addr[30]),
    .S(_17225_),
    .X(_03087_));
 sky130_fd_sc_hd__mux2_2 _23246_ (.A0(mem_la_addr[29]),
    .A1(mem_addr[29]),
    .S(_17225_),
    .X(_03086_));
 sky130_fd_sc_hd__buf_1 _23247_ (.A(_17223_),
    .X(_19125_));
 sky130_fd_sc_hd__buf_1 _23248_ (.A(_19125_),
    .X(_19126_));
 sky130_fd_sc_hd__mux2_2 _23249_ (.A0(mem_la_addr[28]),
    .A1(mem_addr[28]),
    .S(_19126_),
    .X(_03085_));
 sky130_fd_sc_hd__mux2_2 _23250_ (.A0(mem_la_addr[27]),
    .A1(mem_addr[27]),
    .S(_19126_),
    .X(_03084_));
 sky130_fd_sc_hd__mux2_2 _23251_ (.A0(mem_la_addr[26]),
    .A1(mem_addr[26]),
    .S(_19126_),
    .X(_03083_));
 sky130_fd_sc_hd__mux2_2 _23252_ (.A0(mem_la_addr[25]),
    .A1(mem_addr[25]),
    .S(_19126_),
    .X(_03082_));
 sky130_fd_sc_hd__buf_1 _23253_ (.A(_19125_),
    .X(_19127_));
 sky130_fd_sc_hd__mux2_2 _23254_ (.A0(mem_la_addr[24]),
    .A1(mem_addr[24]),
    .S(_19127_),
    .X(_03081_));
 sky130_fd_sc_hd__mux2_2 _23255_ (.A0(mem_la_addr[23]),
    .A1(mem_addr[23]),
    .S(_19127_),
    .X(_03080_));
 sky130_fd_sc_hd__mux2_2 _23256_ (.A0(mem_la_addr[22]),
    .A1(mem_addr[22]),
    .S(_19127_),
    .X(_03079_));
 sky130_fd_sc_hd__mux2_2 _23257_ (.A0(mem_la_addr[21]),
    .A1(mem_addr[21]),
    .S(_19127_),
    .X(_03078_));
 sky130_fd_sc_hd__buf_1 _23258_ (.A(_19125_),
    .X(_19128_));
 sky130_fd_sc_hd__mux2_2 _23259_ (.A0(mem_la_addr[20]),
    .A1(mem_addr[20]),
    .S(_19128_),
    .X(_03077_));
 sky130_fd_sc_hd__mux2_2 _23260_ (.A0(mem_la_addr[19]),
    .A1(mem_addr[19]),
    .S(_19128_),
    .X(_03076_));
 sky130_fd_sc_hd__mux2_2 _23261_ (.A0(mem_la_addr[18]),
    .A1(mem_addr[18]),
    .S(_19128_),
    .X(_03075_));
 sky130_fd_sc_hd__mux2_2 _23262_ (.A0(mem_la_addr[17]),
    .A1(mem_addr[17]),
    .S(_19128_),
    .X(_03074_));
 sky130_fd_sc_hd__buf_1 _23263_ (.A(_19125_),
    .X(_19129_));
 sky130_fd_sc_hd__mux2_2 _23264_ (.A0(mem_la_addr[16]),
    .A1(mem_addr[16]),
    .S(_19129_),
    .X(_03073_));
 sky130_fd_sc_hd__mux2_2 _23265_ (.A0(mem_la_addr[15]),
    .A1(mem_addr[15]),
    .S(_19129_),
    .X(_03072_));
 sky130_fd_sc_hd__mux2_2 _23266_ (.A0(mem_la_addr[14]),
    .A1(mem_addr[14]),
    .S(_19129_),
    .X(_03071_));
 sky130_fd_sc_hd__mux2_2 _23267_ (.A0(mem_la_addr[13]),
    .A1(mem_addr[13]),
    .S(_19129_),
    .X(_03070_));
 sky130_fd_sc_hd__buf_1 _23268_ (.A(_17223_),
    .X(_19130_));
 sky130_fd_sc_hd__mux2_2 _23269_ (.A0(mem_la_addr[12]),
    .A1(mem_addr[12]),
    .S(_19130_),
    .X(_03069_));
 sky130_fd_sc_hd__mux2_2 _23270_ (.A0(mem_la_addr[11]),
    .A1(mem_addr[11]),
    .S(_19130_),
    .X(_03068_));
 sky130_fd_sc_hd__mux2_2 _23271_ (.A0(mem_la_addr[10]),
    .A1(mem_addr[10]),
    .S(_19130_),
    .X(_03067_));
 sky130_fd_sc_hd__mux2_2 _23272_ (.A0(mem_la_addr[9]),
    .A1(mem_addr[9]),
    .S(_19130_),
    .X(_03066_));
 sky130_fd_sc_hd__buf_1 _23273_ (.A(_17223_),
    .X(_19131_));
 sky130_fd_sc_hd__mux2_2 _23274_ (.A0(mem_la_addr[8]),
    .A1(mem_addr[8]),
    .S(_19131_),
    .X(_03065_));
 sky130_fd_sc_hd__mux2_2 _23275_ (.A0(mem_la_addr[7]),
    .A1(mem_addr[7]),
    .S(_19131_),
    .X(_03064_));
 sky130_fd_sc_hd__mux2_2 _23276_ (.A0(mem_la_addr[6]),
    .A1(mem_addr[6]),
    .S(_19131_),
    .X(_03063_));
 sky130_fd_sc_hd__mux2_2 _23277_ (.A0(mem_la_addr[5]),
    .A1(mem_addr[5]),
    .S(_19131_),
    .X(_03062_));
 sky130_fd_sc_hd__mux2_2 _23278_ (.A0(mem_la_addr[4]),
    .A1(mem_addr[4]),
    .S(_17224_),
    .X(_03061_));
 sky130_fd_sc_hd__mux2_2 _23279_ (.A0(mem_la_addr[3]),
    .A1(mem_addr[3]),
    .S(_17224_),
    .X(_03060_));
 sky130_fd_sc_hd__mux2_2 _23280_ (.A0(mem_la_addr[2]),
    .A1(mem_addr[2]),
    .S(_17224_),
    .X(_03059_));
 sky130_fd_sc_hd__buf_1 _23281_ (.A(\pcpi_mul.rs1[31] ),
    .X(_19132_));
 sky130_fd_sc_hd__buf_1 _23282_ (.A(_19132_),
    .X(_19133_));
 sky130_fd_sc_hd__buf_1 _23283_ (.A(_19133_),
    .X(_19134_));
 sky130_fd_sc_hd__buf_1 _23284_ (.A(_19134_),
    .X(_19135_));
 sky130_fd_sc_hd__buf_1 _23285_ (.A(_19135_),
    .X(_19136_));
 sky130_fd_sc_hd__buf_1 _23286_ (.A(_19136_),
    .X(_19137_));
 sky130_fd_sc_hd__a21o_2 _23287_ (.A1(_19137_),
    .A2(_18700_),
    .B1(_16959_),
    .X(_03058_));
 sky130_fd_sc_hd__buf_1 _23288_ (.A(\pcpi_mul.rs1[30] ),
    .X(_19138_));
 sky130_fd_sc_hd__buf_1 _23289_ (.A(_19138_),
    .X(_19139_));
 sky130_vsdinv _23290_ (.A(_19139_),
    .Y(_19140_));
 sky130_fd_sc_hd__buf_1 _23291_ (.A(_19140_),
    .X(_19141_));
 sky130_fd_sc_hd__nand2_2 _23292_ (.A(_18863_),
    .B(_19042_),
    .Y(_19142_));
 sky130_fd_sc_hd__o21ai_2 _23293_ (.A1(_19141_),
    .A2(_18861_),
    .B1(_19142_),
    .Y(_03057_));
 sky130_fd_sc_hd__buf_1 _23294_ (.A(\pcpi_mul.rs1[29] ),
    .X(_19143_));
 sky130_fd_sc_hd__buf_1 _23295_ (.A(_19143_),
    .X(_19144_));
 sky130_vsdinv _23296_ (.A(_19144_),
    .Y(_19145_));
 sky130_fd_sc_hd__buf_1 _23297_ (.A(_19145_),
    .X(_19146_));
 sky130_fd_sc_hd__buf_1 _23298_ (.A(_19146_),
    .X(_19147_));
 sky130_fd_sc_hd__nand2_2 _23299_ (.A(_18863_),
    .B(_19044_),
    .Y(_19148_));
 sky130_fd_sc_hd__o21ai_2 _23300_ (.A1(_19147_),
    .A2(_18861_),
    .B1(_19148_),
    .Y(_03056_));
 sky130_fd_sc_hd__buf_1 _23301_ (.A(\pcpi_mul.rs1[28] ),
    .X(_19149_));
 sky130_vsdinv _23302_ (.A(_19149_),
    .Y(_19150_));
 sky130_fd_sc_hd__buf_1 _23303_ (.A(_19150_),
    .X(_19151_));
 sky130_fd_sc_hd__buf_1 _23304_ (.A(_19151_),
    .X(_19152_));
 sky130_fd_sc_hd__buf_1 _23305_ (.A(_18860_),
    .X(_19153_));
 sky130_fd_sc_hd__buf_1 _23306_ (.A(_18862_),
    .X(_19154_));
 sky130_fd_sc_hd__nand2_2 _23307_ (.A(_19154_),
    .B(_19046_),
    .Y(_19155_));
 sky130_fd_sc_hd__o21ai_2 _23308_ (.A1(_19152_),
    .A2(_19153_),
    .B1(_19155_),
    .Y(_03055_));
 sky130_fd_sc_hd__buf_1 _23309_ (.A(\pcpi_mul.rs1[27] ),
    .X(_19156_));
 sky130_vsdinv _23310_ (.A(_19156_),
    .Y(_19157_));
 sky130_fd_sc_hd__buf_1 _23311_ (.A(_19157_),
    .X(_19158_));
 sky130_fd_sc_hd__buf_1 _23312_ (.A(_19158_),
    .X(_19159_));
 sky130_fd_sc_hd__nand2_2 _23313_ (.A(_19154_),
    .B(_19048_),
    .Y(_19160_));
 sky130_fd_sc_hd__o21ai_2 _23314_ (.A1(_19159_),
    .A2(_19153_),
    .B1(_19160_),
    .Y(_03054_));
 sky130_fd_sc_hd__buf_1 _23315_ (.A(\pcpi_mul.rs1[26] ),
    .X(_19161_));
 sky130_fd_sc_hd__buf_1 _23316_ (.A(_19161_),
    .X(_19162_));
 sky130_vsdinv _23317_ (.A(_19162_),
    .Y(_19163_));
 sky130_fd_sc_hd__buf_1 _23318_ (.A(_19163_),
    .X(_19164_));
 sky130_fd_sc_hd__nand2_2 _23319_ (.A(_19154_),
    .B(_19051_),
    .Y(_19165_));
 sky130_fd_sc_hd__o21ai_2 _23320_ (.A1(_19164_),
    .A2(_19153_),
    .B1(_19165_),
    .Y(_03053_));
 sky130_fd_sc_hd__buf_1 _23321_ (.A(\pcpi_mul.rs1[25] ),
    .X(_19166_));
 sky130_fd_sc_hd__buf_1 _23322_ (.A(_19166_),
    .X(_19167_));
 sky130_vsdinv _23323_ (.A(_19167_),
    .Y(_19168_));
 sky130_fd_sc_hd__buf_1 _23324_ (.A(_19168_),
    .X(_19169_));
 sky130_fd_sc_hd__nand2_2 _23325_ (.A(_19154_),
    .B(_19053_),
    .Y(_19170_));
 sky130_fd_sc_hd__o21ai_2 _23326_ (.A1(_19169_),
    .A2(_19153_),
    .B1(_19170_),
    .Y(_03052_));
 sky130_fd_sc_hd__buf_1 _23327_ (.A(\pcpi_mul.rs1[24] ),
    .X(_19171_));
 sky130_fd_sc_hd__buf_1 _23328_ (.A(_19171_),
    .X(_19172_));
 sky130_vsdinv _23329_ (.A(_19172_),
    .Y(_19173_));
 sky130_fd_sc_hd__buf_1 _23330_ (.A(_19173_),
    .X(_19174_));
 sky130_fd_sc_hd__buf_1 _23331_ (.A(_19174_),
    .X(_19175_));
 sky130_fd_sc_hd__buf_1 _23332_ (.A(_18860_),
    .X(_19176_));
 sky130_fd_sc_hd__buf_1 _23333_ (.A(_18862_),
    .X(_19177_));
 sky130_fd_sc_hd__nand2_2 _23334_ (.A(_19177_),
    .B(_19055_),
    .Y(_19178_));
 sky130_fd_sc_hd__o21ai_2 _23335_ (.A1(_19175_),
    .A2(_19176_),
    .B1(_19178_),
    .Y(_03051_));
 sky130_fd_sc_hd__buf_1 _23336_ (.A(\pcpi_mul.rs1[23] ),
    .X(_19179_));
 sky130_fd_sc_hd__buf_1 _23337_ (.A(_19179_),
    .X(_19180_));
 sky130_vsdinv _23338_ (.A(_19180_),
    .Y(_19181_));
 sky130_fd_sc_hd__buf_1 _23339_ (.A(_19181_),
    .X(_19182_));
 sky130_fd_sc_hd__nand2_2 _23340_ (.A(_19177_),
    .B(_19057_),
    .Y(_19183_));
 sky130_fd_sc_hd__o21ai_2 _23341_ (.A1(_19182_),
    .A2(_19176_),
    .B1(_19183_),
    .Y(_03050_));
 sky130_fd_sc_hd__buf_1 _23342_ (.A(\pcpi_mul.rs1[22] ),
    .X(_19184_));
 sky130_fd_sc_hd__buf_1 _23343_ (.A(_19184_),
    .X(_19185_));
 sky130_vsdinv _23344_ (.A(_19185_),
    .Y(_19186_));
 sky130_fd_sc_hd__buf_1 _23345_ (.A(_19186_),
    .X(_19187_));
 sky130_fd_sc_hd__buf_1 _23346_ (.A(_19187_),
    .X(_19188_));
 sky130_fd_sc_hd__nand2_2 _23347_ (.A(_19177_),
    .B(_19060_),
    .Y(_19189_));
 sky130_fd_sc_hd__o21ai_2 _23348_ (.A1(_19188_),
    .A2(_19176_),
    .B1(_19189_),
    .Y(_03049_));
 sky130_fd_sc_hd__buf_1 _23349_ (.A(\pcpi_mul.rs1[21] ),
    .X(_19190_));
 sky130_vsdinv _23350_ (.A(_19190_),
    .Y(_19191_));
 sky130_fd_sc_hd__buf_1 _23351_ (.A(_19191_),
    .X(_19192_));
 sky130_fd_sc_hd__buf_1 _23352_ (.A(_19192_),
    .X(_19193_));
 sky130_fd_sc_hd__nand2_2 _23353_ (.A(_19177_),
    .B(_19062_),
    .Y(_19194_));
 sky130_fd_sc_hd__o21ai_2 _23354_ (.A1(_19193_),
    .A2(_19176_),
    .B1(_19194_),
    .Y(_03048_));
 sky130_fd_sc_hd__buf_1 _23355_ (.A(\pcpi_mul.rs1[20] ),
    .X(_19195_));
 sky130_fd_sc_hd__buf_1 _23356_ (.A(_19195_),
    .X(_19196_));
 sky130_vsdinv _23357_ (.A(_19196_),
    .Y(_19197_));
 sky130_fd_sc_hd__buf_1 _23358_ (.A(_19197_),
    .X(_19198_));
 sky130_fd_sc_hd__buf_1 _23359_ (.A(_18860_),
    .X(_19199_));
 sky130_fd_sc_hd__buf_1 _23360_ (.A(_18862_),
    .X(_19200_));
 sky130_fd_sc_hd__nand2_2 _23361_ (.A(_19200_),
    .B(_19064_),
    .Y(_19201_));
 sky130_fd_sc_hd__o21ai_2 _23362_ (.A1(_19198_),
    .A2(_19199_),
    .B1(_19201_),
    .Y(_03047_));
 sky130_fd_sc_hd__buf_1 _23363_ (.A(\pcpi_mul.rs1[19] ),
    .X(_19202_));
 sky130_fd_sc_hd__buf_1 _23364_ (.A(_19202_),
    .X(_19203_));
 sky130_vsdinv _23365_ (.A(_19203_),
    .Y(_19204_));
 sky130_fd_sc_hd__buf_1 _23366_ (.A(_19204_),
    .X(_19205_));
 sky130_fd_sc_hd__nand2_2 _23367_ (.A(_19200_),
    .B(_19066_),
    .Y(_19206_));
 sky130_fd_sc_hd__o21ai_2 _23368_ (.A1(_19205_),
    .A2(_19199_),
    .B1(_19206_),
    .Y(_03046_));
 sky130_fd_sc_hd__buf_1 _23369_ (.A(\pcpi_mul.rs1[18] ),
    .X(_19207_));
 sky130_vsdinv _23370_ (.A(_19207_),
    .Y(_19208_));
 sky130_fd_sc_hd__buf_1 _23371_ (.A(_19208_),
    .X(_19209_));
 sky130_fd_sc_hd__nand2_2 _23372_ (.A(_19200_),
    .B(_19069_),
    .Y(_19210_));
 sky130_fd_sc_hd__o21ai_2 _23373_ (.A1(_19209_),
    .A2(_19199_),
    .B1(_19210_),
    .Y(_03045_));
 sky130_fd_sc_hd__buf_1 _23374_ (.A(\pcpi_mul.rs1[17] ),
    .X(_19211_));
 sky130_vsdinv _23375_ (.A(_19211_),
    .Y(_19212_));
 sky130_fd_sc_hd__buf_1 _23376_ (.A(_19212_),
    .X(_19213_));
 sky130_fd_sc_hd__nand2_2 _23377_ (.A(_19200_),
    .B(_19072_),
    .Y(_19214_));
 sky130_fd_sc_hd__o21ai_2 _23378_ (.A1(_19213_),
    .A2(_19199_),
    .B1(_19214_),
    .Y(_03044_));
 sky130_fd_sc_hd__buf_1 _23379_ (.A(\pcpi_mul.rs1[16] ),
    .X(_19215_));
 sky130_fd_sc_hd__buf_1 _23380_ (.A(_19215_),
    .X(_19216_));
 sky130_vsdinv _23381_ (.A(_19216_),
    .Y(_19217_));
 sky130_fd_sc_hd__buf_1 _23382_ (.A(_19217_),
    .X(_19218_));
 sky130_fd_sc_hd__buf_1 _23383_ (.A(_16956_),
    .X(_19219_));
 sky130_fd_sc_hd__buf_1 _23384_ (.A(_19219_),
    .X(_19220_));
 sky130_fd_sc_hd__buf_1 _23385_ (.A(_16964_),
    .X(_19221_));
 sky130_fd_sc_hd__buf_1 _23386_ (.A(_19221_),
    .X(_19222_));
 sky130_fd_sc_hd__nand2_2 _23387_ (.A(_19222_),
    .B(_19075_),
    .Y(_19223_));
 sky130_fd_sc_hd__o21ai_2 _23388_ (.A1(_19218_),
    .A2(_19220_),
    .B1(_19223_),
    .Y(_03043_));
 sky130_fd_sc_hd__buf_1 _23389_ (.A(\pcpi_mul.rs1[15] ),
    .X(_19224_));
 sky130_fd_sc_hd__buf_1 _23390_ (.A(_19224_),
    .X(_19225_));
 sky130_vsdinv _23391_ (.A(_19225_),
    .Y(_19226_));
 sky130_fd_sc_hd__buf_1 _23392_ (.A(_19226_),
    .X(_19227_));
 sky130_fd_sc_hd__buf_1 _23393_ (.A(_19227_),
    .X(_19228_));
 sky130_fd_sc_hd__nand2_2 _23394_ (.A(_19222_),
    .B(_19077_),
    .Y(_19229_));
 sky130_fd_sc_hd__o21ai_2 _23395_ (.A1(_19228_),
    .A2(_19220_),
    .B1(_19229_),
    .Y(_03042_));
 sky130_fd_sc_hd__buf_1 _23396_ (.A(\pcpi_mul.rs1[14] ),
    .X(_19230_));
 sky130_fd_sc_hd__buf_1 _23397_ (.A(_19230_),
    .X(_19231_));
 sky130_vsdinv _23398_ (.A(_19231_),
    .Y(_19232_));
 sky130_fd_sc_hd__buf_1 _23399_ (.A(_19232_),
    .X(_19233_));
 sky130_fd_sc_hd__buf_1 _23400_ (.A(_19233_),
    .X(_19234_));
 sky130_fd_sc_hd__nand2_2 _23401_ (.A(_19222_),
    .B(_19081_),
    .Y(_19235_));
 sky130_fd_sc_hd__o21ai_2 _23402_ (.A1(_19234_),
    .A2(_19220_),
    .B1(_19235_),
    .Y(_03041_));
 sky130_fd_sc_hd__buf_1 _23403_ (.A(\pcpi_mul.rs1[13] ),
    .X(_19236_));
 sky130_fd_sc_hd__buf_1 _23404_ (.A(_19236_),
    .X(_19237_));
 sky130_vsdinv _23405_ (.A(_19237_),
    .Y(_19238_));
 sky130_fd_sc_hd__buf_1 _23406_ (.A(_19238_),
    .X(_19239_));
 sky130_fd_sc_hd__nand2_2 _23407_ (.A(_19222_),
    .B(_19083_),
    .Y(_19240_));
 sky130_fd_sc_hd__o21ai_2 _23408_ (.A1(_19239_),
    .A2(_19220_),
    .B1(_19240_),
    .Y(_03040_));
 sky130_fd_sc_hd__buf_1 _23409_ (.A(\pcpi_mul.rs1[12] ),
    .X(_19241_));
 sky130_fd_sc_hd__buf_1 _23410_ (.A(_19241_),
    .X(_19242_));
 sky130_vsdinv _23411_ (.A(_19242_),
    .Y(_19243_));
 sky130_fd_sc_hd__buf_1 _23412_ (.A(_19243_),
    .X(_19244_));
 sky130_fd_sc_hd__buf_1 _23413_ (.A(_19219_),
    .X(_19245_));
 sky130_fd_sc_hd__buf_1 _23414_ (.A(_19221_),
    .X(_19246_));
 sky130_fd_sc_hd__nand2_2 _23415_ (.A(_19246_),
    .B(_19085_),
    .Y(_19247_));
 sky130_fd_sc_hd__o21ai_2 _23416_ (.A1(_19244_),
    .A2(_19245_),
    .B1(_19247_),
    .Y(_03039_));
 sky130_fd_sc_hd__buf_1 _23417_ (.A(\pcpi_mul.rs1[11] ),
    .X(_19248_));
 sky130_vsdinv _23418_ (.A(_19248_),
    .Y(_19249_));
 sky130_fd_sc_hd__buf_1 _23419_ (.A(_19249_),
    .X(_19250_));
 sky130_fd_sc_hd__nand2_2 _23420_ (.A(_19246_),
    .B(_19087_),
    .Y(_19251_));
 sky130_fd_sc_hd__o21ai_2 _23421_ (.A1(_19250_),
    .A2(_19245_),
    .B1(_19251_),
    .Y(_03038_));
 sky130_fd_sc_hd__buf_1 _23422_ (.A(\pcpi_mul.rs1[10] ),
    .X(_19252_));
 sky130_vsdinv _23423_ (.A(_19252_),
    .Y(_19253_));
 sky130_fd_sc_hd__buf_1 _23424_ (.A(_19253_),
    .X(_19254_));
 sky130_fd_sc_hd__nand2_2 _23425_ (.A(_19246_),
    .B(_19090_),
    .Y(_19255_));
 sky130_fd_sc_hd__o21ai_2 _23426_ (.A1(_19254_),
    .A2(_19245_),
    .B1(_19255_),
    .Y(_03037_));
 sky130_fd_sc_hd__buf_1 _23427_ (.A(\pcpi_mul.rs1[9] ),
    .X(_19256_));
 sky130_fd_sc_hd__buf_1 _23428_ (.A(_19256_),
    .X(_19257_));
 sky130_vsdinv _23429_ (.A(_19257_),
    .Y(_19258_));
 sky130_fd_sc_hd__buf_1 _23430_ (.A(_19258_),
    .X(_19259_));
 sky130_fd_sc_hd__nand2_2 _23431_ (.A(_19246_),
    .B(_19093_),
    .Y(_19260_));
 sky130_fd_sc_hd__o21ai_2 _23432_ (.A1(_19259_),
    .A2(_19245_),
    .B1(_19260_),
    .Y(_03036_));
 sky130_fd_sc_hd__buf_1 _23433_ (.A(\pcpi_mul.rs1[8] ),
    .X(_19261_));
 sky130_vsdinv _23434_ (.A(_19261_),
    .Y(_19262_));
 sky130_fd_sc_hd__buf_1 _23435_ (.A(_19262_),
    .X(_19263_));
 sky130_fd_sc_hd__buf_1 _23436_ (.A(_19219_),
    .X(_19264_));
 sky130_fd_sc_hd__buf_1 _23437_ (.A(_19221_),
    .X(_19265_));
 sky130_fd_sc_hd__nand2_2 _23438_ (.A(_19265_),
    .B(_19096_),
    .Y(_19266_));
 sky130_fd_sc_hd__o21ai_2 _23439_ (.A1(_19263_),
    .A2(_19264_),
    .B1(_19266_),
    .Y(_03035_));
 sky130_fd_sc_hd__buf_1 _23440_ (.A(\pcpi_mul.rs1[7] ),
    .X(_19267_));
 sky130_vsdinv _23441_ (.A(_19267_),
    .Y(_19268_));
 sky130_fd_sc_hd__buf_1 _23442_ (.A(_19268_),
    .X(_19269_));
 sky130_fd_sc_hd__nand2_2 _23443_ (.A(_19265_),
    .B(_19099_),
    .Y(_19270_));
 sky130_fd_sc_hd__o21ai_2 _23444_ (.A1(_19269_),
    .A2(_19264_),
    .B1(_19270_),
    .Y(_03034_));
 sky130_fd_sc_hd__buf_1 _23445_ (.A(\pcpi_mul.rs1[6] ),
    .X(_19271_));
 sky130_fd_sc_hd__buf_1 _23446_ (.A(_19271_),
    .X(_19272_));
 sky130_fd_sc_hd__buf_1 _23447_ (.A(_19272_),
    .X(_19273_));
 sky130_vsdinv _23448_ (.A(_19273_),
    .Y(_19274_));
 sky130_fd_sc_hd__buf_1 _23449_ (.A(_19274_),
    .X(_19275_));
 sky130_fd_sc_hd__nand2_2 _23450_ (.A(_19265_),
    .B(_19103_),
    .Y(_19276_));
 sky130_fd_sc_hd__o21ai_2 _23451_ (.A1(_19275_),
    .A2(_19264_),
    .B1(_19276_),
    .Y(_03033_));
 sky130_fd_sc_hd__buf_1 _23452_ (.A(\pcpi_mul.rs1[5] ),
    .X(_19277_));
 sky130_vsdinv _23453_ (.A(_19277_),
    .Y(_19278_));
 sky130_fd_sc_hd__buf_1 _23454_ (.A(_19278_),
    .X(_19279_));
 sky130_fd_sc_hd__nand2_2 _23455_ (.A(_19265_),
    .B(_19105_),
    .Y(_19280_));
 sky130_fd_sc_hd__o21ai_2 _23456_ (.A1(_19279_),
    .A2(_19264_),
    .B1(_19280_),
    .Y(_03032_));
 sky130_fd_sc_hd__buf_1 _23457_ (.A(\pcpi_mul.rs1[4] ),
    .X(_19281_));
 sky130_vsdinv _23458_ (.A(_19281_),
    .Y(_19282_));
 sky130_fd_sc_hd__buf_1 _23459_ (.A(_19282_),
    .X(_19283_));
 sky130_fd_sc_hd__buf_1 _23460_ (.A(_19219_),
    .X(_19284_));
 sky130_fd_sc_hd__buf_1 _23461_ (.A(_19221_),
    .X(_19285_));
 sky130_fd_sc_hd__nand2_2 _23462_ (.A(_19285_),
    .B(_19108_),
    .Y(_19286_));
 sky130_fd_sc_hd__o21ai_2 _23463_ (.A1(_19283_),
    .A2(_19284_),
    .B1(_19286_),
    .Y(_03031_));
 sky130_fd_sc_hd__buf_1 _23464_ (.A(\pcpi_mul.rs1[3] ),
    .X(_19287_));
 sky130_vsdinv _23465_ (.A(_19287_),
    .Y(_19288_));
 sky130_fd_sc_hd__buf_1 _23466_ (.A(_19288_),
    .X(_19289_));
 sky130_fd_sc_hd__buf_1 _23467_ (.A(_19289_),
    .X(_19290_));
 sky130_fd_sc_hd__nand2_2 _23468_ (.A(_19285_),
    .B(_19110_),
    .Y(_19291_));
 sky130_fd_sc_hd__o21ai_2 _23469_ (.A1(_19290_),
    .A2(_19284_),
    .B1(_19291_),
    .Y(_03030_));
 sky130_fd_sc_hd__buf_1 _23470_ (.A(\pcpi_mul.rs1[2] ),
    .X(_19292_));
 sky130_fd_sc_hd__buf_1 _23471_ (.A(_19292_),
    .X(_19293_));
 sky130_vsdinv _23472_ (.A(_19293_),
    .Y(_19294_));
 sky130_fd_sc_hd__buf_1 _23473_ (.A(_19294_),
    .X(_19295_));
 sky130_fd_sc_hd__nand2_2 _23474_ (.A(_19285_),
    .B(_19113_),
    .Y(_19296_));
 sky130_fd_sc_hd__o21ai_2 _23475_ (.A1(_19295_),
    .A2(_19284_),
    .B1(_19296_),
    .Y(_03029_));
 sky130_fd_sc_hd__buf_1 _23476_ (.A(\pcpi_mul.rs1[1] ),
    .X(_19297_));
 sky130_vsdinv _23477_ (.A(_19297_),
    .Y(_19298_));
 sky130_fd_sc_hd__nand2_2 _23478_ (.A(_19285_),
    .B(_19118_),
    .Y(_19299_));
 sky130_fd_sc_hd__o21ai_2 _23479_ (.A1(_19298_),
    .A2(_19284_),
    .B1(_19299_),
    .Y(_03028_));
 sky130_fd_sc_hd__buf_1 _23480_ (.A(\pcpi_mul.rs1[0] ),
    .X(_19300_));
 sky130_fd_sc_hd__buf_1 _23481_ (.A(_19300_),
    .X(_19301_));
 sky130_vsdinv _23482_ (.A(_19301_),
    .Y(_19302_));
 sky130_fd_sc_hd__nand2_2 _23483_ (.A(_16975_),
    .B(_19124_),
    .Y(_19303_));
 sky130_fd_sc_hd__o21ai_2 _23484_ (.A1(_19302_),
    .A2(_16966_),
    .B1(_19303_),
    .Y(_03027_));
 sky130_fd_sc_hd__buf_1 _23485_ (.A(_18280_),
    .X(_19304_));
 sky130_fd_sc_hd__buf_1 _23486_ (.A(_18293_),
    .X(_19305_));
 sky130_fd_sc_hd__o2111ai_2 _23487_ (.A1(_18890_),
    .A2(_19304_),
    .B1(_18290_),
    .C1(_18370_),
    .D1(_19305_),
    .Y(_19306_));
 sky130_fd_sc_hd__buf_1 _23488_ (.A(_19306_),
    .X(_19307_));
 sky130_fd_sc_hd__buf_1 _23489_ (.A(_19307_),
    .X(_19308_));
 sky130_fd_sc_hd__mux2_2 _23490_ (.A0(_18650_),
    .A1(\cpuregs[5][31] ),
    .S(_19308_),
    .X(_03026_));
 sky130_fd_sc_hd__mux2_2 _23491_ (.A0(_18654_),
    .A1(\cpuregs[5][30] ),
    .S(_19308_),
    .X(_03025_));
 sky130_fd_sc_hd__mux2_2 _23492_ (.A0(_18655_),
    .A1(\cpuregs[5][29] ),
    .S(_19308_),
    .X(_03024_));
 sky130_fd_sc_hd__mux2_2 _23493_ (.A0(_18656_),
    .A1(\cpuregs[5][28] ),
    .S(_19308_),
    .X(_03023_));
 sky130_fd_sc_hd__buf_1 _23494_ (.A(_19307_),
    .X(_19309_));
 sky130_fd_sc_hd__mux2_2 _23495_ (.A0(_18657_),
    .A1(\cpuregs[5][27] ),
    .S(_19309_),
    .X(_03022_));
 sky130_fd_sc_hd__mux2_2 _23496_ (.A0(_18659_),
    .A1(\cpuregs[5][26] ),
    .S(_19309_),
    .X(_03021_));
 sky130_fd_sc_hd__mux2_2 _23497_ (.A0(_18660_),
    .A1(\cpuregs[5][25] ),
    .S(_19309_),
    .X(_03020_));
 sky130_fd_sc_hd__mux2_2 _23498_ (.A0(_18661_),
    .A1(\cpuregs[5][24] ),
    .S(_19309_),
    .X(_03019_));
 sky130_fd_sc_hd__buf_1 _23499_ (.A(_19307_),
    .X(_19310_));
 sky130_fd_sc_hd__mux2_2 _23500_ (.A0(_18662_),
    .A1(\cpuregs[5][23] ),
    .S(_19310_),
    .X(_03018_));
 sky130_fd_sc_hd__mux2_2 _23501_ (.A0(_18664_),
    .A1(\cpuregs[5][22] ),
    .S(_19310_),
    .X(_03017_));
 sky130_fd_sc_hd__mux2_2 _23502_ (.A0(_18665_),
    .A1(\cpuregs[5][21] ),
    .S(_19310_),
    .X(_03016_));
 sky130_fd_sc_hd__mux2_2 _23503_ (.A0(_18666_),
    .A1(\cpuregs[5][20] ),
    .S(_19310_),
    .X(_03015_));
 sky130_fd_sc_hd__buf_1 _23504_ (.A(_19307_),
    .X(_19311_));
 sky130_fd_sc_hd__mux2_2 _23505_ (.A0(_18667_),
    .A1(\cpuregs[5][19] ),
    .S(_19311_),
    .X(_03014_));
 sky130_fd_sc_hd__mux2_2 _23506_ (.A0(_18669_),
    .A1(\cpuregs[5][18] ),
    .S(_19311_),
    .X(_03013_));
 sky130_fd_sc_hd__mux2_2 _23507_ (.A0(_18670_),
    .A1(\cpuregs[5][17] ),
    .S(_19311_),
    .X(_03012_));
 sky130_fd_sc_hd__mux2_2 _23508_ (.A0(_18671_),
    .A1(\cpuregs[5][16] ),
    .S(_19311_),
    .X(_03011_));
 sky130_fd_sc_hd__buf_1 _23509_ (.A(_19306_),
    .X(_19312_));
 sky130_fd_sc_hd__buf_1 _23510_ (.A(_19312_),
    .X(_19313_));
 sky130_fd_sc_hd__mux2_2 _23511_ (.A0(_18672_),
    .A1(\cpuregs[5][15] ),
    .S(_19313_),
    .X(_03010_));
 sky130_fd_sc_hd__mux2_2 _23512_ (.A0(_18675_),
    .A1(\cpuregs[5][14] ),
    .S(_19313_),
    .X(_03009_));
 sky130_fd_sc_hd__mux2_2 _23513_ (.A0(_18676_),
    .A1(\cpuregs[5][13] ),
    .S(_19313_),
    .X(_03008_));
 sky130_fd_sc_hd__mux2_2 _23514_ (.A0(_18677_),
    .A1(\cpuregs[5][12] ),
    .S(_19313_),
    .X(_03007_));
 sky130_fd_sc_hd__buf_1 _23515_ (.A(_19312_),
    .X(_19314_));
 sky130_fd_sc_hd__mux2_2 _23516_ (.A0(_18678_),
    .A1(\cpuregs[5][11] ),
    .S(_19314_),
    .X(_03006_));
 sky130_fd_sc_hd__mux2_2 _23517_ (.A0(_18680_),
    .A1(\cpuregs[5][10] ),
    .S(_19314_),
    .X(_03005_));
 sky130_fd_sc_hd__mux2_2 _23518_ (.A0(_18681_),
    .A1(\cpuregs[5][9] ),
    .S(_19314_),
    .X(_03004_));
 sky130_fd_sc_hd__mux2_2 _23519_ (.A0(_18682_),
    .A1(\cpuregs[5][8] ),
    .S(_19314_),
    .X(_03003_));
 sky130_fd_sc_hd__buf_1 _23520_ (.A(_19312_),
    .X(_19315_));
 sky130_fd_sc_hd__mux2_2 _23521_ (.A0(_18683_),
    .A1(\cpuregs[5][7] ),
    .S(_19315_),
    .X(_03002_));
 sky130_fd_sc_hd__mux2_2 _23522_ (.A0(_18685_),
    .A1(\cpuregs[5][6] ),
    .S(_19315_),
    .X(_03001_));
 sky130_fd_sc_hd__mux2_2 _23523_ (.A0(_18686_),
    .A1(\cpuregs[5][5] ),
    .S(_19315_),
    .X(_03000_));
 sky130_fd_sc_hd__mux2_2 _23524_ (.A0(_18687_),
    .A1(\cpuregs[5][4] ),
    .S(_19315_),
    .X(_02999_));
 sky130_fd_sc_hd__buf_1 _23525_ (.A(_19312_),
    .X(_19316_));
 sky130_fd_sc_hd__mux2_2 _23526_ (.A0(_18688_),
    .A1(\cpuregs[5][3] ),
    .S(_19316_),
    .X(_02998_));
 sky130_fd_sc_hd__mux2_2 _23527_ (.A0(_18690_),
    .A1(\cpuregs[5][2] ),
    .S(_19316_),
    .X(_02997_));
 sky130_fd_sc_hd__mux2_2 _23528_ (.A0(_18691_),
    .A1(\cpuregs[5][1] ),
    .S(_19316_),
    .X(_02996_));
 sky130_fd_sc_hd__mux2_2 _23529_ (.A0(_18692_),
    .A1(\cpuregs[5][0] ),
    .S(_19316_),
    .X(_02995_));
 sky130_fd_sc_hd__and3b_2 _23530_ (.A_N(_18281_),
    .B(_18457_),
    .C(_18285_),
    .X(_19317_));
 sky130_fd_sc_hd__buf_1 _23531_ (.A(_19317_),
    .X(_19318_));
 sky130_fd_sc_hd__buf_1 _23532_ (.A(_19318_),
    .X(_19319_));
 sky130_fd_sc_hd__mux2_2 _23533_ (.A0(\cpuregs[2][31] ),
    .A1(_18272_),
    .S(_19319_),
    .X(_02994_));
 sky130_fd_sc_hd__mux2_2 _23534_ (.A0(\cpuregs[2][30] ),
    .A1(_18298_),
    .S(_19319_),
    .X(_02993_));
 sky130_fd_sc_hd__mux2_2 _23535_ (.A0(\cpuregs[2][29] ),
    .A1(_18300_),
    .S(_19319_),
    .X(_02992_));
 sky130_fd_sc_hd__mux2_2 _23536_ (.A0(\cpuregs[2][28] ),
    .A1(_18302_),
    .S(_19319_),
    .X(_02991_));
 sky130_fd_sc_hd__buf_1 _23537_ (.A(_19318_),
    .X(_19320_));
 sky130_fd_sc_hd__mux2_2 _23538_ (.A0(\cpuregs[2][27] ),
    .A1(_18304_),
    .S(_19320_),
    .X(_02990_));
 sky130_fd_sc_hd__mux2_2 _23539_ (.A0(\cpuregs[2][26] ),
    .A1(_18307_),
    .S(_19320_),
    .X(_02989_));
 sky130_fd_sc_hd__mux2_2 _23540_ (.A0(\cpuregs[2][25] ),
    .A1(_18309_),
    .S(_19320_),
    .X(_02988_));
 sky130_fd_sc_hd__mux2_2 _23541_ (.A0(\cpuregs[2][24] ),
    .A1(_18311_),
    .S(_19320_),
    .X(_02987_));
 sky130_fd_sc_hd__buf_1 _23542_ (.A(_19318_),
    .X(_19321_));
 sky130_fd_sc_hd__mux2_2 _23543_ (.A0(\cpuregs[2][23] ),
    .A1(_18313_),
    .S(_19321_),
    .X(_02986_));
 sky130_fd_sc_hd__mux2_2 _23544_ (.A0(\cpuregs[2][22] ),
    .A1(_18316_),
    .S(_19321_),
    .X(_02985_));
 sky130_fd_sc_hd__mux2_2 _23545_ (.A0(\cpuregs[2][21] ),
    .A1(_18318_),
    .S(_19321_),
    .X(_02984_));
 sky130_fd_sc_hd__mux2_2 _23546_ (.A0(\cpuregs[2][20] ),
    .A1(_18320_),
    .S(_19321_),
    .X(_02983_));
 sky130_fd_sc_hd__buf_1 _23547_ (.A(_19318_),
    .X(_19322_));
 sky130_fd_sc_hd__mux2_2 _23548_ (.A0(\cpuregs[2][19] ),
    .A1(_18322_),
    .S(_19322_),
    .X(_02982_));
 sky130_fd_sc_hd__mux2_2 _23549_ (.A0(\cpuregs[2][18] ),
    .A1(_18325_),
    .S(_19322_),
    .X(_02981_));
 sky130_fd_sc_hd__mux2_2 _23550_ (.A0(\cpuregs[2][17] ),
    .A1(_18327_),
    .S(_19322_),
    .X(_02980_));
 sky130_fd_sc_hd__mux2_2 _23551_ (.A0(\cpuregs[2][16] ),
    .A1(_18329_),
    .S(_19322_),
    .X(_02979_));
 sky130_fd_sc_hd__buf_1 _23552_ (.A(_19317_),
    .X(_19323_));
 sky130_fd_sc_hd__buf_1 _23553_ (.A(_19323_),
    .X(_19324_));
 sky130_fd_sc_hd__mux2_2 _23554_ (.A0(\cpuregs[2][15] ),
    .A1(_18331_),
    .S(_19324_),
    .X(_02978_));
 sky130_fd_sc_hd__mux2_2 _23555_ (.A0(\cpuregs[2][14] ),
    .A1(_18335_),
    .S(_19324_),
    .X(_02977_));
 sky130_fd_sc_hd__mux2_2 _23556_ (.A0(\cpuregs[2][13] ),
    .A1(_18337_),
    .S(_19324_),
    .X(_02976_));
 sky130_fd_sc_hd__mux2_2 _23557_ (.A0(\cpuregs[2][12] ),
    .A1(_18339_),
    .S(_19324_),
    .X(_02975_));
 sky130_fd_sc_hd__buf_1 _23558_ (.A(_19323_),
    .X(_19325_));
 sky130_fd_sc_hd__mux2_2 _23559_ (.A0(\cpuregs[2][11] ),
    .A1(_18341_),
    .S(_19325_),
    .X(_02974_));
 sky130_fd_sc_hd__mux2_2 _23560_ (.A0(\cpuregs[2][10] ),
    .A1(_18344_),
    .S(_19325_),
    .X(_02973_));
 sky130_fd_sc_hd__mux2_2 _23561_ (.A0(\cpuregs[2][9] ),
    .A1(_18346_),
    .S(_19325_),
    .X(_02972_));
 sky130_fd_sc_hd__mux2_2 _23562_ (.A0(\cpuregs[2][8] ),
    .A1(_18348_),
    .S(_19325_),
    .X(_02971_));
 sky130_fd_sc_hd__buf_1 _23563_ (.A(_19323_),
    .X(_19326_));
 sky130_fd_sc_hd__mux2_2 _23564_ (.A0(\cpuregs[2][7] ),
    .A1(_18350_),
    .S(_19326_),
    .X(_02970_));
 sky130_fd_sc_hd__mux2_2 _23565_ (.A0(\cpuregs[2][6] ),
    .A1(_18353_),
    .S(_19326_),
    .X(_02969_));
 sky130_fd_sc_hd__mux2_2 _23566_ (.A0(\cpuregs[2][5] ),
    .A1(_18355_),
    .S(_19326_),
    .X(_02968_));
 sky130_fd_sc_hd__mux2_2 _23567_ (.A0(\cpuregs[2][4] ),
    .A1(_18357_),
    .S(_19326_),
    .X(_02967_));
 sky130_fd_sc_hd__buf_1 _23568_ (.A(_19323_),
    .X(_19327_));
 sky130_fd_sc_hd__mux2_2 _23569_ (.A0(\cpuregs[2][3] ),
    .A1(_18359_),
    .S(_19327_),
    .X(_02966_));
 sky130_fd_sc_hd__mux2_2 _23570_ (.A0(\cpuregs[2][2] ),
    .A1(_18362_),
    .S(_19327_),
    .X(_02965_));
 sky130_fd_sc_hd__mux2_2 _23571_ (.A0(\cpuregs[2][1] ),
    .A1(_18364_),
    .S(_19327_),
    .X(_02964_));
 sky130_fd_sc_hd__mux2_2 _23572_ (.A0(\cpuregs[2][0] ),
    .A1(_18366_),
    .S(_19327_),
    .X(_02963_));
 sky130_fd_sc_hd__buf_1 _23573_ (.A(_16796_),
    .X(_19328_));
 sky130_fd_sc_hd__buf_1 _23574_ (.A(_19328_),
    .X(mem_xfer));
 sky130_fd_sc_hd__mux2_2 _23575_ (.A0(_18917_),
    .A1(mem_rdata[31]),
    .S(mem_xfer),
    .X(_02962_));
 sky130_fd_sc_hd__mux2_2 _23576_ (.A0(_18915_),
    .A1(mem_rdata[30]),
    .S(mem_xfer),
    .X(_02961_));
 sky130_fd_sc_hd__mux2_2 _23577_ (.A0(_17282_),
    .A1(mem_rdata[29]),
    .S(mem_xfer),
    .X(_02960_));
 sky130_fd_sc_hd__buf_1 _23578_ (.A(_19328_),
    .X(_19329_));
 sky130_fd_sc_hd__mux2_2 _23579_ (.A0(_18959_),
    .A1(mem_rdata[28]),
    .S(_19329_),
    .X(_02959_));
 sky130_fd_sc_hd__mux2_2 _23580_ (.A0(_18949_),
    .A1(mem_rdata[27]),
    .S(_19329_),
    .X(_02958_));
 sky130_fd_sc_hd__mux2_2 _23581_ (.A0(_18960_),
    .A1(mem_rdata[26]),
    .S(_19329_),
    .X(_02957_));
 sky130_fd_sc_hd__mux2_2 _23582_ (.A0(_18946_),
    .A1(mem_rdata[25]),
    .S(_19329_),
    .X(_02956_));
 sky130_fd_sc_hd__buf_1 _23583_ (.A(_19328_),
    .X(_19330_));
 sky130_fd_sc_hd__mux2_2 _23584_ (.A0(_18979_),
    .A1(mem_rdata[24]),
    .S(_19330_),
    .X(_02955_));
 sky130_fd_sc_hd__mux2_2 _23585_ (.A0(_19028_),
    .A1(mem_rdata[23]),
    .S(_19330_),
    .X(_02954_));
 sky130_fd_sc_hd__mux2_2 _23586_ (.A0(_19029_),
    .A1(mem_rdata[22]),
    .S(_19330_),
    .X(_02953_));
 sky130_fd_sc_hd__mux2_2 _23587_ (.A0(_19032_),
    .A1(mem_rdata[21]),
    .S(_19330_),
    .X(_02952_));
 sky130_fd_sc_hd__buf_1 _23588_ (.A(_16796_),
    .X(_19331_));
 sky130_fd_sc_hd__buf_1 _23589_ (.A(_19331_),
    .X(_19332_));
 sky130_fd_sc_hd__mux2_2 _23590_ (.A0(\mem_rdata_q[20] ),
    .A1(mem_rdata[20]),
    .S(_19332_),
    .X(_02951_));
 sky130_fd_sc_hd__mux2_2 _23591_ (.A0(\mem_rdata_q[19] ),
    .A1(mem_rdata[19]),
    .S(_19332_),
    .X(_02950_));
 sky130_fd_sc_hd__mux2_2 _23592_ (.A0(\mem_rdata_q[18] ),
    .A1(mem_rdata[18]),
    .S(_19332_),
    .X(_02949_));
 sky130_fd_sc_hd__mux2_2 _23593_ (.A0(\mem_rdata_q[17] ),
    .A1(mem_rdata[17]),
    .S(_19332_),
    .X(_02948_));
 sky130_fd_sc_hd__buf_1 _23594_ (.A(_19331_),
    .X(_19333_));
 sky130_fd_sc_hd__mux2_2 _23595_ (.A0(\mem_rdata_q[16] ),
    .A1(mem_rdata[16]),
    .S(_19333_),
    .X(_02947_));
 sky130_fd_sc_hd__mux2_2 _23596_ (.A0(\mem_rdata_q[15] ),
    .A1(mem_rdata[15]),
    .S(_19333_),
    .X(_02946_));
 sky130_fd_sc_hd__mux2_2 _23597_ (.A0(_17242_),
    .A1(mem_rdata[14]),
    .S(_19333_),
    .X(_02945_));
 sky130_fd_sc_hd__mux2_2 _23598_ (.A0(_18912_),
    .A1(mem_rdata[13]),
    .S(_19333_),
    .X(_02944_));
 sky130_fd_sc_hd__buf_1 _23599_ (.A(_19331_),
    .X(_19334_));
 sky130_fd_sc_hd__mux2_2 _23600_ (.A0(_18913_),
    .A1(mem_rdata[12]),
    .S(_19334_),
    .X(_02943_));
 sky130_fd_sc_hd__mux2_2 _23601_ (.A0(\mem_rdata_q[11] ),
    .A1(mem_rdata[11]),
    .S(_19334_),
    .X(_02942_));
 sky130_fd_sc_hd__mux2_2 _23602_ (.A0(\mem_rdata_q[10] ),
    .A1(mem_rdata[10]),
    .S(_19334_),
    .X(_02941_));
 sky130_fd_sc_hd__mux2_2 _23603_ (.A0(\mem_rdata_q[9] ),
    .A1(mem_rdata[9]),
    .S(_19334_),
    .X(_02940_));
 sky130_fd_sc_hd__buf_1 _23604_ (.A(_19331_),
    .X(_19335_));
 sky130_fd_sc_hd__mux2_2 _23605_ (.A0(\mem_rdata_q[8] ),
    .A1(mem_rdata[8]),
    .S(_19335_),
    .X(_02939_));
 sky130_fd_sc_hd__mux2_2 _23606_ (.A0(_18937_),
    .A1(mem_rdata[7]),
    .S(_19335_),
    .X(_02938_));
 sky130_fd_sc_hd__mux2_2 _23607_ (.A0(\mem_rdata_q[6] ),
    .A1(mem_rdata[6]),
    .S(_19335_),
    .X(_02937_));
 sky130_fd_sc_hd__mux2_2 _23608_ (.A0(\mem_rdata_q[5] ),
    .A1(mem_rdata[5]),
    .S(_19335_),
    .X(_02936_));
 sky130_fd_sc_hd__buf_1 _23609_ (.A(_16796_),
    .X(_19336_));
 sky130_fd_sc_hd__mux2_2 _23610_ (.A0(\mem_rdata_q[4] ),
    .A1(mem_rdata[4]),
    .S(_19336_),
    .X(_02935_));
 sky130_fd_sc_hd__mux2_2 _23611_ (.A0(\mem_rdata_q[3] ),
    .A1(mem_rdata[3]),
    .S(_19336_),
    .X(_02934_));
 sky130_fd_sc_hd__mux2_2 _23612_ (.A0(\mem_rdata_q[2] ),
    .A1(mem_rdata[2]),
    .S(_19336_),
    .X(_02933_));
 sky130_fd_sc_hd__mux2_2 _23613_ (.A0(\mem_rdata_q[1] ),
    .A1(mem_rdata[1]),
    .S(_19336_),
    .X(_02932_));
 sky130_fd_sc_hd__mux2_2 _23614_ (.A0(\mem_rdata_q[0] ),
    .A1(mem_rdata[0]),
    .S(_19328_),
    .X(_02931_));
 sky130_fd_sc_hd__o2111ai_2 _23615_ (.A1(_18890_),
    .A2(_19304_),
    .B1(_18286_),
    .C1(_18501_),
    .D1(_19305_),
    .Y(_19337_));
 sky130_fd_sc_hd__buf_1 _23616_ (.A(_19337_),
    .X(_19338_));
 sky130_fd_sc_hd__buf_1 _23617_ (.A(_19338_),
    .X(_19339_));
 sky130_fd_sc_hd__mux2_2 _23618_ (.A0(_18650_),
    .A1(\cpuregs[18][31] ),
    .S(_19339_),
    .X(_02930_));
 sky130_fd_sc_hd__mux2_2 _23619_ (.A0(_18654_),
    .A1(\cpuregs[18][30] ),
    .S(_19339_),
    .X(_02929_));
 sky130_fd_sc_hd__mux2_2 _23620_ (.A0(_18655_),
    .A1(\cpuregs[18][29] ),
    .S(_19339_),
    .X(_02928_));
 sky130_fd_sc_hd__mux2_2 _23621_ (.A0(_18656_),
    .A1(\cpuregs[18][28] ),
    .S(_19339_),
    .X(_02927_));
 sky130_fd_sc_hd__buf_1 _23622_ (.A(_19338_),
    .X(_19340_));
 sky130_fd_sc_hd__mux2_2 _23623_ (.A0(_18657_),
    .A1(\cpuregs[18][27] ),
    .S(_19340_),
    .X(_02926_));
 sky130_fd_sc_hd__mux2_2 _23624_ (.A0(_18659_),
    .A1(\cpuregs[18][26] ),
    .S(_19340_),
    .X(_02925_));
 sky130_fd_sc_hd__mux2_2 _23625_ (.A0(_18660_),
    .A1(\cpuregs[18][25] ),
    .S(_19340_),
    .X(_02924_));
 sky130_fd_sc_hd__mux2_2 _23626_ (.A0(_18661_),
    .A1(\cpuregs[18][24] ),
    .S(_19340_),
    .X(_02923_));
 sky130_fd_sc_hd__buf_1 _23627_ (.A(_19338_),
    .X(_19341_));
 sky130_fd_sc_hd__mux2_2 _23628_ (.A0(_18662_),
    .A1(\cpuregs[18][23] ),
    .S(_19341_),
    .X(_02922_));
 sky130_fd_sc_hd__mux2_2 _23629_ (.A0(_18664_),
    .A1(\cpuregs[18][22] ),
    .S(_19341_),
    .X(_02921_));
 sky130_fd_sc_hd__mux2_2 _23630_ (.A0(_18665_),
    .A1(\cpuregs[18][21] ),
    .S(_19341_),
    .X(_02920_));
 sky130_fd_sc_hd__mux2_2 _23631_ (.A0(_18666_),
    .A1(\cpuregs[18][20] ),
    .S(_19341_),
    .X(_02919_));
 sky130_fd_sc_hd__buf_1 _23632_ (.A(_19338_),
    .X(_19342_));
 sky130_fd_sc_hd__mux2_2 _23633_ (.A0(_18667_),
    .A1(\cpuregs[18][19] ),
    .S(_19342_),
    .X(_02918_));
 sky130_fd_sc_hd__mux2_2 _23634_ (.A0(_18669_),
    .A1(\cpuregs[18][18] ),
    .S(_19342_),
    .X(_02917_));
 sky130_fd_sc_hd__mux2_2 _23635_ (.A0(_18670_),
    .A1(\cpuregs[18][17] ),
    .S(_19342_),
    .X(_02916_));
 sky130_fd_sc_hd__mux2_2 _23636_ (.A0(_18671_),
    .A1(\cpuregs[18][16] ),
    .S(_19342_),
    .X(_02915_));
 sky130_fd_sc_hd__buf_1 _23637_ (.A(_19337_),
    .X(_19343_));
 sky130_fd_sc_hd__buf_1 _23638_ (.A(_19343_),
    .X(_19344_));
 sky130_fd_sc_hd__mux2_2 _23639_ (.A0(_18672_),
    .A1(\cpuregs[18][15] ),
    .S(_19344_),
    .X(_02914_));
 sky130_fd_sc_hd__mux2_2 _23640_ (.A0(_18675_),
    .A1(\cpuregs[18][14] ),
    .S(_19344_),
    .X(_02913_));
 sky130_fd_sc_hd__mux2_2 _23641_ (.A0(_18676_),
    .A1(\cpuregs[18][13] ),
    .S(_19344_),
    .X(_02912_));
 sky130_fd_sc_hd__mux2_2 _23642_ (.A0(_18677_),
    .A1(\cpuregs[18][12] ),
    .S(_19344_),
    .X(_02911_));
 sky130_fd_sc_hd__buf_1 _23643_ (.A(_19343_),
    .X(_19345_));
 sky130_fd_sc_hd__mux2_2 _23644_ (.A0(_18678_),
    .A1(\cpuregs[18][11] ),
    .S(_19345_),
    .X(_02910_));
 sky130_fd_sc_hd__mux2_2 _23645_ (.A0(_18680_),
    .A1(\cpuregs[18][10] ),
    .S(_19345_),
    .X(_02909_));
 sky130_fd_sc_hd__mux2_2 _23646_ (.A0(_18681_),
    .A1(\cpuregs[18][9] ),
    .S(_19345_),
    .X(_02908_));
 sky130_fd_sc_hd__mux2_2 _23647_ (.A0(_18682_),
    .A1(\cpuregs[18][8] ),
    .S(_19345_),
    .X(_02907_));
 sky130_fd_sc_hd__buf_1 _23648_ (.A(_19343_),
    .X(_19346_));
 sky130_fd_sc_hd__mux2_2 _23649_ (.A0(_18683_),
    .A1(\cpuregs[18][7] ),
    .S(_19346_),
    .X(_02906_));
 sky130_fd_sc_hd__mux2_2 _23650_ (.A0(_18685_),
    .A1(\cpuregs[18][6] ),
    .S(_19346_),
    .X(_02905_));
 sky130_fd_sc_hd__mux2_2 _23651_ (.A0(_18686_),
    .A1(\cpuregs[18][5] ),
    .S(_19346_),
    .X(_02904_));
 sky130_fd_sc_hd__mux2_2 _23652_ (.A0(_18687_),
    .A1(\cpuregs[18][4] ),
    .S(_19346_),
    .X(_02903_));
 sky130_fd_sc_hd__buf_1 _23653_ (.A(_19343_),
    .X(_19347_));
 sky130_fd_sc_hd__mux2_2 _23654_ (.A0(_18688_),
    .A1(\cpuregs[18][3] ),
    .S(_19347_),
    .X(_02902_));
 sky130_fd_sc_hd__mux2_2 _23655_ (.A0(_18690_),
    .A1(\cpuregs[18][2] ),
    .S(_19347_),
    .X(_02901_));
 sky130_fd_sc_hd__mux2_2 _23656_ (.A0(_18691_),
    .A1(\cpuregs[18][1] ),
    .S(_19347_),
    .X(_02900_));
 sky130_fd_sc_hd__mux2_2 _23657_ (.A0(_18692_),
    .A1(\cpuregs[18][0] ),
    .S(_19347_),
    .X(_02899_));
 sky130_fd_sc_hd__o2111ai_2 _23658_ (.A1(_18890_),
    .A2(_19304_),
    .B1(_18286_),
    .C1(_18368_),
    .D1(_19305_),
    .Y(_19348_));
 sky130_fd_sc_hd__buf_1 _23659_ (.A(_19348_),
    .X(_19349_));
 sky130_fd_sc_hd__buf_1 _23660_ (.A(_19349_),
    .X(_19350_));
 sky130_fd_sc_hd__mux2_2 _23661_ (.A0(_18456_),
    .A1(\cpuregs[10][31] ),
    .S(_19350_),
    .X(_02898_));
 sky130_fd_sc_hd__mux2_2 _23662_ (.A0(_18462_),
    .A1(\cpuregs[10][30] ),
    .S(_19350_),
    .X(_02897_));
 sky130_fd_sc_hd__mux2_2 _23663_ (.A0(_18463_),
    .A1(\cpuregs[10][29] ),
    .S(_19350_),
    .X(_02896_));
 sky130_fd_sc_hd__mux2_2 _23664_ (.A0(_18464_),
    .A1(\cpuregs[10][28] ),
    .S(_19350_),
    .X(_02895_));
 sky130_fd_sc_hd__buf_1 _23665_ (.A(_19349_),
    .X(_19351_));
 sky130_fd_sc_hd__mux2_2 _23666_ (.A0(_18465_),
    .A1(\cpuregs[10][27] ),
    .S(_19351_),
    .X(_02894_));
 sky130_fd_sc_hd__mux2_2 _23667_ (.A0(_18467_),
    .A1(\cpuregs[10][26] ),
    .S(_19351_),
    .X(_02893_));
 sky130_fd_sc_hd__mux2_2 _23668_ (.A0(_18468_),
    .A1(\cpuregs[10][25] ),
    .S(_19351_),
    .X(_02892_));
 sky130_fd_sc_hd__mux2_2 _23669_ (.A0(_18469_),
    .A1(\cpuregs[10][24] ),
    .S(_19351_),
    .X(_02891_));
 sky130_fd_sc_hd__buf_1 _23670_ (.A(_19349_),
    .X(_19352_));
 sky130_fd_sc_hd__mux2_2 _23671_ (.A0(_18470_),
    .A1(\cpuregs[10][23] ),
    .S(_19352_),
    .X(_02890_));
 sky130_fd_sc_hd__mux2_2 _23672_ (.A0(_18472_),
    .A1(\cpuregs[10][22] ),
    .S(_19352_),
    .X(_02889_));
 sky130_fd_sc_hd__mux2_2 _23673_ (.A0(_18473_),
    .A1(\cpuregs[10][21] ),
    .S(_19352_),
    .X(_02888_));
 sky130_fd_sc_hd__mux2_2 _23674_ (.A0(_18474_),
    .A1(\cpuregs[10][20] ),
    .S(_19352_),
    .X(_02887_));
 sky130_fd_sc_hd__buf_1 _23675_ (.A(_19349_),
    .X(_19353_));
 sky130_fd_sc_hd__mux2_2 _23676_ (.A0(_18475_),
    .A1(\cpuregs[10][19] ),
    .S(_19353_),
    .X(_02886_));
 sky130_fd_sc_hd__mux2_2 _23677_ (.A0(_18477_),
    .A1(\cpuregs[10][18] ),
    .S(_19353_),
    .X(_02885_));
 sky130_fd_sc_hd__mux2_2 _23678_ (.A0(_18478_),
    .A1(\cpuregs[10][17] ),
    .S(_19353_),
    .X(_02884_));
 sky130_fd_sc_hd__mux2_2 _23679_ (.A0(_18479_),
    .A1(\cpuregs[10][16] ),
    .S(_19353_),
    .X(_02883_));
 sky130_fd_sc_hd__buf_1 _23680_ (.A(_19348_),
    .X(_19354_));
 sky130_fd_sc_hd__buf_1 _23681_ (.A(_19354_),
    .X(_19355_));
 sky130_fd_sc_hd__mux2_2 _23682_ (.A0(_18480_),
    .A1(\cpuregs[10][15] ),
    .S(_19355_),
    .X(_02882_));
 sky130_fd_sc_hd__mux2_2 _23683_ (.A0(_18483_),
    .A1(\cpuregs[10][14] ),
    .S(_19355_),
    .X(_02881_));
 sky130_fd_sc_hd__mux2_2 _23684_ (.A0(_18484_),
    .A1(\cpuregs[10][13] ),
    .S(_19355_),
    .X(_02880_));
 sky130_fd_sc_hd__mux2_2 _23685_ (.A0(_18485_),
    .A1(\cpuregs[10][12] ),
    .S(_19355_),
    .X(_02879_));
 sky130_fd_sc_hd__buf_1 _23686_ (.A(_19354_),
    .X(_19356_));
 sky130_fd_sc_hd__mux2_2 _23687_ (.A0(_18486_),
    .A1(\cpuregs[10][11] ),
    .S(_19356_),
    .X(_02878_));
 sky130_fd_sc_hd__mux2_2 _23688_ (.A0(_18488_),
    .A1(\cpuregs[10][10] ),
    .S(_19356_),
    .X(_02877_));
 sky130_fd_sc_hd__mux2_2 _23689_ (.A0(_18489_),
    .A1(\cpuregs[10][9] ),
    .S(_19356_),
    .X(_02876_));
 sky130_fd_sc_hd__mux2_2 _23690_ (.A0(_18490_),
    .A1(\cpuregs[10][8] ),
    .S(_19356_),
    .X(_02875_));
 sky130_fd_sc_hd__buf_1 _23691_ (.A(_19354_),
    .X(_19357_));
 sky130_fd_sc_hd__mux2_2 _23692_ (.A0(_18491_),
    .A1(\cpuregs[10][7] ),
    .S(_19357_),
    .X(_02874_));
 sky130_fd_sc_hd__mux2_2 _23693_ (.A0(_18493_),
    .A1(\cpuregs[10][6] ),
    .S(_19357_),
    .X(_02873_));
 sky130_fd_sc_hd__mux2_2 _23694_ (.A0(_18494_),
    .A1(\cpuregs[10][5] ),
    .S(_19357_),
    .X(_02872_));
 sky130_fd_sc_hd__mux2_2 _23695_ (.A0(_18495_),
    .A1(\cpuregs[10][4] ),
    .S(_19357_),
    .X(_02871_));
 sky130_fd_sc_hd__buf_1 _23696_ (.A(_19354_),
    .X(_19358_));
 sky130_fd_sc_hd__mux2_2 _23697_ (.A0(_18496_),
    .A1(\cpuregs[10][3] ),
    .S(_19358_),
    .X(_02870_));
 sky130_fd_sc_hd__mux2_2 _23698_ (.A0(_18498_),
    .A1(\cpuregs[10][2] ),
    .S(_19358_),
    .X(_02869_));
 sky130_fd_sc_hd__mux2_2 _23699_ (.A0(_18499_),
    .A1(\cpuregs[10][1] ),
    .S(_19358_),
    .X(_02868_));
 sky130_fd_sc_hd__mux2_2 _23700_ (.A0(_18500_),
    .A1(\cpuregs[10][0] ),
    .S(_19358_),
    .X(_02867_));
 sky130_fd_sc_hd__buf_1 _23701_ (.A(\cpuregs[0][31] ),
    .X(_02866_));
 sky130_fd_sc_hd__buf_1 _23702_ (.A(\cpuregs[0][30] ),
    .X(_02865_));
 sky130_fd_sc_hd__buf_1 _23703_ (.A(\cpuregs[0][29] ),
    .X(_02864_));
 sky130_fd_sc_hd__buf_1 _23704_ (.A(\cpuregs[0][28] ),
    .X(_02863_));
 sky130_fd_sc_hd__buf_1 _23705_ (.A(\cpuregs[0][27] ),
    .X(_02862_));
 sky130_fd_sc_hd__buf_1 _23706_ (.A(\cpuregs[0][26] ),
    .X(_02861_));
 sky130_fd_sc_hd__buf_1 _23707_ (.A(\cpuregs[0][25] ),
    .X(_02860_));
 sky130_fd_sc_hd__buf_1 _23708_ (.A(\cpuregs[0][24] ),
    .X(_02859_));
 sky130_fd_sc_hd__buf_1 _23709_ (.A(\cpuregs[0][23] ),
    .X(_02858_));
 sky130_fd_sc_hd__buf_1 _23710_ (.A(\cpuregs[0][22] ),
    .X(_02857_));
 sky130_fd_sc_hd__buf_1 _23711_ (.A(\cpuregs[0][21] ),
    .X(_02856_));
 sky130_fd_sc_hd__buf_1 _23712_ (.A(\cpuregs[0][20] ),
    .X(_02855_));
 sky130_fd_sc_hd__buf_1 _23713_ (.A(\cpuregs[0][19] ),
    .X(_02854_));
 sky130_fd_sc_hd__buf_1 _23714_ (.A(\cpuregs[0][18] ),
    .X(_02853_));
 sky130_fd_sc_hd__buf_1 _23715_ (.A(\cpuregs[0][17] ),
    .X(_02852_));
 sky130_fd_sc_hd__buf_1 _23716_ (.A(\cpuregs[0][16] ),
    .X(_02851_));
 sky130_fd_sc_hd__buf_1 _23717_ (.A(\cpuregs[0][15] ),
    .X(_02850_));
 sky130_fd_sc_hd__buf_1 _23718_ (.A(\cpuregs[0][14] ),
    .X(_02849_));
 sky130_fd_sc_hd__buf_1 _23719_ (.A(\cpuregs[0][13] ),
    .X(_02848_));
 sky130_fd_sc_hd__buf_1 _23720_ (.A(\cpuregs[0][12] ),
    .X(_02847_));
 sky130_fd_sc_hd__buf_1 _23721_ (.A(\cpuregs[0][11] ),
    .X(_02846_));
 sky130_fd_sc_hd__buf_1 _23722_ (.A(\cpuregs[0][10] ),
    .X(_02845_));
 sky130_fd_sc_hd__buf_1 _23723_ (.A(\cpuregs[0][9] ),
    .X(_02844_));
 sky130_fd_sc_hd__buf_1 _23724_ (.A(\cpuregs[0][8] ),
    .X(_02843_));
 sky130_fd_sc_hd__buf_1 _23725_ (.A(\cpuregs[0][7] ),
    .X(_02842_));
 sky130_fd_sc_hd__buf_1 _23726_ (.A(\cpuregs[0][6] ),
    .X(_02841_));
 sky130_fd_sc_hd__buf_1 _23727_ (.A(\cpuregs[0][5] ),
    .X(_02840_));
 sky130_fd_sc_hd__buf_1 _23728_ (.A(\cpuregs[0][4] ),
    .X(_02839_));
 sky130_fd_sc_hd__buf_1 _23729_ (.A(\cpuregs[0][3] ),
    .X(_02838_));
 sky130_fd_sc_hd__buf_1 _23730_ (.A(\cpuregs[0][2] ),
    .X(_02837_));
 sky130_fd_sc_hd__buf_1 _23731_ (.A(\cpuregs[0][1] ),
    .X(_02836_));
 sky130_fd_sc_hd__buf_1 _23732_ (.A(\cpuregs[0][0] ),
    .X(_02835_));
 sky130_fd_sc_hd__o2111ai_2 _23733_ (.A1(_18626_),
    .A2(_19304_),
    .B1(_18286_),
    .C1(_18549_),
    .D1(_19305_),
    .Y(_19359_));
 sky130_fd_sc_hd__buf_1 _23734_ (.A(_19359_),
    .X(_19360_));
 sky130_fd_sc_hd__buf_1 _23735_ (.A(_19360_),
    .X(_19361_));
 sky130_fd_sc_hd__mux2_2 _23736_ (.A0(_18456_),
    .A1(\cpuregs[14][31] ),
    .S(_19361_),
    .X(_02834_));
 sky130_fd_sc_hd__mux2_2 _23737_ (.A0(_18462_),
    .A1(\cpuregs[14][30] ),
    .S(_19361_),
    .X(_02833_));
 sky130_fd_sc_hd__mux2_2 _23738_ (.A0(_18463_),
    .A1(\cpuregs[14][29] ),
    .S(_19361_),
    .X(_02832_));
 sky130_fd_sc_hd__mux2_2 _23739_ (.A0(_18464_),
    .A1(\cpuregs[14][28] ),
    .S(_19361_),
    .X(_02831_));
 sky130_fd_sc_hd__buf_1 _23740_ (.A(_19360_),
    .X(_19362_));
 sky130_fd_sc_hd__mux2_2 _23741_ (.A0(_18465_),
    .A1(\cpuregs[14][27] ),
    .S(_19362_),
    .X(_02830_));
 sky130_fd_sc_hd__mux2_2 _23742_ (.A0(_18467_),
    .A1(\cpuregs[14][26] ),
    .S(_19362_),
    .X(_02829_));
 sky130_fd_sc_hd__mux2_2 _23743_ (.A0(_18468_),
    .A1(\cpuregs[14][25] ),
    .S(_19362_),
    .X(_02828_));
 sky130_fd_sc_hd__mux2_2 _23744_ (.A0(_18469_),
    .A1(\cpuregs[14][24] ),
    .S(_19362_),
    .X(_02827_));
 sky130_fd_sc_hd__buf_1 _23745_ (.A(_19360_),
    .X(_19363_));
 sky130_fd_sc_hd__mux2_2 _23746_ (.A0(_18470_),
    .A1(\cpuregs[14][23] ),
    .S(_19363_),
    .X(_02826_));
 sky130_fd_sc_hd__mux2_2 _23747_ (.A0(_18472_),
    .A1(\cpuregs[14][22] ),
    .S(_19363_),
    .X(_02825_));
 sky130_fd_sc_hd__mux2_2 _23748_ (.A0(_18473_),
    .A1(\cpuregs[14][21] ),
    .S(_19363_),
    .X(_02824_));
 sky130_fd_sc_hd__mux2_2 _23749_ (.A0(_18474_),
    .A1(\cpuregs[14][20] ),
    .S(_19363_),
    .X(_02823_));
 sky130_fd_sc_hd__buf_1 _23750_ (.A(_19360_),
    .X(_19364_));
 sky130_fd_sc_hd__mux2_2 _23751_ (.A0(_18475_),
    .A1(\cpuregs[14][19] ),
    .S(_19364_),
    .X(_02822_));
 sky130_fd_sc_hd__mux2_2 _23752_ (.A0(_18477_),
    .A1(\cpuregs[14][18] ),
    .S(_19364_),
    .X(_02821_));
 sky130_fd_sc_hd__mux2_2 _23753_ (.A0(_18478_),
    .A1(\cpuregs[14][17] ),
    .S(_19364_),
    .X(_02820_));
 sky130_fd_sc_hd__mux2_2 _23754_ (.A0(_18479_),
    .A1(\cpuregs[14][16] ),
    .S(_19364_),
    .X(_02819_));
 sky130_fd_sc_hd__buf_1 _23755_ (.A(_19359_),
    .X(_19365_));
 sky130_fd_sc_hd__buf_1 _23756_ (.A(_19365_),
    .X(_19366_));
 sky130_fd_sc_hd__mux2_2 _23757_ (.A0(_18480_),
    .A1(\cpuregs[14][15] ),
    .S(_19366_),
    .X(_02818_));
 sky130_fd_sc_hd__mux2_2 _23758_ (.A0(_18483_),
    .A1(\cpuregs[14][14] ),
    .S(_19366_),
    .X(_02817_));
 sky130_fd_sc_hd__mux2_2 _23759_ (.A0(_18484_),
    .A1(\cpuregs[14][13] ),
    .S(_19366_),
    .X(_02816_));
 sky130_fd_sc_hd__mux2_2 _23760_ (.A0(_18485_),
    .A1(\cpuregs[14][12] ),
    .S(_19366_),
    .X(_02815_));
 sky130_fd_sc_hd__buf_1 _23761_ (.A(_19365_),
    .X(_19367_));
 sky130_fd_sc_hd__mux2_2 _23762_ (.A0(_18486_),
    .A1(\cpuregs[14][11] ),
    .S(_19367_),
    .X(_02814_));
 sky130_fd_sc_hd__mux2_2 _23763_ (.A0(_18488_),
    .A1(\cpuregs[14][10] ),
    .S(_19367_),
    .X(_02813_));
 sky130_fd_sc_hd__mux2_2 _23764_ (.A0(_18489_),
    .A1(\cpuregs[14][9] ),
    .S(_19367_),
    .X(_02812_));
 sky130_fd_sc_hd__mux2_2 _23765_ (.A0(_18490_),
    .A1(\cpuregs[14][8] ),
    .S(_19367_),
    .X(_02811_));
 sky130_fd_sc_hd__buf_1 _23766_ (.A(_19365_),
    .X(_19368_));
 sky130_fd_sc_hd__mux2_2 _23767_ (.A0(_18491_),
    .A1(\cpuregs[14][7] ),
    .S(_19368_),
    .X(_02810_));
 sky130_fd_sc_hd__mux2_2 _23768_ (.A0(_18493_),
    .A1(\cpuregs[14][6] ),
    .S(_19368_),
    .X(_02809_));
 sky130_fd_sc_hd__mux2_2 _23769_ (.A0(_18494_),
    .A1(\cpuregs[14][5] ),
    .S(_19368_),
    .X(_02808_));
 sky130_fd_sc_hd__mux2_2 _23770_ (.A0(_18495_),
    .A1(\cpuregs[14][4] ),
    .S(_19368_),
    .X(_02807_));
 sky130_fd_sc_hd__buf_1 _23771_ (.A(_19365_),
    .X(_19369_));
 sky130_fd_sc_hd__mux2_2 _23772_ (.A0(_18496_),
    .A1(\cpuregs[14][3] ),
    .S(_19369_),
    .X(_02806_));
 sky130_fd_sc_hd__mux2_2 _23773_ (.A0(_18498_),
    .A1(\cpuregs[14][2] ),
    .S(_19369_),
    .X(_02805_));
 sky130_fd_sc_hd__mux2_2 _23774_ (.A0(_18499_),
    .A1(\cpuregs[14][1] ),
    .S(_19369_),
    .X(_02804_));
 sky130_fd_sc_hd__mux2_2 _23775_ (.A0(_18500_),
    .A1(\cpuregs[14][0] ),
    .S(_19369_),
    .X(_02803_));
 sky130_fd_sc_hd__nand3b_2 _23776_ (.A_N(_18626_),
    .B(_18458_),
    .C(_18368_),
    .Y(_19370_));
 sky130_fd_sc_hd__buf_1 _23777_ (.A(_19370_),
    .X(_19371_));
 sky130_fd_sc_hd__buf_1 _23778_ (.A(_19371_),
    .X(_19372_));
 sky130_fd_sc_hd__mux2_2 _23779_ (.A0(_18456_),
    .A1(\cpuregs[8][31] ),
    .S(_19372_),
    .X(_02802_));
 sky130_fd_sc_hd__mux2_2 _23780_ (.A0(_18462_),
    .A1(\cpuregs[8][30] ),
    .S(_19372_),
    .X(_02801_));
 sky130_fd_sc_hd__mux2_2 _23781_ (.A0(_18463_),
    .A1(\cpuregs[8][29] ),
    .S(_19372_),
    .X(_02800_));
 sky130_fd_sc_hd__mux2_2 _23782_ (.A0(_18464_),
    .A1(\cpuregs[8][28] ),
    .S(_19372_),
    .X(_02799_));
 sky130_fd_sc_hd__buf_1 _23783_ (.A(_19371_),
    .X(_19373_));
 sky130_fd_sc_hd__mux2_2 _23784_ (.A0(_18465_),
    .A1(\cpuregs[8][27] ),
    .S(_19373_),
    .X(_02798_));
 sky130_fd_sc_hd__mux2_2 _23785_ (.A0(_18467_),
    .A1(\cpuregs[8][26] ),
    .S(_19373_),
    .X(_02797_));
 sky130_fd_sc_hd__mux2_2 _23786_ (.A0(_18468_),
    .A1(\cpuregs[8][25] ),
    .S(_19373_),
    .X(_02796_));
 sky130_fd_sc_hd__mux2_2 _23787_ (.A0(_18469_),
    .A1(\cpuregs[8][24] ),
    .S(_19373_),
    .X(_02795_));
 sky130_fd_sc_hd__buf_1 _23788_ (.A(_19371_),
    .X(_19374_));
 sky130_fd_sc_hd__mux2_2 _23789_ (.A0(_18470_),
    .A1(\cpuregs[8][23] ),
    .S(_19374_),
    .X(_02794_));
 sky130_fd_sc_hd__mux2_2 _23790_ (.A0(_18472_),
    .A1(\cpuregs[8][22] ),
    .S(_19374_),
    .X(_02793_));
 sky130_fd_sc_hd__mux2_2 _23791_ (.A0(_18473_),
    .A1(\cpuregs[8][21] ),
    .S(_19374_),
    .X(_02792_));
 sky130_fd_sc_hd__mux2_2 _23792_ (.A0(_18474_),
    .A1(\cpuregs[8][20] ),
    .S(_19374_),
    .X(_02791_));
 sky130_fd_sc_hd__buf_1 _23793_ (.A(_19371_),
    .X(_19375_));
 sky130_fd_sc_hd__mux2_2 _23794_ (.A0(_18475_),
    .A1(\cpuregs[8][19] ),
    .S(_19375_),
    .X(_02790_));
 sky130_fd_sc_hd__mux2_2 _23795_ (.A0(_18477_),
    .A1(\cpuregs[8][18] ),
    .S(_19375_),
    .X(_02789_));
 sky130_fd_sc_hd__mux2_2 _23796_ (.A0(_18478_),
    .A1(\cpuregs[8][17] ),
    .S(_19375_),
    .X(_02788_));
 sky130_fd_sc_hd__mux2_2 _23797_ (.A0(_18479_),
    .A1(\cpuregs[8][16] ),
    .S(_19375_),
    .X(_02787_));
 sky130_fd_sc_hd__buf_1 _23798_ (.A(_19370_),
    .X(_19376_));
 sky130_fd_sc_hd__buf_1 _23799_ (.A(_19376_),
    .X(_19377_));
 sky130_fd_sc_hd__mux2_2 _23800_ (.A0(_18480_),
    .A1(\cpuregs[8][15] ),
    .S(_19377_),
    .X(_02786_));
 sky130_fd_sc_hd__mux2_2 _23801_ (.A0(_18483_),
    .A1(\cpuregs[8][14] ),
    .S(_19377_),
    .X(_02785_));
 sky130_fd_sc_hd__mux2_2 _23802_ (.A0(_18484_),
    .A1(\cpuregs[8][13] ),
    .S(_19377_),
    .X(_02784_));
 sky130_fd_sc_hd__mux2_2 _23803_ (.A0(_18485_),
    .A1(\cpuregs[8][12] ),
    .S(_19377_),
    .X(_02783_));
 sky130_fd_sc_hd__buf_1 _23804_ (.A(_19376_),
    .X(_19378_));
 sky130_fd_sc_hd__mux2_2 _23805_ (.A0(_18486_),
    .A1(\cpuregs[8][11] ),
    .S(_19378_),
    .X(_02782_));
 sky130_fd_sc_hd__mux2_2 _23806_ (.A0(_18488_),
    .A1(\cpuregs[8][10] ),
    .S(_19378_),
    .X(_02781_));
 sky130_fd_sc_hd__mux2_2 _23807_ (.A0(_18489_),
    .A1(\cpuregs[8][9] ),
    .S(_19378_),
    .X(_02780_));
 sky130_fd_sc_hd__mux2_2 _23808_ (.A0(_18490_),
    .A1(\cpuregs[8][8] ),
    .S(_19378_),
    .X(_02779_));
 sky130_fd_sc_hd__buf_1 _23809_ (.A(_19376_),
    .X(_19379_));
 sky130_fd_sc_hd__mux2_2 _23810_ (.A0(_18491_),
    .A1(\cpuregs[8][7] ),
    .S(_19379_),
    .X(_02778_));
 sky130_fd_sc_hd__mux2_2 _23811_ (.A0(_18493_),
    .A1(\cpuregs[8][6] ),
    .S(_19379_),
    .X(_02777_));
 sky130_fd_sc_hd__mux2_2 _23812_ (.A0(_18494_),
    .A1(\cpuregs[8][5] ),
    .S(_19379_),
    .X(_02776_));
 sky130_fd_sc_hd__mux2_2 _23813_ (.A0(_18495_),
    .A1(\cpuregs[8][4] ),
    .S(_19379_),
    .X(_02775_));
 sky130_fd_sc_hd__buf_1 _23814_ (.A(_19376_),
    .X(_19380_));
 sky130_fd_sc_hd__mux2_2 _23815_ (.A0(_18496_),
    .A1(\cpuregs[8][3] ),
    .S(_19380_),
    .X(_02774_));
 sky130_fd_sc_hd__mux2_2 _23816_ (.A0(_18498_),
    .A1(\cpuregs[8][2] ),
    .S(_19380_),
    .X(_02773_));
 sky130_fd_sc_hd__mux2_2 _23817_ (.A0(_18499_),
    .A1(\cpuregs[8][1] ),
    .S(_19380_),
    .X(_02772_));
 sky130_fd_sc_hd__mux2_2 _23818_ (.A0(_18500_),
    .A1(\cpuregs[8][0] ),
    .S(_19380_),
    .X(_02771_));
 sky130_fd_sc_hd__nor2_2 _23819_ (.A(_16833_),
    .B(_17037_),
    .Y(_00292_));
 sky130_fd_sc_hd__and2b_2 _23820_ (.A_N(_16987_),
    .B(_16833_),
    .X(_19381_));
 sky130_fd_sc_hd__buf_1 _23821_ (.A(\reg_next_pc[0] ),
    .X(_19382_));
 sky130_fd_sc_hd__o311a_2 _23822_ (.A1(_17392_),
    .A2(_00292_),
    .A3(_19381_),
    .B1(_16832_),
    .C1(_19382_),
    .X(_02770_));
 sky130_fd_sc_hd__and2_2 _23823_ (.A(_18271_),
    .B(_00008_),
    .X(_02769_));
 sky130_fd_sc_hd__and2_2 _23824_ (.A(_18271_),
    .B(_19818_),
    .X(_02768_));
 sky130_fd_sc_hd__and2_2 _23825_ (.A(_18271_),
    .B(_00031_),
    .X(_02767_));
 sky130_fd_sc_hd__buf_1 _23826_ (.A(_18038_),
    .X(_19383_));
 sky130_fd_sc_hd__and2_2 _23827_ (.A(_19383_),
    .B(_00032_),
    .X(_02766_));
 sky130_fd_sc_hd__and2_2 _23828_ (.A(_19383_),
    .B(_00033_),
    .X(_02765_));
 sky130_fd_sc_hd__and2_2 _23829_ (.A(_19383_),
    .B(_00034_),
    .X(_02764_));
 sky130_fd_sc_hd__and2_2 _23830_ (.A(_19383_),
    .B(_00035_),
    .X(_02763_));
 sky130_fd_sc_hd__buf_1 _23831_ (.A(_17324_),
    .X(_19384_));
 sky130_fd_sc_hd__buf_1 _23832_ (.A(_19384_),
    .X(_19385_));
 sky130_fd_sc_hd__and2_2 _23833_ (.A(_19385_),
    .B(_00036_),
    .X(_02762_));
 sky130_fd_sc_hd__and2_2 _23834_ (.A(_19385_),
    .B(_00037_),
    .X(_02761_));
 sky130_fd_sc_hd__and2_2 _23835_ (.A(_19385_),
    .B(_00009_),
    .X(_02760_));
 sky130_fd_sc_hd__and2_2 _23836_ (.A(_19385_),
    .B(_00010_),
    .X(_02759_));
 sky130_fd_sc_hd__buf_1 _23837_ (.A(_19384_),
    .X(_19386_));
 sky130_fd_sc_hd__and2_2 _23838_ (.A(_19386_),
    .B(_00011_),
    .X(_02758_));
 sky130_fd_sc_hd__and2_2 _23839_ (.A(_19386_),
    .B(_00012_),
    .X(_02757_));
 sky130_fd_sc_hd__and2_2 _23840_ (.A(_19386_),
    .B(_00013_),
    .X(_02756_));
 sky130_fd_sc_hd__and2_2 _23841_ (.A(_19386_),
    .B(_00014_),
    .X(_02755_));
 sky130_fd_sc_hd__buf_1 _23842_ (.A(_19384_),
    .X(_19387_));
 sky130_fd_sc_hd__and2_2 _23843_ (.A(_19387_),
    .B(_00015_),
    .X(_02754_));
 sky130_fd_sc_hd__and2_2 _23844_ (.A(_19387_),
    .B(_00016_),
    .X(_02753_));
 sky130_fd_sc_hd__and2_2 _23845_ (.A(_19387_),
    .B(_00017_),
    .X(_02752_));
 sky130_fd_sc_hd__and2_2 _23846_ (.A(_19387_),
    .B(_00018_),
    .X(_02751_));
 sky130_fd_sc_hd__buf_1 _23847_ (.A(_19384_),
    .X(_19388_));
 sky130_fd_sc_hd__and2_2 _23848_ (.A(_19388_),
    .B(_00019_),
    .X(_02750_));
 sky130_fd_sc_hd__and2_2 _23849_ (.A(_19388_),
    .B(_00020_),
    .X(_02749_));
 sky130_fd_sc_hd__and2_2 _23850_ (.A(_19388_),
    .B(_00021_),
    .X(_02748_));
 sky130_fd_sc_hd__and2_2 _23851_ (.A(_19388_),
    .B(_00022_),
    .X(_02747_));
 sky130_fd_sc_hd__buf_1 _23852_ (.A(_16831_),
    .X(_19389_));
 sky130_fd_sc_hd__and2_2 _23853_ (.A(_19389_),
    .B(_00023_),
    .X(_02746_));
 sky130_fd_sc_hd__and2_2 _23854_ (.A(_19389_),
    .B(_00024_),
    .X(_02745_));
 sky130_fd_sc_hd__and2_2 _23855_ (.A(_19389_),
    .B(_00025_),
    .X(_02744_));
 sky130_fd_sc_hd__and2_2 _23856_ (.A(_19389_),
    .B(_00026_),
    .X(_02743_));
 sky130_fd_sc_hd__buf_1 _23857_ (.A(_16831_),
    .X(_19390_));
 sky130_fd_sc_hd__and2_2 _23858_ (.A(_19390_),
    .B(_00027_),
    .X(_02742_));
 sky130_fd_sc_hd__and2_2 _23859_ (.A(_19390_),
    .B(_00028_),
    .X(_02741_));
 sky130_fd_sc_hd__and2_2 _23860_ (.A(_19390_),
    .B(_00029_),
    .X(_02740_));
 sky130_fd_sc_hd__and2_2 _23861_ (.A(_19390_),
    .B(_00030_),
    .X(_02739_));
 sky130_fd_sc_hd__nor2_2 _23862_ (.A(_16980_),
    .B(is_sb_sh_sw),
    .Y(_19391_));
 sky130_vsdinv _23863_ (.A(_19391_),
    .Y(_19392_));
 sky130_vsdinv _23864_ (.A(_18939_),
    .Y(_19393_));
 sky130_fd_sc_hd__buf_1 _23865_ (.A(_17082_),
    .X(_19394_));
 sky130_fd_sc_hd__and2_2 _23866_ (.A(_18935_),
    .B(_19394_),
    .X(_19395_));
 sky130_fd_sc_hd__a221o_2 _23867_ (.A1(\mem_rdata_q[8] ),
    .A2(_19392_),
    .B1(_19393_),
    .B2(_19032_),
    .C1(_19395_),
    .X(_19396_));
 sky130_fd_sc_hd__buf_1 _23868_ (.A(\decoded_imm[1] ),
    .X(_19397_));
 sky130_fd_sc_hd__mux2_2 _23869_ (.A0(_19396_),
    .A1(_19397_),
    .S(_18910_),
    .X(_02738_));
 sky130_fd_sc_hd__and2_2 _23870_ (.A(\decoded_imm_uj[2] ),
    .B(_19394_),
    .X(_19398_));
 sky130_fd_sc_hd__a221o_2 _23871_ (.A1(\mem_rdata_q[9] ),
    .A2(_19392_),
    .B1(_19393_),
    .B2(_19029_),
    .C1(_19398_),
    .X(_19399_));
 sky130_fd_sc_hd__buf_1 _23872_ (.A(\decoded_imm[2] ),
    .X(_19400_));
 sky130_fd_sc_hd__buf_1 _23873_ (.A(_17341_),
    .X(_19401_));
 sky130_fd_sc_hd__mux2_2 _23874_ (.A0(_19399_),
    .A1(_19400_),
    .S(_19401_),
    .X(_02737_));
 sky130_fd_sc_hd__and2_2 _23875_ (.A(_18934_),
    .B(_19394_),
    .X(_19402_));
 sky130_fd_sc_hd__a221o_2 _23876_ (.A1(\mem_rdata_q[10] ),
    .A2(_19392_),
    .B1(_19393_),
    .B2(_19028_),
    .C1(_19402_),
    .X(_19403_));
 sky130_fd_sc_hd__buf_1 _23877_ (.A(\decoded_imm[3] ),
    .X(_19404_));
 sky130_fd_sc_hd__mux2_2 _23878_ (.A0(_19403_),
    .A1(_19404_),
    .S(_19401_),
    .X(_02736_));
 sky130_fd_sc_hd__and2_2 _23879_ (.A(_18932_),
    .B(_19394_),
    .X(_19405_));
 sky130_fd_sc_hd__a221o_2 _23880_ (.A1(\mem_rdata_q[11] ),
    .A2(_19392_),
    .B1(_19393_),
    .B2(_18979_),
    .C1(_19405_),
    .X(_19406_));
 sky130_fd_sc_hd__buf_1 _23881_ (.A(\decoded_imm[4] ),
    .X(_19407_));
 sky130_fd_sc_hd__mux2_2 _23882_ (.A0(_19406_),
    .A1(_19407_),
    .S(_19401_),
    .X(_02735_));
 sky130_fd_sc_hd__nand3_2 _23883_ (.A(_18939_),
    .B(_18542_),
    .C(_17061_),
    .Y(_19408_));
 sky130_fd_sc_hd__buf_1 _23884_ (.A(_19408_),
    .X(_19409_));
 sky130_fd_sc_hd__buf_1 _23885_ (.A(_19409_),
    .X(_19410_));
 sky130_vsdinv _23886_ (.A(\decoded_imm_uj[5] ),
    .Y(_19411_));
 sky130_fd_sc_hd__o2bb2ai_2 _23887_ (.A1_N(_18946_),
    .A2_N(_19410_),
    .B1(_19411_),
    .B2(_00323_),
    .Y(_19412_));
 sky130_fd_sc_hd__buf_1 _23888_ (.A(\decoded_imm[5] ),
    .X(_19413_));
 sky130_fd_sc_hd__mux2_2 _23889_ (.A0(_19412_),
    .A1(_19413_),
    .S(_19401_),
    .X(_02734_));
 sky130_fd_sc_hd__a22o_2 _23890_ (.A1(\decoded_imm_uj[6] ),
    .A2(_17084_),
    .B1(_19410_),
    .B2(_18960_),
    .X(_19414_));
 sky130_fd_sc_hd__buf_1 _23891_ (.A(\decoded_imm[6] ),
    .X(_19415_));
 sky130_fd_sc_hd__buf_1 _23892_ (.A(_18972_),
    .X(_19416_));
 sky130_fd_sc_hd__mux2_2 _23893_ (.A0(_19414_),
    .A1(_19415_),
    .S(_19416_),
    .X(_02733_));
 sky130_vsdinv _23894_ (.A(\decoded_imm_uj[7] ),
    .Y(_19417_));
 sky130_fd_sc_hd__o2bb2ai_2 _23895_ (.A1_N(_18949_),
    .A2_N(_19410_),
    .B1(_19417_),
    .B2(_00323_),
    .Y(_19418_));
 sky130_fd_sc_hd__buf_1 _23896_ (.A(\decoded_imm[7] ),
    .X(_19419_));
 sky130_fd_sc_hd__mux2_2 _23897_ (.A0(_19418_),
    .A1(_19419_),
    .S(_19416_),
    .X(_02732_));
 sky130_fd_sc_hd__buf_1 _23898_ (.A(_19408_),
    .X(_19420_));
 sky130_fd_sc_hd__a22o_2 _23899_ (.A1(_18930_),
    .A2(_17084_),
    .B1(_19420_),
    .B2(\mem_rdata_q[28] ),
    .X(_19421_));
 sky130_fd_sc_hd__buf_1 _23900_ (.A(\decoded_imm[8] ),
    .X(_19422_));
 sky130_fd_sc_hd__mux2_2 _23901_ (.A0(_19421_),
    .A1(_19422_),
    .S(_19416_),
    .X(_02731_));
 sky130_vsdinv _23902_ (.A(\decoded_imm_uj[9] ),
    .Y(_19423_));
 sky130_fd_sc_hd__o2bb2ai_2 _23903_ (.A1_N(_17282_),
    .A2_N(_19410_),
    .B1(_19423_),
    .B2(_16989_),
    .Y(_19424_));
 sky130_fd_sc_hd__buf_1 _23904_ (.A(\decoded_imm[9] ),
    .X(_19425_));
 sky130_fd_sc_hd__mux2_2 _23905_ (.A0(_19424_),
    .A1(_19425_),
    .S(_19416_),
    .X(_02730_));
 sky130_fd_sc_hd__a22o_2 _23906_ (.A1(_18929_),
    .A2(_17083_),
    .B1(_19420_),
    .B2(_18915_),
    .X(_19426_));
 sky130_fd_sc_hd__buf_1 _23907_ (.A(\decoded_imm[10] ),
    .X(_19427_));
 sky130_fd_sc_hd__buf_1 _23908_ (.A(_18972_),
    .X(_19428_));
 sky130_fd_sc_hd__mux2_2 _23909_ (.A0(_19426_),
    .A1(_19427_),
    .S(_19428_),
    .X(_02729_));
 sky130_fd_sc_hd__buf_1 _23910_ (.A(\decoded_imm[11] ),
    .X(_19429_));
 sky130_fd_sc_hd__nand2_2 _23911_ (.A(_18939_),
    .B(_17062_),
    .Y(_19430_));
 sky130_fd_sc_hd__and2_2 _23912_ (.A(_16980_),
    .B(_18937_),
    .X(_19431_));
 sky130_fd_sc_hd__a221oi_2 _23913_ (.A1(\decoded_imm_uj[11] ),
    .A2(_17084_),
    .B1(_19430_),
    .B2(_18917_),
    .C1(_19431_),
    .Y(_19432_));
 sky130_fd_sc_hd__nor2_2 _23914_ (.A(_17342_),
    .B(_19432_),
    .Y(_19433_));
 sky130_fd_sc_hd__a21o_2 _23915_ (.A1(_19429_),
    .A2(_18955_),
    .B1(_19433_),
    .X(_02728_));
 sky130_vsdinv _23916_ (.A(_16988_),
    .Y(_19434_));
 sky130_fd_sc_hd__buf_1 _23917_ (.A(_19434_),
    .X(_19435_));
 sky130_fd_sc_hd__buf_1 _23918_ (.A(_18916_),
    .X(_19436_));
 sky130_fd_sc_hd__buf_1 _23919_ (.A(_17082_),
    .X(_19437_));
 sky130_fd_sc_hd__and2_2 _23920_ (.A(\decoded_imm_uj[12] ),
    .B(_19437_),
    .X(_19438_));
 sky130_fd_sc_hd__a221o_2 _23921_ (.A1(_18913_),
    .A2(_19435_),
    .B1(_19420_),
    .B2(_19436_),
    .C1(_19438_),
    .X(_19439_));
 sky130_fd_sc_hd__buf_1 _23922_ (.A(\decoded_imm[12] ),
    .X(_19440_));
 sky130_fd_sc_hd__mux2_2 _23923_ (.A0(_19439_),
    .A1(_19440_),
    .S(_19428_),
    .X(_02727_));
 sky130_fd_sc_hd__buf_1 _23924_ (.A(_19408_),
    .X(_19441_));
 sky130_fd_sc_hd__and2_2 _23925_ (.A(\decoded_imm_uj[13] ),
    .B(_19437_),
    .X(_19442_));
 sky130_fd_sc_hd__a221o_2 _23926_ (.A1(_18912_),
    .A2(_19435_),
    .B1(_19441_),
    .B2(_19436_),
    .C1(_19442_),
    .X(_19443_));
 sky130_fd_sc_hd__buf_1 _23927_ (.A(\decoded_imm[13] ),
    .X(_19444_));
 sky130_fd_sc_hd__mux2_2 _23928_ (.A0(_19443_),
    .A1(_19444_),
    .S(_19428_),
    .X(_02726_));
 sky130_fd_sc_hd__buf_1 _23929_ (.A(\decoded_imm[14] ),
    .X(_19445_));
 sky130_vsdinv _23930_ (.A(_19445_),
    .Y(_19446_));
 sky130_fd_sc_hd__buf_1 _23931_ (.A(_18916_),
    .X(_19447_));
 sky130_fd_sc_hd__buf_1 _23932_ (.A(_17082_),
    .X(_19448_));
 sky130_fd_sc_hd__and2_2 _23933_ (.A(\decoded_imm_uj[14] ),
    .B(_19448_),
    .X(_19449_));
 sky130_fd_sc_hd__a221oi_2 _23934_ (.A1(_17272_),
    .A2(_19434_),
    .B1(_19409_),
    .B2(_19447_),
    .C1(_19449_),
    .Y(_19450_));
 sky130_fd_sc_hd__or2b_2 _23935_ (.A(_19450_),
    .B_N(_17331_),
    .X(_19451_));
 sky130_fd_sc_hd__o21ai_2 _23936_ (.A1(_19446_),
    .A2(_18903_),
    .B1(_19451_),
    .Y(_02725_));
 sky130_fd_sc_hd__and2_2 _23937_ (.A(\decoded_imm_uj[15] ),
    .B(_19437_),
    .X(_19452_));
 sky130_fd_sc_hd__a221o_2 _23938_ (.A1(\mem_rdata_q[15] ),
    .A2(_19435_),
    .B1(_19441_),
    .B2(_19436_),
    .C1(_19452_),
    .X(_19453_));
 sky130_fd_sc_hd__buf_1 _23939_ (.A(\decoded_imm[15] ),
    .X(_19454_));
 sky130_fd_sc_hd__mux2_2 _23940_ (.A0(_19453_),
    .A1(_19454_),
    .S(_19428_),
    .X(_02724_));
 sky130_fd_sc_hd__buf_1 _23941_ (.A(_19434_),
    .X(_19455_));
 sky130_fd_sc_hd__and2_2 _23942_ (.A(\decoded_imm_uj[16] ),
    .B(_19437_),
    .X(_19456_));
 sky130_fd_sc_hd__a221o_2 _23943_ (.A1(\mem_rdata_q[16] ),
    .A2(_19455_),
    .B1(_19441_),
    .B2(_19436_),
    .C1(_19456_),
    .X(_19457_));
 sky130_fd_sc_hd__buf_1 _23944_ (.A(\decoded_imm[16] ),
    .X(_19458_));
 sky130_fd_sc_hd__buf_1 _23945_ (.A(_18972_),
    .X(_19459_));
 sky130_fd_sc_hd__mux2_2 _23946_ (.A0(_19457_),
    .A1(_19458_),
    .S(_19459_),
    .X(_02723_));
 sky130_fd_sc_hd__and2_2 _23947_ (.A(\decoded_imm_uj[17] ),
    .B(_19448_),
    .X(_19460_));
 sky130_fd_sc_hd__a221o_2 _23948_ (.A1(\mem_rdata_q[17] ),
    .A2(_19455_),
    .B1(_19441_),
    .B2(_19447_),
    .C1(_19460_),
    .X(_19461_));
 sky130_fd_sc_hd__buf_1 _23949_ (.A(\decoded_imm[17] ),
    .X(_19462_));
 sky130_fd_sc_hd__mux2_2 _23950_ (.A0(_19461_),
    .A1(_19462_),
    .S(_19459_),
    .X(_02722_));
 sky130_fd_sc_hd__and2_2 _23951_ (.A(_18926_),
    .B(_19448_),
    .X(_19463_));
 sky130_fd_sc_hd__a221o_2 _23952_ (.A1(\mem_rdata_q[18] ),
    .A2(_19455_),
    .B1(_19409_),
    .B2(_19447_),
    .C1(_19463_),
    .X(_19464_));
 sky130_fd_sc_hd__buf_1 _23953_ (.A(\decoded_imm[18] ),
    .X(_19465_));
 sky130_fd_sc_hd__mux2_2 _23954_ (.A0(_19464_),
    .A1(_19465_),
    .S(_19459_),
    .X(_02721_));
 sky130_fd_sc_hd__and2_2 _23955_ (.A(\decoded_imm_uj[19] ),
    .B(_19448_),
    .X(_19466_));
 sky130_fd_sc_hd__a221o_2 _23956_ (.A1(\mem_rdata_q[19] ),
    .A2(_19455_),
    .B1(_19409_),
    .B2(_19447_),
    .C1(_19466_),
    .X(_19467_));
 sky130_fd_sc_hd__buf_1 _23957_ (.A(\decoded_imm[19] ),
    .X(_19468_));
 sky130_fd_sc_hd__mux2_2 _23958_ (.A0(_19467_),
    .A1(_19468_),
    .S(_19459_),
    .X(_02720_));
 sky130_fd_sc_hd__a2bb2oi_2 _23959_ (.A1_N(_17248_),
    .A2_N(_19391_),
    .B1(_18923_),
    .B2(_17083_),
    .Y(_19469_));
 sky130_fd_sc_hd__buf_1 _23960_ (.A(_19469_),
    .X(_19470_));
 sky130_fd_sc_hd__buf_1 _23961_ (.A(_19470_),
    .X(_19471_));
 sky130_fd_sc_hd__buf_1 _23962_ (.A(_16988_),
    .X(_19472_));
 sky130_fd_sc_hd__buf_1 _23963_ (.A(_19472_),
    .X(_19473_));
 sky130_fd_sc_hd__o21a_2 _23964_ (.A1(_18938_),
    .A2(_19473_),
    .B1(_18026_),
    .X(_19474_));
 sky130_fd_sc_hd__o31ai_2 _23965_ (.A1(is_alu_reg_imm),
    .A2(is_lb_lh_lw_lbu_lhu),
    .A3(_17086_),
    .B1(_18916_),
    .Y(_19475_));
 sky130_fd_sc_hd__buf_1 _23966_ (.A(_19475_),
    .X(_19476_));
 sky130_fd_sc_hd__buf_1 _23967_ (.A(_19476_),
    .X(_19477_));
 sky130_vsdinv _23968_ (.A(\decoded_imm[20] ),
    .Y(_19478_));
 sky130_fd_sc_hd__a32oi_2 _23969_ (.A1(_19471_),
    .A2(_19474_),
    .A3(_19477_),
    .B1(_19478_),
    .B2(_18989_),
    .Y(_02719_));
 sky130_fd_sc_hd__buf_1 _23970_ (.A(_19434_),
    .X(_19479_));
 sky130_fd_sc_hd__buf_1 _23971_ (.A(_17289_),
    .X(_19480_));
 sky130_fd_sc_hd__a21boi_2 _23972_ (.A1(_19479_),
    .A2(_19032_),
    .B1_N(_19480_),
    .Y(_19481_));
 sky130_fd_sc_hd__buf_1 _23973_ (.A(_19469_),
    .X(_19482_));
 sky130_fd_sc_hd__buf_1 _23974_ (.A(\decoded_imm[21] ),
    .X(_19483_));
 sky130_vsdinv _23975_ (.A(_19483_),
    .Y(_19484_));
 sky130_fd_sc_hd__buf_1 _23976_ (.A(_18954_),
    .X(_19485_));
 sky130_fd_sc_hd__a32oi_2 _23977_ (.A1(_19481_),
    .A2(_19482_),
    .A3(_19477_),
    .B1(_19484_),
    .B2(_19485_),
    .Y(_02718_));
 sky130_fd_sc_hd__a21boi_2 _23978_ (.A1(_19479_),
    .A2(_19029_),
    .B1_N(_17290_),
    .Y(_19486_));
 sky130_vsdinv _23979_ (.A(\decoded_imm[22] ),
    .Y(_19487_));
 sky130_fd_sc_hd__a32oi_2 _23980_ (.A1(_19486_),
    .A2(_19482_),
    .A3(_19477_),
    .B1(_19487_),
    .B2(_19485_),
    .Y(_02717_));
 sky130_fd_sc_hd__a21boi_2 _23981_ (.A1(_19479_),
    .A2(_19028_),
    .B1_N(_17290_),
    .Y(_19488_));
 sky130_fd_sc_hd__buf_1 _23982_ (.A(\decoded_imm[23] ),
    .X(_19489_));
 sky130_vsdinv _23983_ (.A(_19489_),
    .Y(_19490_));
 sky130_fd_sc_hd__a32oi_2 _23984_ (.A1(_19488_),
    .A2(_19482_),
    .A3(_19477_),
    .B1(_19490_),
    .B2(_19485_),
    .Y(_02716_));
 sky130_fd_sc_hd__buf_1 _23985_ (.A(\decoded_imm[24] ),
    .X(_19491_));
 sky130_fd_sc_hd__o21a_2 _23986_ (.A1(_18980_),
    .A2(_19472_),
    .B1(_19026_),
    .X(_19492_));
 sky130_fd_sc_hd__nand3_2 _23987_ (.A(_19482_),
    .B(_19492_),
    .C(_19476_),
    .Y(_19493_));
 sky130_fd_sc_hd__o21a_2 _23988_ (.A1(_19491_),
    .A2(_18027_),
    .B1(_19493_),
    .X(_02715_));
 sky130_fd_sc_hd__o21a_2 _23989_ (.A1(_18947_),
    .A2(_19473_),
    .B1(_19480_),
    .X(_19494_));
 sky130_fd_sc_hd__buf_1 _23990_ (.A(_19475_),
    .X(_19495_));
 sky130_fd_sc_hd__buf_1 _23991_ (.A(\decoded_imm[25] ),
    .X(_19496_));
 sky130_vsdinv _23992_ (.A(_19496_),
    .Y(_19497_));
 sky130_fd_sc_hd__a32oi_2 _23993_ (.A1(_19471_),
    .A2(_19494_),
    .A3(_19495_),
    .B1(_19497_),
    .B2(_19485_),
    .Y(_02714_));
 sky130_fd_sc_hd__o21a_2 _23994_ (.A1(_18993_),
    .A2(_19473_),
    .B1(_19480_),
    .X(_19498_));
 sky130_fd_sc_hd__buf_1 _23995_ (.A(\decoded_imm[26] ),
    .X(_19499_));
 sky130_vsdinv _23996_ (.A(_19499_),
    .Y(_19500_));
 sky130_fd_sc_hd__a32oi_2 _23997_ (.A1(_19471_),
    .A2(_19498_),
    .A3(_19495_),
    .B1(_19500_),
    .B2(_18965_),
    .Y(_02713_));
 sky130_fd_sc_hd__buf_1 _23998_ (.A(\decoded_imm[27] ),
    .X(_19501_));
 sky130_fd_sc_hd__o21a_2 _23999_ (.A1(_18977_),
    .A2(_19472_),
    .B1(_19026_),
    .X(_19502_));
 sky130_fd_sc_hd__nand3_2 _24000_ (.A(_19470_),
    .B(_19502_),
    .C(_19476_),
    .Y(_19503_));
 sky130_fd_sc_hd__o21a_2 _24001_ (.A1(_19501_),
    .A2(_19025_),
    .B1(_19503_),
    .X(_02712_));
 sky130_fd_sc_hd__buf_1 _24002_ (.A(\decoded_imm[28] ),
    .X(_19504_));
 sky130_fd_sc_hd__a21boi_2 _24003_ (.A1(_19479_),
    .A2(_18959_),
    .B1_N(_17290_),
    .Y(_19505_));
 sky130_fd_sc_hd__nand3_2 _24004_ (.A(_19505_),
    .B(_19495_),
    .C(_19470_),
    .Y(_19506_));
 sky130_fd_sc_hd__o21a_2 _24005_ (.A1(_19504_),
    .A2(_19025_),
    .B1(_19506_),
    .X(_02711_));
 sky130_fd_sc_hd__o21a_2 _24006_ (.A1(_17250_),
    .A2(_19473_),
    .B1(_19480_),
    .X(_19507_));
 sky130_fd_sc_hd__buf_1 _24007_ (.A(\decoded_imm[29] ),
    .X(_19508_));
 sky130_vsdinv _24008_ (.A(_19508_),
    .Y(_19509_));
 sky130_fd_sc_hd__a32oi_2 _24009_ (.A1(_19471_),
    .A2(_19507_),
    .A3(_19495_),
    .B1(_19509_),
    .B2(_18965_),
    .Y(_02710_));
 sky130_fd_sc_hd__buf_1 _24010_ (.A(\decoded_imm[30] ),
    .X(_19510_));
 sky130_fd_sc_hd__o21a_2 _24011_ (.A1(_17249_),
    .A2(_19472_),
    .B1(_19026_),
    .X(_19511_));
 sky130_fd_sc_hd__nand3_2 _24012_ (.A(_19470_),
    .B(_19511_),
    .C(_19476_),
    .Y(_19512_));
 sky130_fd_sc_hd__o21a_2 _24013_ (.A1(_19510_),
    .A2(_19025_),
    .B1(_19512_),
    .X(_02709_));
 sky130_fd_sc_hd__nor2_2 _24014_ (.A(_19435_),
    .B(_19420_),
    .Y(_19513_));
 sky130_fd_sc_hd__buf_1 _24015_ (.A(_18922_),
    .X(_19514_));
 sky130_fd_sc_hd__and2_2 _24016_ (.A(_19514_),
    .B(_17083_),
    .X(_19515_));
 sky130_fd_sc_hd__o21bai_2 _24017_ (.A1(_17248_),
    .A2(_19513_),
    .B1_N(_19515_),
    .Y(_19516_));
 sky130_fd_sc_hd__mux2_2 _24018_ (.A0(_19516_),
    .A1(\decoded_imm[31] ),
    .S(_18954_),
    .X(_02708_));
 sky130_fd_sc_hd__buf_1 _24019_ (.A(_17057_),
    .X(_19517_));
 sky130_fd_sc_hd__nor3b_2 _24020_ (.A(_19517_),
    .B(_17859_),
    .C_N(_19778_),
    .Y(_19518_));
 sky130_fd_sc_hd__and2_2 _24021_ (.A(_18544_),
    .B(_17020_),
    .X(_19519_));
 sky130_fd_sc_hd__mux2_2 _24022_ (.A0(_18283_),
    .A1(_19518_),
    .S(_19519_),
    .X(_02707_));
 sky130_fd_sc_hd__nand2_2 _24023_ (.A(_16983_),
    .B(_17020_),
    .Y(_02542_));
 sky130_fd_sc_hd__buf_1 _24024_ (.A(_19519_),
    .X(_19520_));
 sky130_vsdinv _24025_ (.A(_19520_),
    .Y(_19521_));
 sky130_fd_sc_hd__and3b_2 _24026_ (.A_N(_02542_),
    .B(_17051_),
    .C(_18022_),
    .X(_19522_));
 sky130_fd_sc_hd__nand3_2 _24027_ (.A(_19522_),
    .B(\decoded_rd[1] ),
    .C(_19519_),
    .Y(_19523_));
 sky130_fd_sc_hd__a21bo_2 _24028_ (.A1(_18284_),
    .A2(_19521_),
    .B1_N(_19523_),
    .X(_02706_));
 sky130_fd_sc_hd__nand3_2 _24029_ (.A(_19522_),
    .B(\decoded_rd[2] ),
    .C(_19520_),
    .Y(_19524_));
 sky130_fd_sc_hd__o21ai_2 _24030_ (.A1(_18277_),
    .A2(_19520_),
    .B1(_19524_),
    .Y(_02705_));
 sky130_fd_sc_hd__nand3_2 _24031_ (.A(_19522_),
    .B(\decoded_rd[3] ),
    .C(_19519_),
    .Y(_19525_));
 sky130_fd_sc_hd__o21ai_2 _24032_ (.A1(_18278_),
    .A2(_19520_),
    .B1(_19525_),
    .Y(_02704_));
 sky130_fd_sc_hd__nand2_2 _24033_ (.A(_17062_),
    .B(_17065_),
    .Y(_19526_));
 sky130_fd_sc_hd__a21oi_2 _24034_ (.A1(_17004_),
    .A2(_17015_),
    .B1(_19526_),
    .Y(_19527_));
 sky130_vsdinv _24035_ (.A(_19527_),
    .Y(_19528_));
 sky130_fd_sc_hd__o31ai_2 _24036_ (.A1(is_jalr_addi_slti_sltiu_xori_ori_andi),
    .A2(is_slli_srli_srai),
    .A3(is_lui_auipc_jal),
    .B1(_16829_),
    .Y(_19529_));
 sky130_fd_sc_hd__a21oi_2 _24037_ (.A1(_19528_),
    .A2(_19529_),
    .B1(_18384_),
    .Y(_02703_));
 sky130_fd_sc_hd__buf_1 _24038_ (.A(_18852_),
    .X(_19530_));
 sky130_fd_sc_hd__nor2b_2 _24039_ (.A(_19530_),
    .B_N(_02558_),
    .Y(_02702_));
 sky130_fd_sc_hd__nor2b_2 _24040_ (.A(_19530_),
    .B_N(_02557_),
    .Y(_02701_));
 sky130_fd_sc_hd__nor2b_2 _24041_ (.A(_19530_),
    .B_N(_02556_),
    .Y(_02700_));
 sky130_fd_sc_hd__nor2b_2 _24042_ (.A(_19530_),
    .B_N(_02555_),
    .Y(_02699_));
 sky130_fd_sc_hd__buf_1 _24043_ (.A(_18852_),
    .X(_19531_));
 sky130_fd_sc_hd__nor2b_2 _24044_ (.A(_19531_),
    .B_N(_02554_),
    .Y(_02698_));
 sky130_fd_sc_hd__nor2b_2 _24045_ (.A(_19531_),
    .B_N(_02553_),
    .Y(_02697_));
 sky130_fd_sc_hd__nor2b_2 _24046_ (.A(_19531_),
    .B_N(_02552_),
    .Y(_02696_));
 sky130_fd_sc_hd__nor2b_2 _24047_ (.A(_19531_),
    .B_N(_02551_),
    .Y(_02695_));
 sky130_fd_sc_hd__buf_1 _24048_ (.A(_18445_),
    .X(_19532_));
 sky130_fd_sc_hd__nor2b_2 _24049_ (.A(_19532_),
    .B_N(_00122_),
    .Y(_02550_));
 sky130_fd_sc_hd__buf_1 _24050_ (.A(_18852_),
    .X(_19533_));
 sky130_fd_sc_hd__buf_1 _24051_ (.A(_18445_),
    .X(_19534_));
 sky130_fd_sc_hd__nor3b_2 _24052_ (.A(_19533_),
    .B(_19534_),
    .C_N(_00122_),
    .Y(_02694_));
 sky130_fd_sc_hd__nor2b_2 _24053_ (.A(_19532_),
    .B_N(_00116_),
    .Y(_02549_));
 sky130_fd_sc_hd__buf_1 _24054_ (.A(_18445_),
    .X(_19535_));
 sky130_fd_sc_hd__nor3b_2 _24055_ (.A(_19533_),
    .B(_19535_),
    .C_N(_00116_),
    .Y(_02693_));
 sky130_fd_sc_hd__nor2b_2 _24056_ (.A(_19532_),
    .B_N(_00110_),
    .Y(_02548_));
 sky130_fd_sc_hd__nor3b_2 _24057_ (.A(_19533_),
    .B(_19535_),
    .C_N(_00110_),
    .Y(_02692_));
 sky130_fd_sc_hd__nor2b_2 _24058_ (.A(_19532_),
    .B_N(_00104_),
    .Y(_02547_));
 sky130_fd_sc_hd__nor3b_2 _24059_ (.A(_18442_),
    .B(_19535_),
    .C_N(_00104_),
    .Y(_02691_));
 sky130_fd_sc_hd__nor3b_2 _24060_ (.A(_19534_),
    .B(_18526_),
    .C_N(_00094_),
    .Y(_02546_));
 sky130_vsdinv _24061_ (.A(mem_la_wdata[4]),
    .Y(_19536_));
 sky130_fd_sc_hd__buf_1 _24062_ (.A(_19536_),
    .X(_19537_));
 sky130_fd_sc_hd__buf_1 _24063_ (.A(_19537_),
    .X(_02327_));
 sky130_vsdinv _24064_ (.A(mem_la_wdata[3]),
    .Y(_19538_));
 sky130_fd_sc_hd__buf_1 _24065_ (.A(_19538_),
    .X(_02324_));
 sky130_vsdinv _24066_ (.A(_18447_),
    .Y(_19539_));
 sky130_fd_sc_hd__buf_1 _24067_ (.A(_19539_),
    .X(_19540_));
 sky130_fd_sc_hd__and4_2 _24068_ (.A(_02327_),
    .B(_02324_),
    .C(_19540_),
    .D(_00094_),
    .X(_02690_));
 sky130_fd_sc_hd__nor3b_2 _24069_ (.A(_19534_),
    .B(_18526_),
    .C_N(_00084_),
    .Y(_02545_));
 sky130_fd_sc_hd__and4_2 _24070_ (.A(_02327_),
    .B(_02324_),
    .C(_19540_),
    .D(_00084_),
    .X(_02689_));
 sky130_fd_sc_hd__buf_1 _24071_ (.A(_19539_),
    .X(_02321_));
 sky130_vsdinv _24072_ (.A(_18449_),
    .Y(_19541_));
 sky130_fd_sc_hd__buf_1 _24073_ (.A(_19541_),
    .X(_02318_));
 sky130_fd_sc_hd__and4_2 _24074_ (.A(_02324_),
    .B(_02321_),
    .C(_02318_),
    .D(_00066_),
    .X(_02544_));
 sky130_fd_sc_hd__nor2b_2 _24075_ (.A(_18451_),
    .B_N(_00066_),
    .Y(_00067_));
 sky130_fd_sc_hd__buf_1 _24076_ (.A(_19538_),
    .X(_19542_));
 sky130_fd_sc_hd__and4_2 _24077_ (.A(_00067_),
    .B(_02327_),
    .C(_19542_),
    .D(_02321_),
    .X(_02688_));
 sky130_fd_sc_hd__nor2b_2 _24078_ (.A(_18452_),
    .B_N(_19119_),
    .Y(_00048_));
 sky130_fd_sc_hd__and4_2 _24079_ (.A(_00048_),
    .B(_19542_),
    .C(_19540_),
    .D(_02318_),
    .X(_02543_));
 sky130_fd_sc_hd__buf_1 _24080_ (.A(_19122_),
    .X(_19543_));
 sky130_fd_sc_hd__nor3b_2 _24081_ (.A(_18450_),
    .B(_18454_),
    .C_N(_19543_),
    .Y(_00049_));
 sky130_fd_sc_hd__and4_2 _24082_ (.A(_00049_),
    .B(_19537_),
    .C(_19542_),
    .D(_19540_),
    .X(_02687_));
 sky130_fd_sc_hd__buf_1 _24083_ (.A(_17073_),
    .X(_00297_));
 sky130_fd_sc_hd__o211a_2 _24084_ (.A1(_17594_),
    .A2(\reg_next_pc[0] ),
    .B1(resetn),
    .C1(mem_do_rinst),
    .X(_19544_));
 sky130_fd_sc_hd__buf_1 _24085_ (.A(_19544_),
    .X(_19545_));
 sky130_fd_sc_hd__buf_1 _24086_ (.A(_19545_),
    .X(_19546_));
 sky130_fd_sc_hd__buf_1 _24087_ (.A(_19546_),
    .X(_19547_));
 sky130_fd_sc_hd__buf_1 _24088_ (.A(_19547_),
    .X(_00307_));
 sky130_fd_sc_hd__buf_1 _24089_ (.A(_16936_),
    .X(_19548_));
 sky130_fd_sc_hd__buf_1 _24090_ (.A(_17990_),
    .X(_19549_));
 sky130_fd_sc_hd__nor3_2 _24091_ (.A(_19548_),
    .B(_17194_),
    .C(_19549_),
    .Y(_00312_));
 sky130_fd_sc_hd__o21a_2 _24092_ (.A1(mem_do_wdata),
    .A2(mem_do_rdata),
    .B1(resetn),
    .X(_19550_));
 sky130_fd_sc_hd__buf_1 _24093_ (.A(_19550_),
    .X(_19551_));
 sky130_fd_sc_hd__buf_1 _24094_ (.A(_19551_),
    .X(_00303_));
 sky130_fd_sc_hd__and2_2 _24095_ (.A(_19120_),
    .B(\mem_wordsize[2] ),
    .X(_19552_));
 sky130_fd_sc_hd__o21a_2 _24096_ (.A1(_19115_),
    .A2(_19119_),
    .B1(\mem_wordsize[0] ),
    .X(_19553_));
 sky130_fd_sc_hd__o21a_2 _24097_ (.A1(_19552_),
    .A2(_19553_),
    .B1(_19550_),
    .X(_19554_));
 sky130_fd_sc_hd__buf_1 _24098_ (.A(_19554_),
    .X(_19555_));
 sky130_fd_sc_hd__buf_1 _24099_ (.A(_16880_),
    .X(_19556_));
 sky130_fd_sc_hd__o21a_2 _24100_ (.A1(_16924_),
    .A2(_18021_),
    .B1(_16881_),
    .X(_19557_));
 sky130_fd_sc_hd__o2111a_2 _24101_ (.A1(_16879_),
    .A2(_19556_),
    .B1(instr_jal),
    .C1(_16927_),
    .D1(_19557_),
    .X(_02062_));
 sky130_fd_sc_hd__nand3b_2 _24102_ (.A_N(_19555_),
    .B(_02062_),
    .C(_18382_),
    .Y(_19558_));
 sky130_fd_sc_hd__nor2_2 _24103_ (.A(irq_active),
    .B(_17989_),
    .Y(_19559_));
 sky130_vsdinv _24104_ (.A(_19559_),
    .Y(_19560_));
 sky130_fd_sc_hd__buf_1 _24105_ (.A(_19552_),
    .X(_19561_));
 sky130_fd_sc_hd__buf_1 _24106_ (.A(_19553_),
    .X(_19562_));
 sky130_fd_sc_hd__nor2_2 _24107_ (.A(_16848_),
    .B(_16811_),
    .Y(_19563_));
 sky130_fd_sc_hd__o21bai_2 _24108_ (.A1(_19561_),
    .A2(_19562_),
    .B1_N(_19563_),
    .Y(_19564_));
 sky130_fd_sc_hd__buf_1 _24109_ (.A(_19557_),
    .X(_19565_));
 sky130_fd_sc_hd__buf_1 _24110_ (.A(_19550_),
    .X(_19566_));
 sky130_vsdinv _24111_ (.A(_19120_),
    .Y(_19567_));
 sky130_vsdinv _24112_ (.A(\mem_wordsize[2] ),
    .Y(_19568_));
 sky130_fd_sc_hd__o2111a_2 _24113_ (.A1(_19567_),
    .A2(_19568_),
    .B1(_19559_),
    .C1(_19550_),
    .D1(_19553_),
    .X(_19569_));
 sky130_vsdinv _24114_ (.A(_19569_),
    .Y(_19570_));
 sky130_fd_sc_hd__o2111ai_2 _24115_ (.A1(_18956_),
    .A2(_19556_),
    .B1(_16814_),
    .C1(_17266_),
    .D1(_19565_),
    .Y(_19571_));
 sky130_fd_sc_hd__a21o_2 _24116_ (.A1(_19566_),
    .A2(_19570_),
    .B1(_19571_),
    .X(_19572_));
 sky130_fd_sc_hd__o41a_2 _24117_ (.A1(_16930_),
    .A2(_19560_),
    .A3(_19564_),
    .A4(_19565_),
    .B1(_19572_),
    .X(_19573_));
 sky130_fd_sc_hd__buf_1 _24118_ (.A(_19561_),
    .X(_19574_));
 sky130_fd_sc_hd__buf_1 _24119_ (.A(_19562_),
    .X(_19575_));
 sky130_fd_sc_hd__buf_1 _24120_ (.A(_19559_),
    .X(_19576_));
 sky130_fd_sc_hd__o211a_2 _24121_ (.A1(_19116_),
    .A2(_19120_),
    .B1(\mem_wordsize[0] ),
    .C1(_19576_),
    .X(_19577_));
 sky130_fd_sc_hd__nand3_2 _24122_ (.A(_02062_),
    .B(_17221_),
    .C(_19577_),
    .Y(_19578_));
 sky130_fd_sc_hd__o21ai_2 _24123_ (.A1(_19575_),
    .A2(_19571_),
    .B1(_19578_),
    .Y(_19579_));
 sky130_fd_sc_hd__nand3b_2 _24124_ (.A_N(_19574_),
    .B(_19579_),
    .C(_00303_),
    .Y(_19580_));
 sky130_fd_sc_hd__o2111a_2 _24125_ (.A1(_18024_),
    .A2(_00303_),
    .B1(_19558_),
    .C1(_19573_),
    .D1(_19580_),
    .X(_19581_));
 sky130_fd_sc_hd__o2111a_2 _24126_ (.A1(_17594_),
    .A2(\reg_next_pc[0] ),
    .B1(_16806_),
    .C1(_16799_),
    .D1(_19559_),
    .X(_19582_));
 sky130_fd_sc_hd__buf_1 _24127_ (.A(_19582_),
    .X(_19583_));
 sky130_fd_sc_hd__buf_1 _24128_ (.A(_19576_),
    .X(_19584_));
 sky130_fd_sc_hd__buf_1 _24129_ (.A(_19561_),
    .X(_00306_));
 sky130_fd_sc_hd__o2111a_2 _24130_ (.A1(_17217_),
    .A2(_17388_),
    .B1(_18382_),
    .C1(_19584_),
    .D1(_00306_),
    .X(_19585_));
 sky130_fd_sc_hd__o211ai_2 _24131_ (.A1(_19583_),
    .A2(_19585_),
    .B1(_17119_),
    .C1(_02062_),
    .Y(_19586_));
 sky130_fd_sc_hd__buf_1 _24132_ (.A(_19560_),
    .X(_19587_));
 sky130_fd_sc_hd__buf_1 _24133_ (.A(_19544_),
    .X(_19588_));
 sky130_vsdinv _24134_ (.A(_19566_),
    .Y(_19589_));
 sky130_fd_sc_hd__a2111o_2 _24135_ (.A1(_19587_),
    .A2(_19575_),
    .B1(_19574_),
    .C1(_19588_),
    .D1(_19589_),
    .X(_19590_));
 sky130_fd_sc_hd__and3_2 _24136_ (.A(_16925_),
    .B(_17221_),
    .C(_16881_),
    .X(_19591_));
 sky130_fd_sc_hd__buf_1 _24137_ (.A(_18023_),
    .X(_00309_));
 sky130_fd_sc_hd__nand3b_2 _24138_ (.A_N(_19590_),
    .B(_19591_),
    .C(_00309_),
    .Y(_19592_));
 sky130_fd_sc_hd__o2111ai_2 _24139_ (.A1(_18956_),
    .A2(_19556_),
    .B1(_17301_),
    .C1(_19583_),
    .D1(_19591_),
    .Y(_19593_));
 sky130_fd_sc_hd__o2111a_2 _24140_ (.A1(_00307_),
    .A2(_19581_),
    .B1(_19586_),
    .C1(_19592_),
    .D1(_19593_),
    .X(_19594_));
 sky130_fd_sc_hd__o2111ai_2 _24141_ (.A1(_18956_),
    .A2(_19556_),
    .B1(_17393_),
    .C1(_17266_),
    .D1(_19591_),
    .Y(_19595_));
 sky130_fd_sc_hd__nor2_2 _24142_ (.A(_16935_),
    .B(_17209_),
    .Y(_19596_));
 sky130_fd_sc_hd__o211a_2 _24143_ (.A1(instr_ecall_ebreak),
    .A2(pcpi_timeout),
    .B1(_16954_),
    .C1(_19596_),
    .X(_19597_));
 sky130_fd_sc_hd__nand3b_2 _24144_ (.A_N(_18000_),
    .B(_16837_),
    .C(_19597_),
    .Y(_19598_));
 sky130_fd_sc_hd__nand3b_2 _24145_ (.A_N(_19545_),
    .B(_19576_),
    .C(_19561_),
    .Y(_19599_));
 sky130_fd_sc_hd__a21oi_2 _24146_ (.A1(_19595_),
    .A2(_19598_),
    .B1(_19599_),
    .Y(_19600_));
 sky130_fd_sc_hd__nor3_2 _24147_ (.A(_16808_),
    .B(_16805_),
    .C(_16804_),
    .Y(_19601_));
 sky130_vsdinv _24148_ (.A(_19601_),
    .Y(_19602_));
 sky130_fd_sc_hd__buf_1 _24149_ (.A(_19562_),
    .X(_00305_));
 sky130_fd_sc_hd__o21a_2 _24150_ (.A1(_00306_),
    .A2(_00305_),
    .B1(_19587_),
    .X(_19603_));
 sky130_fd_sc_hd__nand3_2 _24151_ (.A(_19591_),
    .B(_17027_),
    .C(_18023_),
    .Y(_19604_));
 sky130_fd_sc_hd__or2_2 _24152_ (.A(_19599_),
    .B(_19604_),
    .X(_19605_));
 sky130_fd_sc_hd__o41ai_2 _24153_ (.A1(_00297_),
    .A2(_19602_),
    .A3(_19547_),
    .A4(_19603_),
    .B1(_19605_),
    .Y(_19606_));
 sky130_fd_sc_hd__buf_1 _24154_ (.A(_19589_),
    .X(_19607_));
 sky130_fd_sc_hd__o21bai_2 _24155_ (.A1(_19600_),
    .A2(_19606_),
    .B1_N(_19607_),
    .Y(_19608_));
 sky130_vsdinv _24156_ (.A(_19582_),
    .Y(_19609_));
 sky130_fd_sc_hd__o21a_2 _24157_ (.A1(_19545_),
    .A2(_19554_),
    .B1(_19609_),
    .X(_19610_));
 sky130_fd_sc_hd__buf_1 _24158_ (.A(_19610_),
    .X(_19611_));
 sky130_fd_sc_hd__buf_1 _24159_ (.A(_19546_),
    .X(_19612_));
 sky130_fd_sc_hd__nand3_2 _24160_ (.A(_19612_),
    .B(_00309_),
    .C(_19584_),
    .Y(_19613_));
 sky130_fd_sc_hd__o31a_2 _24161_ (.A1(_17147_),
    .A2(_19611_),
    .A3(_19565_),
    .B1(_19613_),
    .X(_19614_));
 sky130_fd_sc_hd__a2111o_2 _24162_ (.A1(_19560_),
    .A2(_19575_),
    .B1(_19574_),
    .C1(_19588_),
    .D1(_19589_),
    .X(_19615_));
 sky130_fd_sc_hd__o21bai_2 _24163_ (.A1(_19552_),
    .A2(_19544_),
    .B1_N(_19560_),
    .Y(_19616_));
 sky130_fd_sc_hd__o21a_2 _24164_ (.A1(_19588_),
    .A2(_19551_),
    .B1(_19616_),
    .X(_19617_));
 sky130_fd_sc_hd__a21oi_2 _24165_ (.A1(_19615_),
    .A2(_19617_),
    .B1(_16954_),
    .Y(_19618_));
 sky130_fd_sc_hd__and2_2 _24166_ (.A(_19566_),
    .B(_19562_),
    .X(_19619_));
 sky130_vsdinv _24167_ (.A(_19544_),
    .Y(_19620_));
 sky130_fd_sc_hd__buf_1 _24168_ (.A(_19620_),
    .X(_19621_));
 sky130_fd_sc_hd__a211oi_2 _24169_ (.A1(_19121_),
    .A2(\mem_wordsize[2] ),
    .B1(_16935_),
    .C1(_17989_),
    .Y(_19622_));
 sky130_fd_sc_hd__nand3_2 _24170_ (.A(_19619_),
    .B(_19621_),
    .C(_19622_),
    .Y(_19623_));
 sky130_fd_sc_hd__a21boi_2 _24171_ (.A1(_19610_),
    .A2(_19623_),
    .B1_N(_19597_),
    .Y(_19624_));
 sky130_fd_sc_hd__buf_1 _24172_ (.A(_17017_),
    .X(_19625_));
 sky130_fd_sc_hd__buf_1 _24173_ (.A(_17064_),
    .X(_00310_));
 sky130_fd_sc_hd__o2111ai_2 _24174_ (.A1(_19618_),
    .A2(_19624_),
    .B1(_17119_),
    .C1(_19625_),
    .D1(_00310_),
    .Y(_19626_));
 sky130_fd_sc_hd__nor2_2 _24175_ (.A(_19551_),
    .B(_19588_),
    .Y(_19627_));
 sky130_fd_sc_hd__nor2_2 _24176_ (.A(_19627_),
    .B(_19616_),
    .Y(_19628_));
 sky130_fd_sc_hd__nand2_2 _24177_ (.A(_19564_),
    .B(_18382_),
    .Y(_19629_));
 sky130_fd_sc_hd__a21oi_2 _24178_ (.A1(_19570_),
    .A2(_19629_),
    .B1(_19612_),
    .Y(_19630_));
 sky130_fd_sc_hd__nand3b_2 _24179_ (.A_N(instr_rdcycle),
    .B(_01717_),
    .C(_01714_),
    .Y(_19631_));
 sky130_fd_sc_hd__o211ai_2 _24180_ (.A1(_19628_),
    .A2(_19630_),
    .B1(_17966_),
    .C1(_19631_),
    .Y(_19632_));
 sky130_vsdinv _24181_ (.A(_17073_),
    .Y(_19633_));
 sky130_fd_sc_hd__o211a_2 _24182_ (.A1(_19583_),
    .A2(_19627_),
    .B1(_19633_),
    .C1(_19601_),
    .X(_19634_));
 sky130_fd_sc_hd__o2111ai_2 _24183_ (.A1(_19575_),
    .A2(_19574_),
    .B1(_19576_),
    .C1(_19551_),
    .D1(_19621_),
    .Y(_19635_));
 sky130_fd_sc_hd__or4b_2 _24184_ (.A(_16930_),
    .B(_16983_),
    .C(_16804_),
    .D_N(_17071_),
    .X(_19636_));
 sky130_fd_sc_hd__a21oi_2 _24185_ (.A1(_19611_),
    .A2(_19635_),
    .B1(_19636_),
    .Y(_19637_));
 sky130_fd_sc_hd__o2111ai_2 _24186_ (.A1(_19567_),
    .A2(_19568_),
    .B1(_19566_),
    .C1(_19577_),
    .D1(_19620_),
    .Y(_19638_));
 sky130_fd_sc_hd__nor3_2 _24187_ (.A(_16809_),
    .B(_18543_),
    .C(_19638_),
    .Y(_19639_));
 sky130_fd_sc_hd__o21a_2 _24188_ (.A1(_19545_),
    .A2(_19554_),
    .B1(_19616_),
    .X(_19640_));
 sky130_fd_sc_hd__nor3_2 _24189_ (.A(_16809_),
    .B(_18543_),
    .C(_19640_),
    .Y(_19641_));
 sky130_fd_sc_hd__or4_2 _24190_ (.A(_16841_),
    .B(_00314_),
    .C(_19639_),
    .D(_19641_),
    .X(_19642_));
 sky130_fd_sc_hd__nor3_2 _24191_ (.A(_19634_),
    .B(_19637_),
    .C(_19642_),
    .Y(_19643_));
 sky130_fd_sc_hd__o2111a_2 _24192_ (.A1(_17403_),
    .A2(_19614_),
    .B1(_19626_),
    .C1(_19632_),
    .D1(_19643_),
    .X(_19644_));
 sky130_fd_sc_hd__o211ai_2 _24193_ (.A1(_00322_),
    .A2(_19594_),
    .B1(_19608_),
    .C1(_19644_),
    .Y(_00039_));
 sky130_fd_sc_hd__a21oi_2 _24194_ (.A1(_19564_),
    .A2(_19621_),
    .B1(_19584_),
    .Y(_19645_));
 sky130_fd_sc_hd__nor3b_2 _24195_ (.A(_17782_),
    .B(_19645_),
    .C_N(_17085_),
    .Y(_00040_));
 sky130_vsdinv _24196_ (.A(_17387_),
    .Y(_19646_));
 sky130_fd_sc_hd__o21a_2 _24197_ (.A1(_19546_),
    .A2(_19555_),
    .B1(_19587_),
    .X(_19647_));
 sky130_fd_sc_hd__nand3b_2 _24198_ (.A_N(_19647_),
    .B(_17060_),
    .C(_17859_),
    .Y(_19648_));
 sky130_fd_sc_hd__o41a_2 _24199_ (.A1(_16823_),
    .A2(_19646_),
    .A3(_00307_),
    .A4(_19555_),
    .B1(_19648_),
    .X(_19649_));
 sky130_fd_sc_hd__nor3_2 _24200_ (.A(_19563_),
    .B(_19612_),
    .C(_19603_),
    .Y(_19650_));
 sky130_fd_sc_hd__o311ai_2 _24201_ (.A1(_19583_),
    .A2(_19627_),
    .A3(_19650_),
    .B1(_16810_),
    .C1(_19602_),
    .Y(_19651_));
 sky130_fd_sc_hd__o2111ai_2 _24202_ (.A1(_19547_),
    .A2(_19555_),
    .B1(_17080_),
    .C1(_19584_),
    .D1(_17069_),
    .Y(_19652_));
 sky130_fd_sc_hd__a21oi_2 _24203_ (.A1(_19651_),
    .A2(_19652_),
    .B1(_16824_),
    .Y(_19653_));
 sky130_fd_sc_hd__o21bai_2 _24204_ (.A1(_17782_),
    .A2(_19649_),
    .B1_N(_19653_),
    .Y(_00044_));
 sky130_fd_sc_hd__a211o_2 _24205_ (.A1(_19640_),
    .A2(_19638_),
    .B1(\pcpi_mul.active[1] ),
    .C1(_18002_),
    .X(_19654_));
 sky130_fd_sc_hd__nand3b_2 _24206_ (.A_N(_17009_),
    .B(_16828_),
    .C(_01717_),
    .Y(_19655_));
 sky130_fd_sc_hd__nor2_2 _24207_ (.A(is_jalr_addi_slti_sltiu_xori_ori_andi),
    .B(is_slli_srli_srai),
    .Y(_01304_));
 sky130_fd_sc_hd__or4b_2 _24208_ (.A(_16931_),
    .B(is_lui_auipc_jal),
    .C(_19655_),
    .D_N(_01304_),
    .X(_19656_));
 sky130_fd_sc_hd__a21oi_2 _24209_ (.A1(_19590_),
    .A2(_19617_),
    .B1(_19656_),
    .Y(_19657_));
 sky130_fd_sc_hd__o21ai_2 _24210_ (.A1(_17059_),
    .A2(_00310_),
    .B1(_19657_),
    .Y(_19658_));
 sky130_fd_sc_hd__o31ai_2 _24211_ (.A1(_18001_),
    .A2(_19654_),
    .A3(_18000_),
    .B1(_19658_),
    .Y(_00041_));
 sky130_fd_sc_hd__o221ai_2 _24212_ (.A1(_16935_),
    .A2(_17209_),
    .B1(instr_ecall_ebreak),
    .B2(pcpi_timeout),
    .C1(_16954_),
    .Y(_19659_));
 sky130_fd_sc_hd__a211oi_2 _24213_ (.A1(_19611_),
    .A2(_19635_),
    .B1(_19659_),
    .C1(_18000_),
    .Y(_19660_));
 sky130_fd_sc_hd__o31a_2 _24214_ (.A1(\cpu_state[0] ),
    .A2(_19645_),
    .A3(_19660_),
    .B1(_17326_),
    .X(_00038_));
 sky130_fd_sc_hd__buf_1 _24215_ (.A(_17065_),
    .X(_19661_));
 sky130_fd_sc_hd__nand3_2 _24216_ (.A(_17803_),
    .B(_18936_),
    .C(_19661_),
    .Y(_19662_));
 sky130_fd_sc_hd__and3_2 _24217_ (.A(_17386_),
    .B(_16816_),
    .C(_17079_),
    .X(_19663_));
 sky130_fd_sc_hd__buf_1 _24218_ (.A(\cpu_state[5] ),
    .X(_19664_));
 sky130_fd_sc_hd__nand3_2 _24219_ (.A(_19663_),
    .B(_19664_),
    .C(_19619_),
    .Y(_19665_));
 sky130_fd_sc_hd__o31ai_2 _24220_ (.A1(_19587_),
    .A2(_19607_),
    .A3(_19662_),
    .B1(_19665_),
    .Y(_19666_));
 sky130_fd_sc_hd__buf_1 _24221_ (.A(\mem_wordsize[2] ),
    .X(_19667_));
 sky130_fd_sc_hd__a2111o_2 _24222_ (.A1(_19121_),
    .A2(_19667_),
    .B1(_00305_),
    .C1(_19546_),
    .D1(_19589_),
    .X(_19668_));
 sky130_fd_sc_hd__a21oi_2 _24223_ (.A1(_19668_),
    .A2(_19617_),
    .B1(_19662_),
    .Y(_19669_));
 sky130_fd_sc_hd__nand3b_2 _24224_ (.A_N(_19601_),
    .B(_16810_),
    .C(_19577_),
    .Y(_19670_));
 sky130_fd_sc_hd__nand3b_2 _24225_ (.A_N(_00305_),
    .B(_17068_),
    .C(_17079_),
    .Y(_19671_));
 sky130_fd_sc_hd__a2111o_2 _24226_ (.A1(_19670_),
    .A2(_19671_),
    .B1(_19547_),
    .C1(_19607_),
    .D1(_00306_),
    .X(_19672_));
 sky130_fd_sc_hd__or2b_2 _24227_ (.A(_19599_),
    .B_N(_00303_),
    .X(_19673_));
 sky130_fd_sc_hd__a2111o_2 _24228_ (.A1(_19673_),
    .A2(_19611_),
    .B1(_16842_),
    .C1(_19601_),
    .D1(_17387_),
    .X(_19674_));
 sky130_fd_sc_hd__nand3b_2 _24229_ (.A_N(_19617_),
    .B(_17068_),
    .C(_17079_),
    .Y(_19675_));
 sky130_fd_sc_hd__a31oi_2 _24230_ (.A1(_19672_),
    .A2(_19674_),
    .A3(_19675_),
    .B1(_18030_),
    .Y(_19676_));
 sky130_fd_sc_hd__a311o_2 _24231_ (.A1(_19621_),
    .A2(_19622_),
    .A3(_19666_),
    .B1(_19669_),
    .C1(_19676_),
    .X(_00043_));
 sky130_fd_sc_hd__o31a_2 _24232_ (.A1(_16845_),
    .A2(_17081_),
    .A3(_17388_),
    .B1(_17222_),
    .X(mem_la_read));
 sky130_fd_sc_hd__and3_2 _24233_ (.A(_00290_),
    .B(_16837_),
    .C(_17218_),
    .X(_19677_));
 sky130_fd_sc_hd__buf_1 _24234_ (.A(_19677_),
    .X(mem_la_write));
 sky130_fd_sc_hd__nand2_2 _24235_ (.A(_16850_),
    .B(_17222_),
    .Y(_00316_));
 sky130_fd_sc_hd__and2_2 _24236_ (.A(_16848_),
    .B(\cpu_state[5] ),
    .X(_00317_));
 sky130_fd_sc_hd__buf_1 _24237_ (.A(_17057_),
    .X(_19678_));
 sky130_fd_sc_hd__buf_1 _24238_ (.A(_19678_),
    .X(_19679_));
 sky130_vsdinv _24239_ (.A(_19628_),
    .Y(_19680_));
 sky130_fd_sc_hd__a2111o_2 _24240_ (.A1(_19668_),
    .A2(_19680_),
    .B1(_18542_),
    .C1(alu_wait),
    .D1(_17056_),
    .X(_19681_));
 sky130_fd_sc_hd__o31ai_2 _24241_ (.A1(_17093_),
    .A2(_00302_),
    .A3(_19647_),
    .B1(_19681_),
    .Y(_19682_));
 sky130_fd_sc_hd__nand3b_2 _24242_ (.A_N(_19612_),
    .B(_17119_),
    .C(_19563_),
    .Y(_19683_));
 sky130_fd_sc_hd__a41oi_2 _24243_ (.A1(_19609_),
    .A2(_19673_),
    .A3(_19590_),
    .A4(_19683_),
    .B1(_19529_),
    .Y(_19684_));
 sky130_fd_sc_hd__a2111oi_2 _24244_ (.A1(_19680_),
    .A2(_19638_),
    .B1(_17189_),
    .C1(_19526_),
    .D1(_00310_),
    .Y(_19685_));
 sky130_fd_sc_hd__nand3_2 _24245_ (.A(_19527_),
    .B(_17803_),
    .C(_19564_),
    .Y(_19686_));
 sky130_fd_sc_hd__o2111ai_2 _24246_ (.A1(_19607_),
    .A2(_19569_),
    .B1(_17057_),
    .C1(_17071_),
    .D1(_17068_),
    .Y(_19687_));
 sky130_fd_sc_hd__a21oi_2 _24247_ (.A1(_19686_),
    .A2(_19687_),
    .B1(_00307_),
    .Y(_19688_));
 sky130_fd_sc_hd__a2111o_2 _24248_ (.A1(_19679_),
    .A2(_19682_),
    .B1(_19684_),
    .C1(_19685_),
    .D1(_19688_),
    .X(_00042_));
 sky130_vsdinv _24249_ (.A(_19565_),
    .Y(_00308_));
 sky130_fd_sc_hd__xnor2_2 _24250_ (.A(_18452_),
    .B(_19119_),
    .Y(_19689_));
 sky130_fd_sc_hd__inv_2 _24251_ (.A(_19689_),
    .Y(_02591_));
 sky130_fd_sc_hd__xor2_2 _24252_ (.A(pcpi_rs2[23]),
    .B(_19056_),
    .X(_19690_));
 sky130_fd_sc_hd__xor2_2 _24253_ (.A(pcpi_rs2[20]),
    .B(_19063_),
    .X(_19691_));
 sky130_fd_sc_hd__xor2_2 _24254_ (.A(pcpi_rs2[21]),
    .B(_19061_),
    .X(_19692_));
 sky130_fd_sc_hd__xor2_2 _24255_ (.A(pcpi_rs2[22]),
    .B(_19059_),
    .X(_19693_));
 sky130_fd_sc_hd__or4_2 _24256_ (.A(_19690_),
    .B(_19691_),
    .C(_19692_),
    .D(_19693_),
    .X(_19694_));
 sky130_fd_sc_hd__xor2_2 _24257_ (.A(_18406_),
    .B(_19065_),
    .X(_19695_));
 sky130_fd_sc_hd__xor2_2 _24258_ (.A(pcpi_rs2[16]),
    .B(_19074_),
    .X(_19696_));
 sky130_fd_sc_hd__xor2_2 _24259_ (.A(pcpi_rs2[17]),
    .B(_19071_),
    .X(_19697_));
 sky130_fd_sc_hd__xor2_2 _24260_ (.A(pcpi_rs2[18]),
    .B(_19068_),
    .X(_19698_));
 sky130_fd_sc_hd__or4_2 _24261_ (.A(_19695_),
    .B(_19696_),
    .C(_19697_),
    .D(_19698_),
    .X(_19699_));
 sky130_fd_sc_hd__xor2_2 _24262_ (.A(pcpi_rs2[27]),
    .B(pcpi_rs1[27]),
    .X(_19700_));
 sky130_fd_sc_hd__buf_1 _24263_ (.A(pcpi_rs1[26]),
    .X(_19701_));
 sky130_fd_sc_hd__xor2_2 _24264_ (.A(pcpi_rs2[26]),
    .B(_19701_),
    .X(_19702_));
 sky130_fd_sc_hd__buf_1 _24265_ (.A(pcpi_rs1[24]),
    .X(_19703_));
 sky130_fd_sc_hd__nor2_2 _24266_ (.A(_18396_),
    .B(_19703_),
    .Y(_19704_));
 sky130_fd_sc_hd__and2_2 _24267_ (.A(pcpi_rs2[24]),
    .B(pcpi_rs1[24]),
    .X(_19705_));
 sky130_fd_sc_hd__nor2_2 _24268_ (.A(pcpi_rs2[25]),
    .B(_19052_),
    .Y(_19706_));
 sky130_fd_sc_hd__and2_2 _24269_ (.A(pcpi_rs2[25]),
    .B(pcpi_rs1[25]),
    .X(_19707_));
 sky130_fd_sc_hd__o22ai_2 _24270_ (.A1(_19704_),
    .A2(_19705_),
    .B1(_19706_),
    .B2(_19707_),
    .Y(_19708_));
 sky130_fd_sc_hd__nor2_2 _24271_ (.A(pcpi_rs2[30]),
    .B(pcpi_rs1[30]),
    .Y(_19709_));
 sky130_fd_sc_hd__and2_2 _24272_ (.A(pcpi_rs2[30]),
    .B(pcpi_rs1[30]),
    .X(_19710_));
 sky130_fd_sc_hd__xor2_2 _24273_ (.A(pcpi_rs1[31]),
    .B(pcpi_rs2[31]),
    .X(_19711_));
 sky130_vsdinv _24274_ (.A(_19711_),
    .Y(_19712_));
 sky130_fd_sc_hd__and2_2 _24275_ (.A(pcpi_rs2[29]),
    .B(pcpi_rs1[29]),
    .X(_19713_));
 sky130_fd_sc_hd__nor2_2 _24276_ (.A(pcpi_rs2[29]),
    .B(pcpi_rs1[29]),
    .Y(_19714_));
 sky130_fd_sc_hd__inv_2 _24277_ (.A(pcpi_rs2[28]),
    .Y(_02399_));
 sky130_vsdinv _24278_ (.A(pcpi_rs1[28]),
    .Y(_19715_));
 sky130_fd_sc_hd__nand2_2 _24279_ (.A(_02399_),
    .B(_19715_),
    .Y(_19716_));
 sky130_fd_sc_hd__nand2_2 _24280_ (.A(pcpi_rs2[28]),
    .B(pcpi_rs1[28]),
    .Y(_19717_));
 sky130_fd_sc_hd__a2bb2oi_2 _24281_ (.A1_N(_19713_),
    .A2_N(_19714_),
    .B1(_19716_),
    .B2(_19717_),
    .Y(_19718_));
 sky130_fd_sc_hd__o211ai_2 _24282_ (.A1(_19709_),
    .A2(_19710_),
    .B1(_19712_),
    .C1(_19718_),
    .Y(_19719_));
 sky130_fd_sc_hd__or4_2 _24283_ (.A(_19700_),
    .B(_19702_),
    .C(_19708_),
    .D(_19719_),
    .X(_19720_));
 sky130_fd_sc_hd__nor3_2 _24284_ (.A(_19694_),
    .B(_19699_),
    .C(_19720_),
    .Y(_19721_));
 sky130_fd_sc_hd__xor2_2 _24285_ (.A(pcpi_rs2[15]),
    .B(_19076_),
    .X(_19722_));
 sky130_fd_sc_hd__xor2_2 _24286_ (.A(pcpi_rs2[12]),
    .B(_19084_),
    .X(_19723_));
 sky130_fd_sc_hd__xor2_2 _24287_ (.A(pcpi_rs2[13]),
    .B(_19082_),
    .X(_19724_));
 sky130_fd_sc_hd__xor2_2 _24288_ (.A(pcpi_rs2[14]),
    .B(_19080_),
    .X(_19725_));
 sky130_fd_sc_hd__or4_2 _24289_ (.A(_19722_),
    .B(_19723_),
    .C(_19724_),
    .D(_19725_),
    .X(_19726_));
 sky130_fd_sc_hd__xnor2_2 _24290_ (.A(mem_la_wdata[3]),
    .B(_19109_),
    .Y(_19727_));
 sky130_vsdinv _24291_ (.A(_19112_),
    .Y(_19728_));
 sky130_fd_sc_hd__nand2_2 _24292_ (.A(_19539_),
    .B(_19728_),
    .Y(_19729_));
 sky130_fd_sc_hd__nand2_2 _24293_ (.A(_18447_),
    .B(_19112_),
    .Y(_19730_));
 sky130_fd_sc_hd__nand2_2 _24294_ (.A(_19729_),
    .B(_19730_),
    .Y(_19731_));
 sky130_fd_sc_hd__nand2_2 _24295_ (.A(_19727_),
    .B(_19731_),
    .Y(_19732_));
 sky130_fd_sc_hd__nor2_2 _24296_ (.A(_18441_),
    .B(_19107_),
    .Y(_19733_));
 sky130_fd_sc_hd__and2_2 _24297_ (.A(mem_la_wdata[4]),
    .B(_19106_),
    .X(_19734_));
 sky130_fd_sc_hd__nor2_2 _24298_ (.A(_18438_),
    .B(_19104_),
    .Y(_19735_));
 sky130_fd_sc_hd__and2_2 _24299_ (.A(_18438_),
    .B(_19104_),
    .X(_19736_));
 sky130_fd_sc_hd__o22ai_2 _24300_ (.A1(_19733_),
    .A2(_19734_),
    .B1(_19735_),
    .B2(_19736_),
    .Y(_19737_));
 sky130_fd_sc_hd__inv_2 _24301_ (.A(_18435_),
    .Y(_02333_));
 sky130_vsdinv _24302_ (.A(_19102_),
    .Y(_19738_));
 sky130_fd_sc_hd__nand2_2 _24303_ (.A(_02333_),
    .B(_19738_),
    .Y(_19739_));
 sky130_fd_sc_hd__nand2_2 _24304_ (.A(_18435_),
    .B(_19102_),
    .Y(_19740_));
 sky130_fd_sc_hd__xor2_2 _24305_ (.A(_18449_),
    .B(_19115_),
    .X(_19741_));
 sky130_fd_sc_hd__xor2_2 _24306_ (.A(_18432_),
    .B(_19098_),
    .X(_19742_));
 sky130_fd_sc_hd__a2111o_2 _24307_ (.A1(_19739_),
    .A2(_19740_),
    .B1(_19741_),
    .C1(_19742_),
    .D1(_02591_),
    .X(_19743_));
 sky130_fd_sc_hd__nor3_2 _24308_ (.A(_19732_),
    .B(_19737_),
    .C(_19743_),
    .Y(_19744_));
 sky130_fd_sc_hd__nor2_2 _24309_ (.A(_18429_),
    .B(_19095_),
    .Y(_19745_));
 sky130_fd_sc_hd__and2_2 _24310_ (.A(_18429_),
    .B(_19095_),
    .X(_19746_));
 sky130_fd_sc_hd__xnor2_2 _24311_ (.A(pcpi_rs2[9]),
    .B(_19092_),
    .Y(_19747_));
 sky130_fd_sc_hd__nor2_2 _24312_ (.A(_18423_),
    .B(_19086_),
    .Y(_19748_));
 sky130_fd_sc_hd__and2_2 _24313_ (.A(pcpi_rs2[11]),
    .B(_19086_),
    .X(_19749_));
 sky130_fd_sc_hd__nor2_2 _24314_ (.A(_19748_),
    .B(_19749_),
    .Y(_19750_));
 sky130_vsdinv _24315_ (.A(_19750_),
    .Y(_19751_));
 sky130_fd_sc_hd__xor2_2 _24316_ (.A(pcpi_rs2[10]),
    .B(_19089_),
    .X(_19752_));
 sky130_vsdinv _24317_ (.A(_19752_),
    .Y(_19753_));
 sky130_fd_sc_hd__o2111a_2 _24318_ (.A1(_19745_),
    .A2(_19746_),
    .B1(_19747_),
    .C1(_19751_),
    .D1(_19753_),
    .X(_19754_));
 sky130_fd_sc_hd__and3b_2 _24319_ (.A_N(_19726_),
    .B(_19744_),
    .C(_19754_),
    .X(_19755_));
 sky130_fd_sc_hd__and2_2 _24320_ (.A(_19721_),
    .B(_19755_),
    .X(_19756_));
 sky130_fd_sc_hd__buf_1 _24321_ (.A(_19756_),
    .X(_00000_));
 sky130_fd_sc_hd__o211a_2 _24322_ (.A1(_16938_),
    .A2(pcpi_insn[12]),
    .B1(_16948_),
    .C1(_16944_),
    .X(\pcpi_mul.instr_any_mulh ));
 sky130_fd_sc_hd__or3_2 _24323_ (.A(instr_slt),
    .B(instr_slti),
    .C(instr_blt),
    .X(_00006_));
 sky130_fd_sc_hd__or3_2 _24324_ (.A(instr_sltu),
    .B(instr_sltiu),
    .C(instr_bltu),
    .X(_00007_));
 sky130_fd_sc_hd__a211o_2 _24325_ (.A1(_18005_),
    .A2(_16800_),
    .B1(_16836_),
    .C1(_18001_),
    .X(_00299_));
 sky130_fd_sc_hd__buf_1 _24326_ (.A(_19667_),
    .X(_19757_));
 sky130_fd_sc_hd__buf_1 _24327_ (.A(_19757_),
    .X(_19758_));
 sky130_fd_sc_hd__buf_1 _24328_ (.A(_16821_),
    .X(_19759_));
 sky130_fd_sc_hd__nor3_2 _24329_ (.A(_17393_),
    .B(_19759_),
    .C(_19664_),
    .Y(_19760_));
 sky130_fd_sc_hd__o21ba_2 _24330_ (.A1(_00319_),
    .A2(_00317_),
    .B1_N(_17387_),
    .X(_19761_));
 sky130_fd_sc_hd__a2111o_2 _24331_ (.A1(_19633_),
    .A2(_19663_),
    .B1(_17048_),
    .C1(_19760_),
    .D1(_19761_),
    .X(_19762_));
 sky130_fd_sc_hd__buf_1 _24332_ (.A(_16849_),
    .X(_19763_));
 sky130_fd_sc_hd__o2111ai_2 _24333_ (.A1(instr_lhu),
    .A2(instr_lh),
    .B1(_17803_),
    .C1(_19763_),
    .D1(_17389_),
    .Y(_19764_));
 sky130_fd_sc_hd__o41a_2 _24334_ (.A1(_17218_),
    .A2(_17148_),
    .A3(_19011_),
    .A4(_18030_),
    .B1(_19764_),
    .X(_19765_));
 sky130_fd_sc_hd__o2bb2ai_2 _24335_ (.A1_N(_19758_),
    .A2_N(_19762_),
    .B1(_00296_),
    .B2(_19765_),
    .Y(_00047_));
 sky130_fd_sc_hd__buf_1 _24336_ (.A(_16847_),
    .X(_00301_));
 sky130_fd_sc_hd__buf_1 _24337_ (.A(_19517_),
    .X(_19766_));
 sky130_fd_sc_hd__nor3_2 _24338_ (.A(_19766_),
    .B(_17390_),
    .C(_19664_),
    .Y(_00336_));
 sky130_fd_sc_hd__a211o_2 _24339_ (.A1(_16858_),
    .A2(_17081_),
    .B1(_17211_),
    .C1(_17386_),
    .X(_00338_));
 sky130_fd_sc_hd__inv_2 _24340_ (.A(alu_eq),
    .Y(_00340_));
 sky130_fd_sc_hd__nor3_2 _24341_ (.A(instr_bne),
    .B(is_slti_blt_slt),
    .C(is_sltiu_bltu_sltu),
    .Y(_19767_));
 sky130_fd_sc_hd__and2_2 _24342_ (.A(_19767_),
    .B(_17012_),
    .X(_00341_));
 sky130_fd_sc_hd__and2b_2 _24343_ (.A_N(alu_lts),
    .B(instr_bge),
    .X(_19768_));
 sky130_fd_sc_hd__and2b_2 _24344_ (.A_N(alu_ltu),
    .B(instr_bgeu),
    .X(_19769_));
 sky130_fd_sc_hd__a221o_2 _24345_ (.A1(is_slti_blt_slt),
    .A2(alu_lts),
    .B1(is_sltiu_bltu_sltu),
    .B2(alu_ltu),
    .C1(_19769_),
    .X(_19770_));
 sky130_fd_sc_hd__a211oi_2 _24346_ (.A1(instr_bne),
    .A2(_00340_),
    .B1(_19768_),
    .C1(_19770_),
    .Y(_00342_));
 sky130_fd_sc_hd__nand2_2 _24347_ (.A(_19783_),
    .B(_00343_),
    .Y(_00344_));
 sky130_fd_sc_hd__buf_1 _24348_ (.A(_16984_),
    .X(_19771_));
 sky130_fd_sc_hd__o22ai_2 _24349_ (.A1(_00346_),
    .A2(_19771_),
    .B1(_00339_),
    .B2(_00297_),
    .Y(_00347_));
 sky130_fd_sc_hd__buf_1 _24350_ (.A(_17037_),
    .X(_19772_));
 sky130_fd_sc_hd__o21ba_2 _24351_ (.A1(_17361_),
    .A2(do_waitirq),
    .B1_N(_19772_),
    .X(_00349_));
 sky130_fd_sc_hd__nor3b_2 _24352_ (.A(_18014_),
    .B(_18019_),
    .C_N(_00349_),
    .Y(_00351_));
 sky130_fd_sc_hd__buf_1 _24353_ (.A(_17966_),
    .X(_19773_));
 sky130_fd_sc_hd__buf_1 _24354_ (.A(_19661_),
    .X(_19774_));
 sky130_fd_sc_hd__nor3_2 _24355_ (.A(_19766_),
    .B(_19773_),
    .C(_19774_),
    .Y(_00354_));
 sky130_fd_sc_hd__a211oi_2 _24356_ (.A1(_19766_),
    .A2(_17081_),
    .B1(_19773_),
    .C1(_19774_),
    .Y(_00355_));
 sky130_fd_sc_hd__inv_2 _24357_ (.A(\decoded_imm_uj[4] ),
    .Y(_00367_));
 sky130_vsdinv _24358_ (.A(\cpuregs[0][1] ),
    .Y(_00371_));
 sky130_vsdinv _24359_ (.A(\cpuregs[1][1] ),
    .Y(_00372_));
 sky130_vsdinv _24360_ (.A(\cpuregs[2][1] ),
    .Y(_00373_));
 sky130_vsdinv _24361_ (.A(\cpuregs[3][1] ),
    .Y(_00374_));
 sky130_vsdinv _24362_ (.A(\cpuregs[4][1] ),
    .Y(_00376_));
 sky130_vsdinv _24363_ (.A(\cpuregs[5][1] ),
    .Y(_00377_));
 sky130_vsdinv _24364_ (.A(\cpuregs[6][1] ),
    .Y(_00378_));
 sky130_vsdinv _24365_ (.A(\cpuregs[7][1] ),
    .Y(_00379_));
 sky130_vsdinv _24366_ (.A(\cpuregs[8][1] ),
    .Y(_00381_));
 sky130_vsdinv _24367_ (.A(\cpuregs[9][1] ),
    .Y(_00382_));
 sky130_vsdinv _24368_ (.A(\cpuregs[10][1] ),
    .Y(_00383_));
 sky130_vsdinv _24369_ (.A(\cpuregs[11][1] ),
    .Y(_00384_));
 sky130_vsdinv _24370_ (.A(\cpuregs[12][1] ),
    .Y(_00386_));
 sky130_vsdinv _24371_ (.A(\cpuregs[13][1] ),
    .Y(_00387_));
 sky130_vsdinv _24372_ (.A(\cpuregs[14][1] ),
    .Y(_00388_));
 sky130_vsdinv _24373_ (.A(\cpuregs[15][1] ),
    .Y(_00389_));
 sky130_vsdinv _24374_ (.A(\cpuregs[16][1] ),
    .Y(_00392_));
 sky130_vsdinv _24375_ (.A(\cpuregs[17][1] ),
    .Y(_00393_));
 sky130_vsdinv _24376_ (.A(\cpuregs[18][1] ),
    .Y(_00394_));
 sky130_vsdinv _24377_ (.A(\cpuregs[19][1] ),
    .Y(_00395_));
 sky130_vsdinv _24378_ (.A(\cpuregs[0][2] ),
    .Y(_00398_));
 sky130_vsdinv _24379_ (.A(\cpuregs[1][2] ),
    .Y(_00399_));
 sky130_vsdinv _24380_ (.A(\cpuregs[2][2] ),
    .Y(_00400_));
 sky130_vsdinv _24381_ (.A(\cpuregs[3][2] ),
    .Y(_00401_));
 sky130_vsdinv _24382_ (.A(\cpuregs[4][2] ),
    .Y(_00403_));
 sky130_vsdinv _24383_ (.A(\cpuregs[5][2] ),
    .Y(_00404_));
 sky130_vsdinv _24384_ (.A(\cpuregs[6][2] ),
    .Y(_00405_));
 sky130_vsdinv _24385_ (.A(\cpuregs[7][2] ),
    .Y(_00406_));
 sky130_vsdinv _24386_ (.A(\cpuregs[8][2] ),
    .Y(_00408_));
 sky130_vsdinv _24387_ (.A(\cpuregs[9][2] ),
    .Y(_00409_));
 sky130_vsdinv _24388_ (.A(\cpuregs[10][2] ),
    .Y(_00410_));
 sky130_vsdinv _24389_ (.A(\cpuregs[11][2] ),
    .Y(_00411_));
 sky130_vsdinv _24390_ (.A(\cpuregs[12][2] ),
    .Y(_00413_));
 sky130_vsdinv _24391_ (.A(\cpuregs[13][2] ),
    .Y(_00414_));
 sky130_vsdinv _24392_ (.A(\cpuregs[14][2] ),
    .Y(_00415_));
 sky130_vsdinv _24393_ (.A(\cpuregs[15][2] ),
    .Y(_00416_));
 sky130_vsdinv _24394_ (.A(\cpuregs[16][2] ),
    .Y(_00419_));
 sky130_vsdinv _24395_ (.A(\cpuregs[17][2] ),
    .Y(_00420_));
 sky130_vsdinv _24396_ (.A(\cpuregs[18][2] ),
    .Y(_00421_));
 sky130_vsdinv _24397_ (.A(\cpuregs[19][2] ),
    .Y(_00422_));
 sky130_vsdinv _24398_ (.A(\cpuregs[0][3] ),
    .Y(_00425_));
 sky130_vsdinv _24399_ (.A(\cpuregs[1][3] ),
    .Y(_00426_));
 sky130_vsdinv _24400_ (.A(\cpuregs[2][3] ),
    .Y(_00427_));
 sky130_vsdinv _24401_ (.A(\cpuregs[3][3] ),
    .Y(_00428_));
 sky130_vsdinv _24402_ (.A(\cpuregs[4][3] ),
    .Y(_00430_));
 sky130_vsdinv _24403_ (.A(\cpuregs[5][3] ),
    .Y(_00431_));
 sky130_vsdinv _24404_ (.A(\cpuregs[6][3] ),
    .Y(_00432_));
 sky130_vsdinv _24405_ (.A(\cpuregs[7][3] ),
    .Y(_00433_));
 sky130_vsdinv _24406_ (.A(\cpuregs[8][3] ),
    .Y(_00435_));
 sky130_vsdinv _24407_ (.A(\cpuregs[9][3] ),
    .Y(_00436_));
 sky130_vsdinv _24408_ (.A(\cpuregs[10][3] ),
    .Y(_00437_));
 sky130_vsdinv _24409_ (.A(\cpuregs[11][3] ),
    .Y(_00438_));
 sky130_vsdinv _24410_ (.A(\cpuregs[12][3] ),
    .Y(_00440_));
 sky130_vsdinv _24411_ (.A(\cpuregs[13][3] ),
    .Y(_00441_));
 sky130_vsdinv _24412_ (.A(\cpuregs[14][3] ),
    .Y(_00442_));
 sky130_vsdinv _24413_ (.A(\cpuregs[15][3] ),
    .Y(_00443_));
 sky130_vsdinv _24414_ (.A(\cpuregs[16][3] ),
    .Y(_00446_));
 sky130_vsdinv _24415_ (.A(\cpuregs[17][3] ),
    .Y(_00447_));
 sky130_vsdinv _24416_ (.A(\cpuregs[18][3] ),
    .Y(_00448_));
 sky130_vsdinv _24417_ (.A(\cpuregs[19][3] ),
    .Y(_00449_));
 sky130_vsdinv _24418_ (.A(\cpuregs[0][4] ),
    .Y(_00452_));
 sky130_vsdinv _24419_ (.A(\cpuregs[1][4] ),
    .Y(_00453_));
 sky130_vsdinv _24420_ (.A(\cpuregs[2][4] ),
    .Y(_00454_));
 sky130_vsdinv _24421_ (.A(\cpuregs[3][4] ),
    .Y(_00455_));
 sky130_vsdinv _24422_ (.A(\cpuregs[4][4] ),
    .Y(_00457_));
 sky130_vsdinv _24423_ (.A(\cpuregs[5][4] ),
    .Y(_00458_));
 sky130_vsdinv _24424_ (.A(\cpuregs[6][4] ),
    .Y(_00459_));
 sky130_vsdinv _24425_ (.A(\cpuregs[7][4] ),
    .Y(_00460_));
 sky130_vsdinv _24426_ (.A(\cpuregs[8][4] ),
    .Y(_00462_));
 sky130_vsdinv _24427_ (.A(\cpuregs[9][4] ),
    .Y(_00463_));
 sky130_vsdinv _24428_ (.A(\cpuregs[10][4] ),
    .Y(_00464_));
 sky130_vsdinv _24429_ (.A(\cpuregs[11][4] ),
    .Y(_00465_));
 sky130_vsdinv _24430_ (.A(\cpuregs[12][4] ),
    .Y(_00467_));
 sky130_vsdinv _24431_ (.A(\cpuregs[13][4] ),
    .Y(_00468_));
 sky130_vsdinv _24432_ (.A(\cpuregs[14][4] ),
    .Y(_00469_));
 sky130_vsdinv _24433_ (.A(\cpuregs[15][4] ),
    .Y(_00470_));
 sky130_vsdinv _24434_ (.A(\cpuregs[16][4] ),
    .Y(_00473_));
 sky130_vsdinv _24435_ (.A(\cpuregs[17][4] ),
    .Y(_00474_));
 sky130_vsdinv _24436_ (.A(\cpuregs[18][4] ),
    .Y(_00475_));
 sky130_vsdinv _24437_ (.A(\cpuregs[19][4] ),
    .Y(_00476_));
 sky130_vsdinv _24438_ (.A(\cpuregs[0][5] ),
    .Y(_00479_));
 sky130_vsdinv _24439_ (.A(\cpuregs[1][5] ),
    .Y(_00480_));
 sky130_vsdinv _24440_ (.A(\cpuregs[2][5] ),
    .Y(_00481_));
 sky130_vsdinv _24441_ (.A(\cpuregs[3][5] ),
    .Y(_00482_));
 sky130_vsdinv _24442_ (.A(\cpuregs[4][5] ),
    .Y(_00484_));
 sky130_vsdinv _24443_ (.A(\cpuregs[5][5] ),
    .Y(_00485_));
 sky130_vsdinv _24444_ (.A(\cpuregs[6][5] ),
    .Y(_00486_));
 sky130_vsdinv _24445_ (.A(\cpuregs[7][5] ),
    .Y(_00487_));
 sky130_vsdinv _24446_ (.A(\cpuregs[8][5] ),
    .Y(_00489_));
 sky130_vsdinv _24447_ (.A(\cpuregs[9][5] ),
    .Y(_00490_));
 sky130_vsdinv _24448_ (.A(\cpuregs[10][5] ),
    .Y(_00491_));
 sky130_vsdinv _24449_ (.A(\cpuregs[11][5] ),
    .Y(_00492_));
 sky130_vsdinv _24450_ (.A(\cpuregs[12][5] ),
    .Y(_00494_));
 sky130_vsdinv _24451_ (.A(\cpuregs[13][5] ),
    .Y(_00495_));
 sky130_vsdinv _24452_ (.A(\cpuregs[14][5] ),
    .Y(_00496_));
 sky130_vsdinv _24453_ (.A(\cpuregs[15][5] ),
    .Y(_00497_));
 sky130_vsdinv _24454_ (.A(\cpuregs[16][5] ),
    .Y(_00500_));
 sky130_vsdinv _24455_ (.A(\cpuregs[17][5] ),
    .Y(_00501_));
 sky130_vsdinv _24456_ (.A(\cpuregs[18][5] ),
    .Y(_00502_));
 sky130_vsdinv _24457_ (.A(\cpuregs[19][5] ),
    .Y(_00503_));
 sky130_vsdinv _24458_ (.A(\cpuregs[0][6] ),
    .Y(_00506_));
 sky130_vsdinv _24459_ (.A(\cpuregs[1][6] ),
    .Y(_00507_));
 sky130_vsdinv _24460_ (.A(\cpuregs[2][6] ),
    .Y(_00508_));
 sky130_vsdinv _24461_ (.A(\cpuregs[3][6] ),
    .Y(_00509_));
 sky130_vsdinv _24462_ (.A(\cpuregs[4][6] ),
    .Y(_00511_));
 sky130_vsdinv _24463_ (.A(\cpuregs[5][6] ),
    .Y(_00512_));
 sky130_vsdinv _24464_ (.A(\cpuregs[6][6] ),
    .Y(_00513_));
 sky130_vsdinv _24465_ (.A(\cpuregs[7][6] ),
    .Y(_00514_));
 sky130_vsdinv _24466_ (.A(\cpuregs[8][6] ),
    .Y(_00516_));
 sky130_vsdinv _24467_ (.A(\cpuregs[9][6] ),
    .Y(_00517_));
 sky130_vsdinv _24468_ (.A(\cpuregs[10][6] ),
    .Y(_00518_));
 sky130_vsdinv _24469_ (.A(\cpuregs[11][6] ),
    .Y(_00519_));
 sky130_vsdinv _24470_ (.A(\cpuregs[12][6] ),
    .Y(_00521_));
 sky130_vsdinv _24471_ (.A(\cpuregs[13][6] ),
    .Y(_00522_));
 sky130_vsdinv _24472_ (.A(\cpuregs[14][6] ),
    .Y(_00523_));
 sky130_vsdinv _24473_ (.A(\cpuregs[15][6] ),
    .Y(_00524_));
 sky130_vsdinv _24474_ (.A(\cpuregs[16][6] ),
    .Y(_00527_));
 sky130_vsdinv _24475_ (.A(\cpuregs[17][6] ),
    .Y(_00528_));
 sky130_vsdinv _24476_ (.A(\cpuregs[18][6] ),
    .Y(_00529_));
 sky130_vsdinv _24477_ (.A(\cpuregs[19][6] ),
    .Y(_00530_));
 sky130_vsdinv _24478_ (.A(\cpuregs[0][7] ),
    .Y(_00533_));
 sky130_vsdinv _24479_ (.A(\cpuregs[1][7] ),
    .Y(_00534_));
 sky130_vsdinv _24480_ (.A(\cpuregs[2][7] ),
    .Y(_00535_));
 sky130_vsdinv _24481_ (.A(\cpuregs[3][7] ),
    .Y(_00536_));
 sky130_vsdinv _24482_ (.A(\cpuregs[4][7] ),
    .Y(_00538_));
 sky130_vsdinv _24483_ (.A(\cpuregs[5][7] ),
    .Y(_00539_));
 sky130_vsdinv _24484_ (.A(\cpuregs[6][7] ),
    .Y(_00540_));
 sky130_vsdinv _24485_ (.A(\cpuregs[7][7] ),
    .Y(_00541_));
 sky130_vsdinv _24486_ (.A(\cpuregs[8][7] ),
    .Y(_00543_));
 sky130_vsdinv _24487_ (.A(\cpuregs[9][7] ),
    .Y(_00544_));
 sky130_vsdinv _24488_ (.A(\cpuregs[10][7] ),
    .Y(_00545_));
 sky130_vsdinv _24489_ (.A(\cpuregs[11][7] ),
    .Y(_00546_));
 sky130_vsdinv _24490_ (.A(\cpuregs[12][7] ),
    .Y(_00548_));
 sky130_vsdinv _24491_ (.A(\cpuregs[13][7] ),
    .Y(_00549_));
 sky130_vsdinv _24492_ (.A(\cpuregs[14][7] ),
    .Y(_00550_));
 sky130_vsdinv _24493_ (.A(\cpuregs[15][7] ),
    .Y(_00551_));
 sky130_vsdinv _24494_ (.A(\cpuregs[16][7] ),
    .Y(_00554_));
 sky130_vsdinv _24495_ (.A(\cpuregs[17][7] ),
    .Y(_00555_));
 sky130_vsdinv _24496_ (.A(\cpuregs[18][7] ),
    .Y(_00556_));
 sky130_vsdinv _24497_ (.A(\cpuregs[19][7] ),
    .Y(_00557_));
 sky130_vsdinv _24498_ (.A(\cpuregs[0][8] ),
    .Y(_00560_));
 sky130_vsdinv _24499_ (.A(\cpuregs[1][8] ),
    .Y(_00561_));
 sky130_vsdinv _24500_ (.A(\cpuregs[2][8] ),
    .Y(_00562_));
 sky130_vsdinv _24501_ (.A(\cpuregs[3][8] ),
    .Y(_00563_));
 sky130_vsdinv _24502_ (.A(\cpuregs[4][8] ),
    .Y(_00565_));
 sky130_vsdinv _24503_ (.A(\cpuregs[5][8] ),
    .Y(_00566_));
 sky130_vsdinv _24504_ (.A(\cpuregs[6][8] ),
    .Y(_00567_));
 sky130_vsdinv _24505_ (.A(\cpuregs[7][8] ),
    .Y(_00568_));
 sky130_vsdinv _24506_ (.A(\cpuregs[8][8] ),
    .Y(_00570_));
 sky130_vsdinv _24507_ (.A(\cpuregs[9][8] ),
    .Y(_00571_));
 sky130_vsdinv _24508_ (.A(\cpuregs[10][8] ),
    .Y(_00572_));
 sky130_vsdinv _24509_ (.A(\cpuregs[11][8] ),
    .Y(_00573_));
 sky130_vsdinv _24510_ (.A(\cpuregs[12][8] ),
    .Y(_00575_));
 sky130_vsdinv _24511_ (.A(\cpuregs[13][8] ),
    .Y(_00576_));
 sky130_vsdinv _24512_ (.A(\cpuregs[14][8] ),
    .Y(_00577_));
 sky130_vsdinv _24513_ (.A(\cpuregs[15][8] ),
    .Y(_00578_));
 sky130_vsdinv _24514_ (.A(\cpuregs[16][8] ),
    .Y(_00581_));
 sky130_vsdinv _24515_ (.A(\cpuregs[17][8] ),
    .Y(_00582_));
 sky130_vsdinv _24516_ (.A(\cpuregs[18][8] ),
    .Y(_00583_));
 sky130_vsdinv _24517_ (.A(\cpuregs[19][8] ),
    .Y(_00584_));
 sky130_vsdinv _24518_ (.A(\cpuregs[0][9] ),
    .Y(_00587_));
 sky130_vsdinv _24519_ (.A(\cpuregs[1][9] ),
    .Y(_00588_));
 sky130_vsdinv _24520_ (.A(\cpuregs[2][9] ),
    .Y(_00589_));
 sky130_vsdinv _24521_ (.A(\cpuregs[3][9] ),
    .Y(_00590_));
 sky130_vsdinv _24522_ (.A(\cpuregs[4][9] ),
    .Y(_00592_));
 sky130_vsdinv _24523_ (.A(\cpuregs[5][9] ),
    .Y(_00593_));
 sky130_vsdinv _24524_ (.A(\cpuregs[6][9] ),
    .Y(_00594_));
 sky130_vsdinv _24525_ (.A(\cpuregs[7][9] ),
    .Y(_00595_));
 sky130_vsdinv _24526_ (.A(\cpuregs[8][9] ),
    .Y(_00597_));
 sky130_vsdinv _24527_ (.A(\cpuregs[9][9] ),
    .Y(_00598_));
 sky130_vsdinv _24528_ (.A(\cpuregs[10][9] ),
    .Y(_00599_));
 sky130_vsdinv _24529_ (.A(\cpuregs[11][9] ),
    .Y(_00600_));
 sky130_vsdinv _24530_ (.A(\cpuregs[12][9] ),
    .Y(_00602_));
 sky130_vsdinv _24531_ (.A(\cpuregs[13][9] ),
    .Y(_00603_));
 sky130_vsdinv _24532_ (.A(\cpuregs[14][9] ),
    .Y(_00604_));
 sky130_vsdinv _24533_ (.A(\cpuregs[15][9] ),
    .Y(_00605_));
 sky130_vsdinv _24534_ (.A(\cpuregs[16][9] ),
    .Y(_00608_));
 sky130_vsdinv _24535_ (.A(\cpuregs[17][9] ),
    .Y(_00609_));
 sky130_vsdinv _24536_ (.A(\cpuregs[18][9] ),
    .Y(_00610_));
 sky130_vsdinv _24537_ (.A(\cpuregs[19][9] ),
    .Y(_00611_));
 sky130_vsdinv _24538_ (.A(\cpuregs[0][10] ),
    .Y(_00614_));
 sky130_vsdinv _24539_ (.A(\cpuregs[1][10] ),
    .Y(_00615_));
 sky130_vsdinv _24540_ (.A(\cpuregs[2][10] ),
    .Y(_00616_));
 sky130_vsdinv _24541_ (.A(\cpuregs[3][10] ),
    .Y(_00617_));
 sky130_vsdinv _24542_ (.A(\cpuregs[4][10] ),
    .Y(_00619_));
 sky130_vsdinv _24543_ (.A(\cpuregs[5][10] ),
    .Y(_00620_));
 sky130_vsdinv _24544_ (.A(\cpuregs[6][10] ),
    .Y(_00621_));
 sky130_vsdinv _24545_ (.A(\cpuregs[7][10] ),
    .Y(_00622_));
 sky130_vsdinv _24546_ (.A(\cpuregs[8][10] ),
    .Y(_00624_));
 sky130_vsdinv _24547_ (.A(\cpuregs[9][10] ),
    .Y(_00625_));
 sky130_vsdinv _24548_ (.A(\cpuregs[10][10] ),
    .Y(_00626_));
 sky130_vsdinv _24549_ (.A(\cpuregs[11][10] ),
    .Y(_00627_));
 sky130_vsdinv _24550_ (.A(\cpuregs[12][10] ),
    .Y(_00629_));
 sky130_vsdinv _24551_ (.A(\cpuregs[13][10] ),
    .Y(_00630_));
 sky130_vsdinv _24552_ (.A(\cpuregs[14][10] ),
    .Y(_00631_));
 sky130_vsdinv _24553_ (.A(\cpuregs[15][10] ),
    .Y(_00632_));
 sky130_vsdinv _24554_ (.A(\cpuregs[16][10] ),
    .Y(_00635_));
 sky130_vsdinv _24555_ (.A(\cpuregs[17][10] ),
    .Y(_00636_));
 sky130_vsdinv _24556_ (.A(\cpuregs[18][10] ),
    .Y(_00637_));
 sky130_vsdinv _24557_ (.A(\cpuregs[19][10] ),
    .Y(_00638_));
 sky130_vsdinv _24558_ (.A(\cpuregs[0][11] ),
    .Y(_00641_));
 sky130_vsdinv _24559_ (.A(\cpuregs[1][11] ),
    .Y(_00642_));
 sky130_vsdinv _24560_ (.A(\cpuregs[2][11] ),
    .Y(_00643_));
 sky130_vsdinv _24561_ (.A(\cpuregs[3][11] ),
    .Y(_00644_));
 sky130_vsdinv _24562_ (.A(\cpuregs[4][11] ),
    .Y(_00646_));
 sky130_vsdinv _24563_ (.A(\cpuregs[5][11] ),
    .Y(_00647_));
 sky130_vsdinv _24564_ (.A(\cpuregs[6][11] ),
    .Y(_00648_));
 sky130_vsdinv _24565_ (.A(\cpuregs[7][11] ),
    .Y(_00649_));
 sky130_vsdinv _24566_ (.A(\cpuregs[8][11] ),
    .Y(_00651_));
 sky130_vsdinv _24567_ (.A(\cpuregs[9][11] ),
    .Y(_00652_));
 sky130_vsdinv _24568_ (.A(\cpuregs[10][11] ),
    .Y(_00653_));
 sky130_vsdinv _24569_ (.A(\cpuregs[11][11] ),
    .Y(_00654_));
 sky130_vsdinv _24570_ (.A(\cpuregs[12][11] ),
    .Y(_00656_));
 sky130_vsdinv _24571_ (.A(\cpuregs[13][11] ),
    .Y(_00657_));
 sky130_vsdinv _24572_ (.A(\cpuregs[14][11] ),
    .Y(_00658_));
 sky130_vsdinv _24573_ (.A(\cpuregs[15][11] ),
    .Y(_00659_));
 sky130_vsdinv _24574_ (.A(\cpuregs[16][11] ),
    .Y(_00662_));
 sky130_vsdinv _24575_ (.A(\cpuregs[17][11] ),
    .Y(_00663_));
 sky130_vsdinv _24576_ (.A(\cpuregs[18][11] ),
    .Y(_00664_));
 sky130_vsdinv _24577_ (.A(\cpuregs[19][11] ),
    .Y(_00665_));
 sky130_vsdinv _24578_ (.A(\cpuregs[0][12] ),
    .Y(_00668_));
 sky130_vsdinv _24579_ (.A(\cpuregs[1][12] ),
    .Y(_00669_));
 sky130_vsdinv _24580_ (.A(\cpuregs[2][12] ),
    .Y(_00670_));
 sky130_vsdinv _24581_ (.A(\cpuregs[3][12] ),
    .Y(_00671_));
 sky130_vsdinv _24582_ (.A(\cpuregs[4][12] ),
    .Y(_00673_));
 sky130_vsdinv _24583_ (.A(\cpuregs[5][12] ),
    .Y(_00674_));
 sky130_vsdinv _24584_ (.A(\cpuregs[6][12] ),
    .Y(_00675_));
 sky130_vsdinv _24585_ (.A(\cpuregs[7][12] ),
    .Y(_00676_));
 sky130_vsdinv _24586_ (.A(\cpuregs[8][12] ),
    .Y(_00678_));
 sky130_vsdinv _24587_ (.A(\cpuregs[9][12] ),
    .Y(_00679_));
 sky130_vsdinv _24588_ (.A(\cpuregs[10][12] ),
    .Y(_00680_));
 sky130_vsdinv _24589_ (.A(\cpuregs[11][12] ),
    .Y(_00681_));
 sky130_vsdinv _24590_ (.A(\cpuregs[12][12] ),
    .Y(_00683_));
 sky130_vsdinv _24591_ (.A(\cpuregs[13][12] ),
    .Y(_00684_));
 sky130_vsdinv _24592_ (.A(\cpuregs[14][12] ),
    .Y(_00685_));
 sky130_vsdinv _24593_ (.A(\cpuregs[15][12] ),
    .Y(_00686_));
 sky130_vsdinv _24594_ (.A(\cpuregs[16][12] ),
    .Y(_00689_));
 sky130_vsdinv _24595_ (.A(\cpuregs[17][12] ),
    .Y(_00690_));
 sky130_vsdinv _24596_ (.A(\cpuregs[18][12] ),
    .Y(_00691_));
 sky130_vsdinv _24597_ (.A(\cpuregs[19][12] ),
    .Y(_00692_));
 sky130_vsdinv _24598_ (.A(\cpuregs[0][13] ),
    .Y(_00695_));
 sky130_vsdinv _24599_ (.A(\cpuregs[1][13] ),
    .Y(_00696_));
 sky130_vsdinv _24600_ (.A(\cpuregs[2][13] ),
    .Y(_00697_));
 sky130_vsdinv _24601_ (.A(\cpuregs[3][13] ),
    .Y(_00698_));
 sky130_vsdinv _24602_ (.A(\cpuregs[4][13] ),
    .Y(_00700_));
 sky130_vsdinv _24603_ (.A(\cpuregs[5][13] ),
    .Y(_00701_));
 sky130_vsdinv _24604_ (.A(\cpuregs[6][13] ),
    .Y(_00702_));
 sky130_vsdinv _24605_ (.A(\cpuregs[7][13] ),
    .Y(_00703_));
 sky130_vsdinv _24606_ (.A(\cpuregs[8][13] ),
    .Y(_00705_));
 sky130_vsdinv _24607_ (.A(\cpuregs[9][13] ),
    .Y(_00706_));
 sky130_vsdinv _24608_ (.A(\cpuregs[10][13] ),
    .Y(_00707_));
 sky130_vsdinv _24609_ (.A(\cpuregs[11][13] ),
    .Y(_00708_));
 sky130_vsdinv _24610_ (.A(\cpuregs[12][13] ),
    .Y(_00710_));
 sky130_vsdinv _24611_ (.A(\cpuregs[13][13] ),
    .Y(_00711_));
 sky130_vsdinv _24612_ (.A(\cpuregs[14][13] ),
    .Y(_00712_));
 sky130_vsdinv _24613_ (.A(\cpuregs[15][13] ),
    .Y(_00713_));
 sky130_vsdinv _24614_ (.A(\cpuregs[16][13] ),
    .Y(_00716_));
 sky130_vsdinv _24615_ (.A(\cpuregs[17][13] ),
    .Y(_00717_));
 sky130_vsdinv _24616_ (.A(\cpuregs[18][13] ),
    .Y(_00718_));
 sky130_vsdinv _24617_ (.A(\cpuregs[19][13] ),
    .Y(_00719_));
 sky130_vsdinv _24618_ (.A(\cpuregs[0][14] ),
    .Y(_00722_));
 sky130_vsdinv _24619_ (.A(\cpuregs[1][14] ),
    .Y(_00723_));
 sky130_vsdinv _24620_ (.A(\cpuregs[2][14] ),
    .Y(_00724_));
 sky130_vsdinv _24621_ (.A(\cpuregs[3][14] ),
    .Y(_00725_));
 sky130_vsdinv _24622_ (.A(\cpuregs[4][14] ),
    .Y(_00727_));
 sky130_vsdinv _24623_ (.A(\cpuregs[5][14] ),
    .Y(_00728_));
 sky130_vsdinv _24624_ (.A(\cpuregs[6][14] ),
    .Y(_00729_));
 sky130_vsdinv _24625_ (.A(\cpuregs[7][14] ),
    .Y(_00730_));
 sky130_vsdinv _24626_ (.A(\cpuregs[8][14] ),
    .Y(_00732_));
 sky130_vsdinv _24627_ (.A(\cpuregs[9][14] ),
    .Y(_00733_));
 sky130_vsdinv _24628_ (.A(\cpuregs[10][14] ),
    .Y(_00734_));
 sky130_vsdinv _24629_ (.A(\cpuregs[11][14] ),
    .Y(_00735_));
 sky130_vsdinv _24630_ (.A(\cpuregs[12][14] ),
    .Y(_00737_));
 sky130_vsdinv _24631_ (.A(\cpuregs[13][14] ),
    .Y(_00738_));
 sky130_vsdinv _24632_ (.A(\cpuregs[14][14] ),
    .Y(_00739_));
 sky130_vsdinv _24633_ (.A(\cpuregs[15][14] ),
    .Y(_00740_));
 sky130_vsdinv _24634_ (.A(\cpuregs[16][14] ),
    .Y(_00743_));
 sky130_vsdinv _24635_ (.A(\cpuregs[17][14] ),
    .Y(_00744_));
 sky130_vsdinv _24636_ (.A(\cpuregs[18][14] ),
    .Y(_00745_));
 sky130_vsdinv _24637_ (.A(\cpuregs[19][14] ),
    .Y(_00746_));
 sky130_vsdinv _24638_ (.A(\cpuregs[0][15] ),
    .Y(_00749_));
 sky130_vsdinv _24639_ (.A(\cpuregs[1][15] ),
    .Y(_00750_));
 sky130_vsdinv _24640_ (.A(\cpuregs[2][15] ),
    .Y(_00751_));
 sky130_vsdinv _24641_ (.A(\cpuregs[3][15] ),
    .Y(_00752_));
 sky130_vsdinv _24642_ (.A(\cpuregs[4][15] ),
    .Y(_00754_));
 sky130_vsdinv _24643_ (.A(\cpuregs[5][15] ),
    .Y(_00755_));
 sky130_vsdinv _24644_ (.A(\cpuregs[6][15] ),
    .Y(_00756_));
 sky130_vsdinv _24645_ (.A(\cpuregs[7][15] ),
    .Y(_00757_));
 sky130_vsdinv _24646_ (.A(\cpuregs[8][15] ),
    .Y(_00759_));
 sky130_vsdinv _24647_ (.A(\cpuregs[9][15] ),
    .Y(_00760_));
 sky130_vsdinv _24648_ (.A(\cpuregs[10][15] ),
    .Y(_00761_));
 sky130_vsdinv _24649_ (.A(\cpuregs[11][15] ),
    .Y(_00762_));
 sky130_vsdinv _24650_ (.A(\cpuregs[12][15] ),
    .Y(_00764_));
 sky130_vsdinv _24651_ (.A(\cpuregs[13][15] ),
    .Y(_00765_));
 sky130_vsdinv _24652_ (.A(\cpuregs[14][15] ),
    .Y(_00766_));
 sky130_vsdinv _24653_ (.A(\cpuregs[15][15] ),
    .Y(_00767_));
 sky130_vsdinv _24654_ (.A(\cpuregs[16][15] ),
    .Y(_00770_));
 sky130_vsdinv _24655_ (.A(\cpuregs[17][15] ),
    .Y(_00771_));
 sky130_vsdinv _24656_ (.A(\cpuregs[18][15] ),
    .Y(_00772_));
 sky130_vsdinv _24657_ (.A(\cpuregs[19][15] ),
    .Y(_00773_));
 sky130_vsdinv _24658_ (.A(\cpuregs[0][16] ),
    .Y(_00776_));
 sky130_vsdinv _24659_ (.A(\cpuregs[1][16] ),
    .Y(_00777_));
 sky130_vsdinv _24660_ (.A(\cpuregs[2][16] ),
    .Y(_00778_));
 sky130_vsdinv _24661_ (.A(\cpuregs[3][16] ),
    .Y(_00779_));
 sky130_vsdinv _24662_ (.A(\cpuregs[4][16] ),
    .Y(_00781_));
 sky130_vsdinv _24663_ (.A(\cpuregs[5][16] ),
    .Y(_00782_));
 sky130_vsdinv _24664_ (.A(\cpuregs[6][16] ),
    .Y(_00783_));
 sky130_vsdinv _24665_ (.A(\cpuregs[7][16] ),
    .Y(_00784_));
 sky130_vsdinv _24666_ (.A(\cpuregs[8][16] ),
    .Y(_00786_));
 sky130_vsdinv _24667_ (.A(\cpuregs[9][16] ),
    .Y(_00787_));
 sky130_vsdinv _24668_ (.A(\cpuregs[10][16] ),
    .Y(_00788_));
 sky130_vsdinv _24669_ (.A(\cpuregs[11][16] ),
    .Y(_00789_));
 sky130_vsdinv _24670_ (.A(\cpuregs[12][16] ),
    .Y(_00791_));
 sky130_vsdinv _24671_ (.A(\cpuregs[13][16] ),
    .Y(_00792_));
 sky130_vsdinv _24672_ (.A(\cpuregs[14][16] ),
    .Y(_00793_));
 sky130_vsdinv _24673_ (.A(\cpuregs[15][16] ),
    .Y(_00794_));
 sky130_vsdinv _24674_ (.A(\cpuregs[16][16] ),
    .Y(_00797_));
 sky130_vsdinv _24675_ (.A(\cpuregs[17][16] ),
    .Y(_00798_));
 sky130_vsdinv _24676_ (.A(\cpuregs[18][16] ),
    .Y(_00799_));
 sky130_vsdinv _24677_ (.A(\cpuregs[19][16] ),
    .Y(_00800_));
 sky130_vsdinv _24678_ (.A(\cpuregs[0][17] ),
    .Y(_00803_));
 sky130_vsdinv _24679_ (.A(\cpuregs[1][17] ),
    .Y(_00804_));
 sky130_vsdinv _24680_ (.A(\cpuregs[2][17] ),
    .Y(_00805_));
 sky130_vsdinv _24681_ (.A(\cpuregs[3][17] ),
    .Y(_00806_));
 sky130_vsdinv _24682_ (.A(\cpuregs[4][17] ),
    .Y(_00808_));
 sky130_vsdinv _24683_ (.A(\cpuregs[5][17] ),
    .Y(_00809_));
 sky130_vsdinv _24684_ (.A(\cpuregs[6][17] ),
    .Y(_00810_));
 sky130_vsdinv _24685_ (.A(\cpuregs[7][17] ),
    .Y(_00811_));
 sky130_vsdinv _24686_ (.A(\cpuregs[8][17] ),
    .Y(_00813_));
 sky130_vsdinv _24687_ (.A(\cpuregs[9][17] ),
    .Y(_00814_));
 sky130_vsdinv _24688_ (.A(\cpuregs[10][17] ),
    .Y(_00815_));
 sky130_vsdinv _24689_ (.A(\cpuregs[11][17] ),
    .Y(_00816_));
 sky130_vsdinv _24690_ (.A(\cpuregs[12][17] ),
    .Y(_00818_));
 sky130_vsdinv _24691_ (.A(\cpuregs[13][17] ),
    .Y(_00819_));
 sky130_vsdinv _24692_ (.A(\cpuregs[14][17] ),
    .Y(_00820_));
 sky130_vsdinv _24693_ (.A(\cpuregs[15][17] ),
    .Y(_00821_));
 sky130_vsdinv _24694_ (.A(\cpuregs[16][17] ),
    .Y(_00824_));
 sky130_vsdinv _24695_ (.A(\cpuregs[17][17] ),
    .Y(_00825_));
 sky130_vsdinv _24696_ (.A(\cpuregs[18][17] ),
    .Y(_00826_));
 sky130_vsdinv _24697_ (.A(\cpuregs[19][17] ),
    .Y(_00827_));
 sky130_vsdinv _24698_ (.A(\cpuregs[0][18] ),
    .Y(_00830_));
 sky130_vsdinv _24699_ (.A(\cpuregs[1][18] ),
    .Y(_00831_));
 sky130_vsdinv _24700_ (.A(\cpuregs[2][18] ),
    .Y(_00832_));
 sky130_vsdinv _24701_ (.A(\cpuregs[3][18] ),
    .Y(_00833_));
 sky130_vsdinv _24702_ (.A(\cpuregs[4][18] ),
    .Y(_00835_));
 sky130_vsdinv _24703_ (.A(\cpuregs[5][18] ),
    .Y(_00836_));
 sky130_vsdinv _24704_ (.A(\cpuregs[6][18] ),
    .Y(_00837_));
 sky130_vsdinv _24705_ (.A(\cpuregs[7][18] ),
    .Y(_00838_));
 sky130_vsdinv _24706_ (.A(\cpuregs[8][18] ),
    .Y(_00840_));
 sky130_vsdinv _24707_ (.A(\cpuregs[9][18] ),
    .Y(_00841_));
 sky130_vsdinv _24708_ (.A(\cpuregs[10][18] ),
    .Y(_00842_));
 sky130_vsdinv _24709_ (.A(\cpuregs[11][18] ),
    .Y(_00843_));
 sky130_vsdinv _24710_ (.A(\cpuregs[12][18] ),
    .Y(_00845_));
 sky130_vsdinv _24711_ (.A(\cpuregs[13][18] ),
    .Y(_00846_));
 sky130_vsdinv _24712_ (.A(\cpuregs[14][18] ),
    .Y(_00847_));
 sky130_vsdinv _24713_ (.A(\cpuregs[15][18] ),
    .Y(_00848_));
 sky130_vsdinv _24714_ (.A(\cpuregs[16][18] ),
    .Y(_00851_));
 sky130_vsdinv _24715_ (.A(\cpuregs[17][18] ),
    .Y(_00852_));
 sky130_vsdinv _24716_ (.A(\cpuregs[18][18] ),
    .Y(_00853_));
 sky130_vsdinv _24717_ (.A(\cpuregs[19][18] ),
    .Y(_00854_));
 sky130_vsdinv _24718_ (.A(\cpuregs[0][19] ),
    .Y(_00857_));
 sky130_vsdinv _24719_ (.A(\cpuregs[1][19] ),
    .Y(_00858_));
 sky130_vsdinv _24720_ (.A(\cpuregs[2][19] ),
    .Y(_00859_));
 sky130_vsdinv _24721_ (.A(\cpuregs[3][19] ),
    .Y(_00860_));
 sky130_vsdinv _24722_ (.A(\cpuregs[4][19] ),
    .Y(_00862_));
 sky130_vsdinv _24723_ (.A(\cpuregs[5][19] ),
    .Y(_00863_));
 sky130_vsdinv _24724_ (.A(\cpuregs[6][19] ),
    .Y(_00864_));
 sky130_vsdinv _24725_ (.A(\cpuregs[7][19] ),
    .Y(_00865_));
 sky130_vsdinv _24726_ (.A(\cpuregs[8][19] ),
    .Y(_00867_));
 sky130_vsdinv _24727_ (.A(\cpuregs[9][19] ),
    .Y(_00868_));
 sky130_vsdinv _24728_ (.A(\cpuregs[10][19] ),
    .Y(_00869_));
 sky130_vsdinv _24729_ (.A(\cpuregs[11][19] ),
    .Y(_00870_));
 sky130_vsdinv _24730_ (.A(\cpuregs[12][19] ),
    .Y(_00872_));
 sky130_vsdinv _24731_ (.A(\cpuregs[13][19] ),
    .Y(_00873_));
 sky130_vsdinv _24732_ (.A(\cpuregs[14][19] ),
    .Y(_00874_));
 sky130_vsdinv _24733_ (.A(\cpuregs[15][19] ),
    .Y(_00875_));
 sky130_vsdinv _24734_ (.A(\cpuregs[16][19] ),
    .Y(_00878_));
 sky130_vsdinv _24735_ (.A(\cpuregs[17][19] ),
    .Y(_00879_));
 sky130_vsdinv _24736_ (.A(\cpuregs[18][19] ),
    .Y(_00880_));
 sky130_vsdinv _24737_ (.A(\cpuregs[19][19] ),
    .Y(_00881_));
 sky130_vsdinv _24738_ (.A(\cpuregs[0][20] ),
    .Y(_00884_));
 sky130_vsdinv _24739_ (.A(\cpuregs[1][20] ),
    .Y(_00885_));
 sky130_vsdinv _24740_ (.A(\cpuregs[2][20] ),
    .Y(_00886_));
 sky130_vsdinv _24741_ (.A(\cpuregs[3][20] ),
    .Y(_00887_));
 sky130_vsdinv _24742_ (.A(\cpuregs[4][20] ),
    .Y(_00889_));
 sky130_vsdinv _24743_ (.A(\cpuregs[5][20] ),
    .Y(_00890_));
 sky130_vsdinv _24744_ (.A(\cpuregs[6][20] ),
    .Y(_00891_));
 sky130_vsdinv _24745_ (.A(\cpuregs[7][20] ),
    .Y(_00892_));
 sky130_vsdinv _24746_ (.A(\cpuregs[8][20] ),
    .Y(_00894_));
 sky130_vsdinv _24747_ (.A(\cpuregs[9][20] ),
    .Y(_00895_));
 sky130_vsdinv _24748_ (.A(\cpuregs[10][20] ),
    .Y(_00896_));
 sky130_vsdinv _24749_ (.A(\cpuregs[11][20] ),
    .Y(_00897_));
 sky130_vsdinv _24750_ (.A(\cpuregs[12][20] ),
    .Y(_00899_));
 sky130_vsdinv _24751_ (.A(\cpuregs[13][20] ),
    .Y(_00900_));
 sky130_vsdinv _24752_ (.A(\cpuregs[14][20] ),
    .Y(_00901_));
 sky130_vsdinv _24753_ (.A(\cpuregs[15][20] ),
    .Y(_00902_));
 sky130_vsdinv _24754_ (.A(\cpuregs[16][20] ),
    .Y(_00905_));
 sky130_vsdinv _24755_ (.A(\cpuregs[17][20] ),
    .Y(_00906_));
 sky130_vsdinv _24756_ (.A(\cpuregs[18][20] ),
    .Y(_00907_));
 sky130_vsdinv _24757_ (.A(\cpuregs[19][20] ),
    .Y(_00908_));
 sky130_vsdinv _24758_ (.A(\cpuregs[0][21] ),
    .Y(_00911_));
 sky130_vsdinv _24759_ (.A(\cpuregs[1][21] ),
    .Y(_00912_));
 sky130_vsdinv _24760_ (.A(\cpuregs[2][21] ),
    .Y(_00913_));
 sky130_vsdinv _24761_ (.A(\cpuregs[3][21] ),
    .Y(_00914_));
 sky130_vsdinv _24762_ (.A(\cpuregs[4][21] ),
    .Y(_00916_));
 sky130_vsdinv _24763_ (.A(\cpuregs[5][21] ),
    .Y(_00917_));
 sky130_vsdinv _24764_ (.A(\cpuregs[6][21] ),
    .Y(_00918_));
 sky130_vsdinv _24765_ (.A(\cpuregs[7][21] ),
    .Y(_00919_));
 sky130_fd_sc_hd__buf_1 _24766_ (.A(_19121_),
    .X(_19775_));
 sky130_fd_sc_hd__nor2_2 _24767_ (.A(_19117_),
    .B(_19775_),
    .Y(_00304_));
 sky130_vsdinv _24768_ (.A(\cpuregs[8][21] ),
    .Y(_00921_));
 sky130_vsdinv _24769_ (.A(\cpuregs[9][21] ),
    .Y(_00922_));
 sky130_vsdinv _24770_ (.A(\cpuregs[10][21] ),
    .Y(_00923_));
 sky130_vsdinv _24771_ (.A(\cpuregs[11][21] ),
    .Y(_00924_));
 sky130_vsdinv _24772_ (.A(\cpuregs[12][21] ),
    .Y(_00926_));
 sky130_vsdinv _24773_ (.A(\cpuregs[13][21] ),
    .Y(_00927_));
 sky130_vsdinv _24774_ (.A(\cpuregs[14][21] ),
    .Y(_00928_));
 sky130_vsdinv _24775_ (.A(\cpuregs[15][21] ),
    .Y(_00929_));
 sky130_vsdinv _24776_ (.A(\cpuregs[16][21] ),
    .Y(_00932_));
 sky130_vsdinv _24777_ (.A(\cpuregs[17][21] ),
    .Y(_00933_));
 sky130_vsdinv _24778_ (.A(\cpuregs[18][21] ),
    .Y(_00934_));
 sky130_vsdinv _24779_ (.A(\cpuregs[19][21] ),
    .Y(_00935_));
 sky130_vsdinv _24780_ (.A(\cpuregs[0][22] ),
    .Y(_00938_));
 sky130_vsdinv _24781_ (.A(\cpuregs[1][22] ),
    .Y(_00939_));
 sky130_vsdinv _24782_ (.A(\cpuregs[2][22] ),
    .Y(_00940_));
 sky130_vsdinv _24783_ (.A(\cpuregs[3][22] ),
    .Y(_00941_));
 sky130_vsdinv _24784_ (.A(\cpuregs[4][22] ),
    .Y(_00943_));
 sky130_vsdinv _24785_ (.A(\cpuregs[5][22] ),
    .Y(_00944_));
 sky130_vsdinv _24786_ (.A(\cpuregs[6][22] ),
    .Y(_00945_));
 sky130_vsdinv _24787_ (.A(\cpuregs[7][22] ),
    .Y(_00946_));
 sky130_fd_sc_hd__and4_2 _24788_ (.A(_16849_),
    .B(_16837_),
    .C(instr_lw),
    .D(_19759_),
    .X(_19776_));
 sky130_fd_sc_hd__a31o_2 _24789_ (.A1(instr_sw),
    .A2(_19664_),
    .A3(_17383_),
    .B1(_19776_),
    .X(_19777_));
 sky130_fd_sc_hd__a221o_2 _24790_ (.A1(_19646_),
    .A2(_19777_),
    .B1(_19762_),
    .B2(\mem_wordsize[0] ),
    .C1(_18291_),
    .X(_00045_));
 sky130_vsdinv _24791_ (.A(\cpuregs[8][22] ),
    .Y(_00948_));
 sky130_vsdinv _24792_ (.A(\cpuregs[9][22] ),
    .Y(_00949_));
 sky130_vsdinv _24793_ (.A(\cpuregs[10][22] ),
    .Y(_00950_));
 sky130_vsdinv _24794_ (.A(\cpuregs[11][22] ),
    .Y(_00951_));
 sky130_vsdinv _24795_ (.A(\cpuregs[12][22] ),
    .Y(_00953_));
 sky130_vsdinv _24796_ (.A(\cpuregs[13][22] ),
    .Y(_00954_));
 sky130_vsdinv _24797_ (.A(\cpuregs[14][22] ),
    .Y(_00955_));
 sky130_vsdinv _24798_ (.A(\cpuregs[15][22] ),
    .Y(_00956_));
 sky130_vsdinv _24799_ (.A(\cpuregs[16][22] ),
    .Y(_00959_));
 sky130_vsdinv _24800_ (.A(\cpuregs[17][22] ),
    .Y(_00960_));
 sky130_vsdinv _24801_ (.A(\cpuregs[18][22] ),
    .Y(_00961_));
 sky130_vsdinv _24802_ (.A(\cpuregs[19][22] ),
    .Y(_00962_));
 sky130_vsdinv _24803_ (.A(\cpuregs[0][23] ),
    .Y(_00965_));
 sky130_vsdinv _24804_ (.A(\cpuregs[1][23] ),
    .Y(_00966_));
 sky130_vsdinv _24805_ (.A(\cpuregs[2][23] ),
    .Y(_00967_));
 sky130_vsdinv _24806_ (.A(\cpuregs[3][23] ),
    .Y(_00968_));
 sky130_vsdinv _24807_ (.A(\cpuregs[4][23] ),
    .Y(_00970_));
 sky130_vsdinv _24808_ (.A(\cpuregs[5][23] ),
    .Y(_00971_));
 sky130_vsdinv _24809_ (.A(\cpuregs[6][23] ),
    .Y(_00972_));
 sky130_vsdinv _24810_ (.A(\cpuregs[7][23] ),
    .Y(_00973_));
 sky130_vsdinv _24811_ (.A(\cpuregs[8][23] ),
    .Y(_00975_));
 sky130_vsdinv _24812_ (.A(\cpuregs[9][23] ),
    .Y(_00976_));
 sky130_vsdinv _24813_ (.A(\cpuregs[10][23] ),
    .Y(_00977_));
 sky130_vsdinv _24814_ (.A(\cpuregs[11][23] ),
    .Y(_00978_));
 sky130_vsdinv _24815_ (.A(\cpuregs[12][23] ),
    .Y(_00980_));
 sky130_vsdinv _24816_ (.A(\cpuregs[13][23] ),
    .Y(_00981_));
 sky130_vsdinv _24817_ (.A(\cpuregs[14][23] ),
    .Y(_00982_));
 sky130_vsdinv _24818_ (.A(\cpuregs[15][23] ),
    .Y(_00983_));
 sky130_vsdinv _24819_ (.A(\cpuregs[16][23] ),
    .Y(_00986_));
 sky130_vsdinv _24820_ (.A(\cpuregs[17][23] ),
    .Y(_00987_));
 sky130_vsdinv _24821_ (.A(\cpuregs[18][23] ),
    .Y(_00988_));
 sky130_vsdinv _24822_ (.A(\cpuregs[19][23] ),
    .Y(_00989_));
 sky130_vsdinv _24823_ (.A(\cpuregs[0][24] ),
    .Y(_00992_));
 sky130_vsdinv _24824_ (.A(\cpuregs[1][24] ),
    .Y(_00993_));
 sky130_vsdinv _24825_ (.A(\cpuregs[2][24] ),
    .Y(_00994_));
 sky130_vsdinv _24826_ (.A(\cpuregs[3][24] ),
    .Y(_00995_));
 sky130_vsdinv _24827_ (.A(\cpuregs[4][24] ),
    .Y(_00997_));
 sky130_vsdinv _24828_ (.A(\cpuregs[5][24] ),
    .Y(_00998_));
 sky130_vsdinv _24829_ (.A(\cpuregs[6][24] ),
    .Y(_00999_));
 sky130_vsdinv _24830_ (.A(\cpuregs[7][24] ),
    .Y(_01000_));
 sky130_vsdinv _24831_ (.A(\cpuregs[8][24] ),
    .Y(_01002_));
 sky130_vsdinv _24832_ (.A(\cpuregs[9][24] ),
    .Y(_01003_));
 sky130_vsdinv _24833_ (.A(\cpuregs[10][24] ),
    .Y(_01004_));
 sky130_vsdinv _24834_ (.A(\cpuregs[11][24] ),
    .Y(_01005_));
 sky130_vsdinv _24835_ (.A(\cpuregs[12][24] ),
    .Y(_01007_));
 sky130_vsdinv _24836_ (.A(\cpuregs[13][24] ),
    .Y(_01008_));
 sky130_vsdinv _24837_ (.A(\cpuregs[14][24] ),
    .Y(_01009_));
 sky130_vsdinv _24838_ (.A(\cpuregs[15][24] ),
    .Y(_01010_));
 sky130_vsdinv _24839_ (.A(\cpuregs[16][24] ),
    .Y(_01013_));
 sky130_vsdinv _24840_ (.A(\cpuregs[17][24] ),
    .Y(_01014_));
 sky130_vsdinv _24841_ (.A(\cpuregs[18][24] ),
    .Y(_01015_));
 sky130_vsdinv _24842_ (.A(\cpuregs[19][24] ),
    .Y(_01016_));
 sky130_vsdinv _24843_ (.A(\cpuregs[0][25] ),
    .Y(_01019_));
 sky130_vsdinv _24844_ (.A(\cpuregs[1][25] ),
    .Y(_01020_));
 sky130_vsdinv _24845_ (.A(\cpuregs[2][25] ),
    .Y(_01021_));
 sky130_vsdinv _24846_ (.A(\cpuregs[3][25] ),
    .Y(_01022_));
 sky130_vsdinv _24847_ (.A(\cpuregs[4][25] ),
    .Y(_01024_));
 sky130_vsdinv _24848_ (.A(\cpuregs[5][25] ),
    .Y(_01025_));
 sky130_vsdinv _24849_ (.A(\cpuregs[6][25] ),
    .Y(_01026_));
 sky130_vsdinv _24850_ (.A(\cpuregs[7][25] ),
    .Y(_01027_));
 sky130_fd_sc_hd__nor2b_2 _24851_ (.A(_16835_),
    .B_N(_16844_),
    .Y(_00289_));
 sky130_fd_sc_hd__nand2_2 _24852_ (.A(_16856_),
    .B(_00289_),
    .Y(_00298_));
 sky130_vsdinv _24853_ (.A(\cpuregs[8][25] ),
    .Y(_01029_));
 sky130_vsdinv _24854_ (.A(\cpuregs[9][25] ),
    .Y(_01030_));
 sky130_vsdinv _24855_ (.A(\cpuregs[10][25] ),
    .Y(_01031_));
 sky130_vsdinv _24856_ (.A(\cpuregs[11][25] ),
    .Y(_01032_));
 sky130_vsdinv _24857_ (.A(\cpuregs[12][25] ),
    .Y(_01034_));
 sky130_vsdinv _24858_ (.A(\cpuregs[13][25] ),
    .Y(_01035_));
 sky130_vsdinv _24859_ (.A(\cpuregs[14][25] ),
    .Y(_01036_));
 sky130_vsdinv _24860_ (.A(\cpuregs[15][25] ),
    .Y(_01037_));
 sky130_vsdinv _24861_ (.A(\cpuregs[16][25] ),
    .Y(_01040_));
 sky130_vsdinv _24862_ (.A(\cpuregs[17][25] ),
    .Y(_01041_));
 sky130_vsdinv _24863_ (.A(\cpuregs[18][25] ),
    .Y(_01042_));
 sky130_vsdinv _24864_ (.A(\cpuregs[19][25] ),
    .Y(_01043_));
 sky130_vsdinv _24865_ (.A(\cpuregs[0][26] ),
    .Y(_01046_));
 sky130_vsdinv _24866_ (.A(\cpuregs[1][26] ),
    .Y(_01047_));
 sky130_vsdinv _24867_ (.A(\cpuregs[2][26] ),
    .Y(_01048_));
 sky130_vsdinv _24868_ (.A(\cpuregs[3][26] ),
    .Y(_01049_));
 sky130_vsdinv _24869_ (.A(\cpuregs[4][26] ),
    .Y(_01051_));
 sky130_vsdinv _24870_ (.A(\cpuregs[5][26] ),
    .Y(_01052_));
 sky130_vsdinv _24871_ (.A(\cpuregs[6][26] ),
    .Y(_01053_));
 sky130_vsdinv _24872_ (.A(\cpuregs[7][26] ),
    .Y(_01054_));
 sky130_vsdinv _24873_ (.A(\cpuregs[8][26] ),
    .Y(_01056_));
 sky130_vsdinv _24874_ (.A(\cpuregs[9][26] ),
    .Y(_01057_));
 sky130_vsdinv _24875_ (.A(\cpuregs[10][26] ),
    .Y(_01058_));
 sky130_vsdinv _24876_ (.A(\cpuregs[11][26] ),
    .Y(_01059_));
 sky130_vsdinv _24877_ (.A(\cpuregs[12][26] ),
    .Y(_01061_));
 sky130_vsdinv _24878_ (.A(\cpuregs[13][26] ),
    .Y(_01062_));
 sky130_vsdinv _24879_ (.A(\cpuregs[14][26] ),
    .Y(_01063_));
 sky130_vsdinv _24880_ (.A(\cpuregs[15][26] ),
    .Y(_01064_));
 sky130_vsdinv _24881_ (.A(\cpuregs[16][26] ),
    .Y(_01067_));
 sky130_vsdinv _24882_ (.A(\cpuregs[17][26] ),
    .Y(_01068_));
 sky130_vsdinv _24883_ (.A(\cpuregs[18][26] ),
    .Y(_01069_));
 sky130_vsdinv _24884_ (.A(\cpuregs[19][26] ),
    .Y(_01070_));
 sky130_fd_sc_hd__buf_1 _24885_ (.A(_19759_),
    .X(_04073_));
 sky130_fd_sc_hd__o211ai_2 _24886_ (.A1(instr_lbu),
    .A2(instr_lb),
    .B1(_19763_),
    .C1(_04073_),
    .Y(_04074_));
 sky130_fd_sc_hd__o31ai_2 _24887_ (.A1(_17218_),
    .A2(_19013_),
    .A3(_18030_),
    .B1(_04074_),
    .Y(_04075_));
 sky130_fd_sc_hd__buf_1 _24888_ (.A(\mem_wordsize[1] ),
    .X(_04076_));
 sky130_fd_sc_hd__buf_1 _24889_ (.A(_04076_),
    .X(_04077_));
 sky130_fd_sc_hd__buf_1 _24890_ (.A(_04077_),
    .X(_04078_));
 sky130_fd_sc_hd__a22o_2 _24891_ (.A1(_16810_),
    .A2(_04075_),
    .B1(_19762_),
    .B2(_04078_),
    .X(_00046_));
 sky130_vsdinv _24892_ (.A(\cpuregs[0][27] ),
    .Y(_01073_));
 sky130_vsdinv _24893_ (.A(\cpuregs[1][27] ),
    .Y(_01074_));
 sky130_vsdinv _24894_ (.A(\cpuregs[2][27] ),
    .Y(_01075_));
 sky130_vsdinv _24895_ (.A(\cpuregs[3][27] ),
    .Y(_01076_));
 sky130_vsdinv _24896_ (.A(\cpuregs[4][27] ),
    .Y(_01078_));
 sky130_vsdinv _24897_ (.A(\cpuregs[5][27] ),
    .Y(_01079_));
 sky130_vsdinv _24898_ (.A(\cpuregs[6][27] ),
    .Y(_01080_));
 sky130_vsdinv _24899_ (.A(\cpuregs[7][27] ),
    .Y(_01081_));
 sky130_vsdinv _24900_ (.A(\cpuregs[8][27] ),
    .Y(_01083_));
 sky130_vsdinv _24901_ (.A(\cpuregs[9][27] ),
    .Y(_01084_));
 sky130_vsdinv _24902_ (.A(\cpuregs[10][27] ),
    .Y(_01085_));
 sky130_vsdinv _24903_ (.A(\cpuregs[11][27] ),
    .Y(_01086_));
 sky130_vsdinv _24904_ (.A(\cpuregs[12][27] ),
    .Y(_01088_));
 sky130_vsdinv _24905_ (.A(\cpuregs[13][27] ),
    .Y(_01089_));
 sky130_vsdinv _24906_ (.A(\cpuregs[14][27] ),
    .Y(_01090_));
 sky130_vsdinv _24907_ (.A(\cpuregs[15][27] ),
    .Y(_01091_));
 sky130_vsdinv _24908_ (.A(\cpuregs[16][27] ),
    .Y(_01094_));
 sky130_vsdinv _24909_ (.A(\cpuregs[17][27] ),
    .Y(_01095_));
 sky130_vsdinv _24910_ (.A(\cpuregs[18][27] ),
    .Y(_01096_));
 sky130_vsdinv _24911_ (.A(\cpuregs[19][27] ),
    .Y(_01097_));
 sky130_vsdinv _24912_ (.A(\cpuregs[0][28] ),
    .Y(_01100_));
 sky130_vsdinv _24913_ (.A(\cpuregs[1][28] ),
    .Y(_01101_));
 sky130_vsdinv _24914_ (.A(\cpuregs[2][28] ),
    .Y(_01102_));
 sky130_vsdinv _24915_ (.A(\cpuregs[3][28] ),
    .Y(_01103_));
 sky130_vsdinv _24916_ (.A(\cpuregs[4][28] ),
    .Y(_01105_));
 sky130_vsdinv _24917_ (.A(\cpuregs[5][28] ),
    .Y(_01106_));
 sky130_vsdinv _24918_ (.A(\cpuregs[6][28] ),
    .Y(_01107_));
 sky130_vsdinv _24919_ (.A(\cpuregs[7][28] ),
    .Y(_01108_));
 sky130_vsdinv _24920_ (.A(\cpuregs[8][28] ),
    .Y(_01110_));
 sky130_vsdinv _24921_ (.A(\cpuregs[9][28] ),
    .Y(_01111_));
 sky130_vsdinv _24922_ (.A(\cpuregs[10][28] ),
    .Y(_01112_));
 sky130_vsdinv _24923_ (.A(\cpuregs[11][28] ),
    .Y(_01113_));
 sky130_vsdinv _24924_ (.A(\cpuregs[12][28] ),
    .Y(_01115_));
 sky130_vsdinv _24925_ (.A(\cpuregs[13][28] ),
    .Y(_01116_));
 sky130_vsdinv _24926_ (.A(\cpuregs[14][28] ),
    .Y(_01117_));
 sky130_vsdinv _24927_ (.A(\cpuregs[15][28] ),
    .Y(_01118_));
 sky130_vsdinv _24928_ (.A(\cpuregs[16][28] ),
    .Y(_01121_));
 sky130_vsdinv _24929_ (.A(\cpuregs[17][28] ),
    .Y(_01122_));
 sky130_vsdinv _24930_ (.A(\cpuregs[18][28] ),
    .Y(_01123_));
 sky130_vsdinv _24931_ (.A(\cpuregs[19][28] ),
    .Y(_01124_));
 sky130_vsdinv _24932_ (.A(\cpuregs[0][29] ),
    .Y(_01127_));
 sky130_vsdinv _24933_ (.A(\cpuregs[1][29] ),
    .Y(_01128_));
 sky130_vsdinv _24934_ (.A(\cpuregs[2][29] ),
    .Y(_01129_));
 sky130_vsdinv _24935_ (.A(\cpuregs[3][29] ),
    .Y(_01130_));
 sky130_vsdinv _24936_ (.A(\cpuregs[4][29] ),
    .Y(_01132_));
 sky130_vsdinv _24937_ (.A(\cpuregs[5][29] ),
    .Y(_01133_));
 sky130_vsdinv _24938_ (.A(\cpuregs[6][29] ),
    .Y(_01134_));
 sky130_vsdinv _24939_ (.A(\cpuregs[7][29] ),
    .Y(_01135_));
 sky130_vsdinv _24940_ (.A(\cpuregs[8][29] ),
    .Y(_01137_));
 sky130_vsdinv _24941_ (.A(\cpuregs[9][29] ),
    .Y(_01138_));
 sky130_vsdinv _24942_ (.A(\cpuregs[10][29] ),
    .Y(_01139_));
 sky130_vsdinv _24943_ (.A(\cpuregs[11][29] ),
    .Y(_01140_));
 sky130_vsdinv _24944_ (.A(\cpuregs[12][29] ),
    .Y(_01142_));
 sky130_vsdinv _24945_ (.A(\cpuregs[13][29] ),
    .Y(_01143_));
 sky130_fd_sc_hd__buf_1 _24946_ (.A(latched_branch),
    .X(_04079_));
 sky130_fd_sc_hd__buf_1 _24947_ (.A(_04079_),
    .X(_04080_));
 sky130_fd_sc_hd__and2_2 _24948_ (.A(_04080_),
    .B(_00294_),
    .X(_00295_));
 sky130_vsdinv _24949_ (.A(\cpuregs[14][29] ),
    .Y(_01144_));
 sky130_vsdinv _24950_ (.A(\cpuregs[15][29] ),
    .Y(_01145_));
 sky130_vsdinv _24951_ (.A(\cpuregs[16][29] ),
    .Y(_01148_));
 sky130_vsdinv _24952_ (.A(\cpuregs[17][29] ),
    .Y(_01149_));
 sky130_vsdinv _24953_ (.A(\cpuregs[18][29] ),
    .Y(_01150_));
 sky130_vsdinv _24954_ (.A(\cpuregs[19][29] ),
    .Y(_01151_));
 sky130_vsdinv _24955_ (.A(\cpuregs[0][30] ),
    .Y(_01154_));
 sky130_vsdinv _24956_ (.A(\cpuregs[1][30] ),
    .Y(_01155_));
 sky130_vsdinv _24957_ (.A(\cpuregs[2][30] ),
    .Y(_01156_));
 sky130_vsdinv _24958_ (.A(\cpuregs[3][30] ),
    .Y(_01157_));
 sky130_vsdinv _24959_ (.A(\cpuregs[4][30] ),
    .Y(_01159_));
 sky130_vsdinv _24960_ (.A(\cpuregs[5][30] ),
    .Y(_01160_));
 sky130_vsdinv _24961_ (.A(\cpuregs[6][30] ),
    .Y(_01161_));
 sky130_vsdinv _24962_ (.A(\cpuregs[7][30] ),
    .Y(_01162_));
 sky130_vsdinv _24963_ (.A(\cpuregs[8][30] ),
    .Y(_01164_));
 sky130_vsdinv _24964_ (.A(\cpuregs[9][30] ),
    .Y(_01165_));
 sky130_vsdinv _24965_ (.A(\cpuregs[10][30] ),
    .Y(_01166_));
 sky130_vsdinv _24966_ (.A(\cpuregs[11][30] ),
    .Y(_01167_));
 sky130_vsdinv _24967_ (.A(\cpuregs[12][30] ),
    .Y(_01169_));
 sky130_vsdinv _24968_ (.A(\cpuregs[13][30] ),
    .Y(_01170_));
 sky130_vsdinv _24969_ (.A(\cpuregs[14][30] ),
    .Y(_01171_));
 sky130_vsdinv _24970_ (.A(\cpuregs[15][30] ),
    .Y(_01172_));
 sky130_vsdinv _24971_ (.A(\cpuregs[16][30] ),
    .Y(_01175_));
 sky130_vsdinv _24972_ (.A(\cpuregs[17][30] ),
    .Y(_01176_));
 sky130_vsdinv _24973_ (.A(\cpuregs[18][30] ),
    .Y(_01177_));
 sky130_vsdinv _24974_ (.A(\cpuregs[19][30] ),
    .Y(_01178_));
 sky130_vsdinv _24975_ (.A(\cpuregs[0][31] ),
    .Y(_01181_));
 sky130_vsdinv _24976_ (.A(\cpuregs[1][31] ),
    .Y(_01182_));
 sky130_vsdinv _24977_ (.A(\cpuregs[2][31] ),
    .Y(_01183_));
 sky130_vsdinv _24978_ (.A(\cpuregs[3][31] ),
    .Y(_01184_));
 sky130_vsdinv _24979_ (.A(\cpuregs[4][31] ),
    .Y(_01186_));
 sky130_vsdinv _24980_ (.A(\cpuregs[5][31] ),
    .Y(_01187_));
 sky130_vsdinv _24981_ (.A(\cpuregs[6][31] ),
    .Y(_01188_));
 sky130_vsdinv _24982_ (.A(\cpuregs[7][31] ),
    .Y(_01189_));
 sky130_vsdinv _24983_ (.A(\cpuregs[8][31] ),
    .Y(_01191_));
 sky130_vsdinv _24984_ (.A(\cpuregs[9][31] ),
    .Y(_01192_));
 sky130_vsdinv _24985_ (.A(\cpuregs[10][31] ),
    .Y(_01193_));
 sky130_vsdinv _24986_ (.A(\cpuregs[11][31] ),
    .Y(_01194_));
 sky130_vsdinv _24987_ (.A(\cpuregs[12][31] ),
    .Y(_01196_));
 sky130_vsdinv _24988_ (.A(\cpuregs[13][31] ),
    .Y(_01197_));
 sky130_vsdinv _24989_ (.A(\cpuregs[14][31] ),
    .Y(_01198_));
 sky130_vsdinv _24990_ (.A(\cpuregs[15][31] ),
    .Y(_01199_));
 sky130_vsdinv _24991_ (.A(\cpuregs[16][31] ),
    .Y(_01202_));
 sky130_vsdinv _24992_ (.A(\cpuregs[17][31] ),
    .Y(_01203_));
 sky130_vsdinv _24993_ (.A(\cpuregs[18][31] ),
    .Y(_01204_));
 sky130_vsdinv _24994_ (.A(\cpuregs[19][31] ),
    .Y(_01205_));
 sky130_fd_sc_hd__nor2_2 _24995_ (.A(\timer[25] ),
    .B(\timer[26] ),
    .Y(_04081_));
 sky130_vsdinv _24996_ (.A(\timer[24] ),
    .Y(_04082_));
 sky130_fd_sc_hd__nand3b_2 _24997_ (.A_N(\timer[27] ),
    .B(_04081_),
    .C(_04082_),
    .Y(_04083_));
 sky130_fd_sc_hd__nor2_2 _24998_ (.A(\timer[17] ),
    .B(\timer[18] ),
    .Y(_04084_));
 sky130_vsdinv _24999_ (.A(\timer[16] ),
    .Y(_04085_));
 sky130_fd_sc_hd__nand3b_2 _25000_ (.A_N(\timer[19] ),
    .B(_04084_),
    .C(_04085_),
    .Y(_04086_));
 sky130_fd_sc_hd__or2_2 _25001_ (.A(\timer[9] ),
    .B(\timer[10] ),
    .X(_04087_));
 sky130_fd_sc_hd__nor3_2 _25002_ (.A(\timer[1] ),
    .B(\timer[0] ),
    .C(\timer[2] ),
    .Y(_04088_));
 sky130_vsdinv _25003_ (.A(\timer[3] ),
    .Y(_04089_));
 sky130_fd_sc_hd__nor2_2 _25004_ (.A(\timer[5] ),
    .B(\timer[4] ),
    .Y(_04090_));
 sky130_fd_sc_hd__nand3_2 _25005_ (.A(_04088_),
    .B(_04089_),
    .C(_04090_),
    .Y(_04091_));
 sky130_fd_sc_hd__or4_2 _25006_ (.A(\timer[7] ),
    .B(\timer[6] ),
    .C(\timer[8] ),
    .D(_04091_),
    .X(_04092_));
 sky130_fd_sc_hd__nor3_2 _25007_ (.A(\timer[11] ),
    .B(_04087_),
    .C(_04092_),
    .Y(_04093_));
 sky130_fd_sc_hd__nor2_2 _25008_ (.A(\timer[13] ),
    .B(\timer[12] ),
    .Y(_04094_));
 sky130_fd_sc_hd__nand3b_2 _25009_ (.A_N(\timer[14] ),
    .B(_04093_),
    .C(_04094_),
    .Y(_04095_));
 sky130_fd_sc_hd__nor3_2 _25010_ (.A(\timer[15] ),
    .B(_04086_),
    .C(_04095_),
    .Y(_04096_));
 sky130_fd_sc_hd__nor2_2 _25011_ (.A(\timer[21] ),
    .B(\timer[20] ),
    .Y(_04097_));
 sky130_fd_sc_hd__nand3b_2 _25012_ (.A_N(\timer[22] ),
    .B(_04096_),
    .C(_04097_),
    .Y(_04098_));
 sky130_fd_sc_hd__nor3_2 _25013_ (.A(\timer[23] ),
    .B(_04083_),
    .C(_04098_),
    .Y(_04099_));
 sky130_fd_sc_hd__nor2_2 _25014_ (.A(\timer[29] ),
    .B(\timer[28] ),
    .Y(_04100_));
 sky130_fd_sc_hd__nand3b_2 _25015_ (.A_N(\timer[30] ),
    .B(_04099_),
    .C(_04100_),
    .Y(_04101_));
 sky130_fd_sc_hd__nor2_2 _25016_ (.A(\timer[31] ),
    .B(_04101_),
    .Y(_01208_));
 sky130_fd_sc_hd__buf_1 _25017_ (.A(\timer[0] ),
    .X(_04102_));
 sky130_fd_sc_hd__xnor2_2 _25018_ (.A(_04102_),
    .B(_01208_),
    .Y(_01209_));
 sky130_fd_sc_hd__buf_1 _25019_ (.A(\timer[1] ),
    .X(_04103_));
 sky130_fd_sc_hd__xnor2_2 _25020_ (.A(_04103_),
    .B(_04102_),
    .Y(_01211_));
 sky130_fd_sc_hd__buf_1 _25021_ (.A(\timer[2] ),
    .X(_04104_));
 sky130_fd_sc_hd__nor2_2 _25022_ (.A(_04103_),
    .B(_04102_),
    .Y(_04105_));
 sky130_fd_sc_hd__xor2_2 _25023_ (.A(_04104_),
    .B(_04105_),
    .X(_01214_));
 sky130_fd_sc_hd__xor2_2 _25024_ (.A(\timer[3] ),
    .B(_04088_),
    .X(_01217_));
 sky130_vsdinv _25025_ (.A(\timer[4] ),
    .Y(_04106_));
 sky130_fd_sc_hd__nand3b_2 _25026_ (.A_N(_04104_),
    .B(_04105_),
    .C(_04089_),
    .Y(_04107_));
 sky130_fd_sc_hd__xor2_2 _25027_ (.A(_04106_),
    .B(_04107_),
    .X(_01220_));
 sky130_fd_sc_hd__nand3_2 _25028_ (.A(_04088_),
    .B(_04089_),
    .C(_04106_),
    .Y(_04108_));
 sky130_fd_sc_hd__buf_1 _25029_ (.A(_04091_),
    .X(_04109_));
 sky130_fd_sc_hd__a21bo_2 _25030_ (.A1(\timer[5] ),
    .A2(_04108_),
    .B1_N(_04109_),
    .X(_01223_));
 sky130_fd_sc_hd__buf_1 _25031_ (.A(\timer[6] ),
    .X(_04110_));
 sky130_fd_sc_hd__xnor2_2 _25032_ (.A(_04110_),
    .B(_04109_),
    .Y(_01226_));
 sky130_fd_sc_hd__buf_1 _25033_ (.A(\timer[7] ),
    .X(_04111_));
 sky130_fd_sc_hd__nor2_2 _25034_ (.A(_04110_),
    .B(_04109_),
    .Y(_04112_));
 sky130_fd_sc_hd__xor2_2 _25035_ (.A(_04111_),
    .B(_04112_),
    .X(_01229_));
 sky130_fd_sc_hd__buf_1 _25036_ (.A(\timer[8] ),
    .X(_04113_));
 sky130_fd_sc_hd__or3_2 _25037_ (.A(_04111_),
    .B(_04110_),
    .C(_04109_),
    .X(_04114_));
 sky130_fd_sc_hd__xnor2_2 _25038_ (.A(_04113_),
    .B(_04114_),
    .Y(_01232_));
 sky130_vsdinv _25039_ (.A(\timer[9] ),
    .Y(_04115_));
 sky130_fd_sc_hd__xor2_2 _25040_ (.A(_04115_),
    .B(_04092_),
    .X(_01235_));
 sky130_fd_sc_hd__or2b_2 _25041_ (.A(_04092_),
    .B_N(_04115_),
    .X(_04116_));
 sky130_fd_sc_hd__o2bb2ai_2 _25042_ (.A1_N(\timer[10] ),
    .A2_N(_04116_),
    .B1(_04092_),
    .B2(_04087_),
    .Y(_01238_));
 sky130_fd_sc_hd__buf_1 _25043_ (.A(\timer[11] ),
    .X(_04117_));
 sky130_fd_sc_hd__nor3_2 _25044_ (.A(_04113_),
    .B(_04087_),
    .C(_04114_),
    .Y(_04118_));
 sky130_fd_sc_hd__xor2_2 _25045_ (.A(_04117_),
    .B(_04118_),
    .X(_01241_));
 sky130_fd_sc_hd__xor2_2 _25046_ (.A(\timer[12] ),
    .B(_04093_),
    .X(_01244_));
 sky130_fd_sc_hd__or2b_2 _25047_ (.A(\timer[12] ),
    .B_N(_04093_),
    .X(_04119_));
 sky130_fd_sc_hd__and3b_2 _25048_ (.A_N(_04117_),
    .B(_04118_),
    .C(_04094_),
    .X(_04120_));
 sky130_fd_sc_hd__a21o_2 _25049_ (.A1(_04119_),
    .A2(\timer[13] ),
    .B1(_04120_),
    .X(_01247_));
 sky130_fd_sc_hd__xor2_2 _25050_ (.A(\timer[14] ),
    .B(_04120_),
    .X(_01250_));
 sky130_fd_sc_hd__buf_1 _25051_ (.A(\timer[15] ),
    .X(_04121_));
 sky130_fd_sc_hd__xnor2_2 _25052_ (.A(_04121_),
    .B(_04095_),
    .Y(_01253_));
 sky130_fd_sc_hd__nor2_2 _25053_ (.A(_04121_),
    .B(_04095_),
    .Y(_04122_));
 sky130_fd_sc_hd__buf_1 _25054_ (.A(_04122_),
    .X(_04123_));
 sky130_fd_sc_hd__xor2_2 _25055_ (.A(\timer[16] ),
    .B(_04123_),
    .X(_01256_));
 sky130_fd_sc_hd__nor3_2 _25056_ (.A(_04121_),
    .B(\timer[16] ),
    .C(_04095_),
    .Y(_04124_));
 sky130_fd_sc_hd__xor2_2 _25057_ (.A(\timer[17] ),
    .B(_04124_),
    .X(_01259_));
 sky130_fd_sc_hd__nand3b_2 _25058_ (.A_N(\timer[17] ),
    .B(_04123_),
    .C(_04085_),
    .Y(_04125_));
 sky130_fd_sc_hd__a22o_2 _25059_ (.A1(_04084_),
    .A2(_04124_),
    .B1(_04125_),
    .B2(\timer[18] ),
    .X(_01262_));
 sky130_fd_sc_hd__nand3_2 _25060_ (.A(_04123_),
    .B(_04085_),
    .C(_04084_),
    .Y(_04126_));
 sky130_vsdinv _25061_ (.A(_04123_),
    .Y(_04127_));
 sky130_fd_sc_hd__o2bb2ai_2 _25062_ (.A1_N(\timer[19] ),
    .A2_N(_04126_),
    .B1(_04127_),
    .B2(_04086_),
    .Y(_01265_));
 sky130_fd_sc_hd__xor2_2 _25063_ (.A(\timer[20] ),
    .B(_04096_),
    .X(_01268_));
 sky130_fd_sc_hd__or2b_2 _25064_ (.A(\timer[20] ),
    .B_N(_04096_),
    .X(_04128_));
 sky130_vsdinv _25065_ (.A(_04096_),
    .Y(_04129_));
 sky130_vsdinv _25066_ (.A(_04097_),
    .Y(_04130_));
 sky130_fd_sc_hd__o2bb2ai_2 _25067_ (.A1_N(\timer[21] ),
    .A2_N(_04128_),
    .B1(_04129_),
    .B2(_04130_),
    .Y(_01271_));
 sky130_fd_sc_hd__nand3b_2 _25068_ (.A_N(_04086_),
    .B(_04122_),
    .C(_04097_),
    .Y(_04131_));
 sky130_fd_sc_hd__xnor2_2 _25069_ (.A(\timer[22] ),
    .B(_04131_),
    .Y(_01274_));
 sky130_fd_sc_hd__buf_1 _25070_ (.A(\timer[23] ),
    .X(_04132_));
 sky130_fd_sc_hd__xnor2_2 _25071_ (.A(_04132_),
    .B(_04098_),
    .Y(_01277_));
 sky130_fd_sc_hd__nor2_2 _25072_ (.A(_04132_),
    .B(_04098_),
    .Y(_04133_));
 sky130_fd_sc_hd__xor2_2 _25073_ (.A(\timer[24] ),
    .B(_04133_),
    .X(_01280_));
 sky130_fd_sc_hd__nor3_2 _25074_ (.A(_04132_),
    .B(\timer[24] ),
    .C(_04098_),
    .Y(_04134_));
 sky130_fd_sc_hd__xor2_2 _25075_ (.A(\timer[25] ),
    .B(_04134_),
    .X(_01283_));
 sky130_fd_sc_hd__nand3b_2 _25076_ (.A_N(\timer[25] ),
    .B(_04133_),
    .C(_04082_),
    .Y(_04135_));
 sky130_fd_sc_hd__a22o_2 _25077_ (.A1(_04081_),
    .A2(_04134_),
    .B1(_04135_),
    .B2(\timer[26] ),
    .X(_01286_));
 sky130_fd_sc_hd__nand3_2 _25078_ (.A(_04133_),
    .B(_04082_),
    .C(_04081_),
    .Y(_04136_));
 sky130_vsdinv _25079_ (.A(_04133_),
    .Y(_04137_));
 sky130_fd_sc_hd__o2bb2ai_2 _25080_ (.A1_N(\timer[27] ),
    .A2_N(_04136_),
    .B1(_04137_),
    .B2(_04083_),
    .Y(_01289_));
 sky130_fd_sc_hd__xor2_2 _25081_ (.A(\timer[28] ),
    .B(_04099_),
    .X(_01292_));
 sky130_fd_sc_hd__or2b_2 _25082_ (.A(\timer[28] ),
    .B_N(_04099_),
    .X(_04138_));
 sky130_fd_sc_hd__and2_2 _25083_ (.A(_04099_),
    .B(_04100_),
    .X(_04139_));
 sky130_fd_sc_hd__a21o_2 _25084_ (.A1(_04138_),
    .A2(\timer[29] ),
    .B1(_04139_),
    .X(_01295_));
 sky130_fd_sc_hd__xor2_2 _25085_ (.A(\timer[30] ),
    .B(_04139_),
    .X(_01298_));
 sky130_fd_sc_hd__xnor2_2 _25086_ (.A(\timer[31] ),
    .B(_04101_),
    .Y(_01301_));
 sky130_fd_sc_hd__nor2b_2 _25087_ (.A(_18909_),
    .B_N(_19413_),
    .Y(_01315_));
 sky130_fd_sc_hd__nor2b_2 _25088_ (.A(_18909_),
    .B_N(_19415_),
    .Y(_01317_));
 sky130_fd_sc_hd__nor2b_2 _25089_ (.A(_18909_),
    .B_N(_19419_),
    .Y(_01319_));
 sky130_fd_sc_hd__buf_1 _25090_ (.A(_18908_),
    .X(_04140_));
 sky130_fd_sc_hd__buf_1 _25091_ (.A(_04140_),
    .X(_04141_));
 sky130_fd_sc_hd__nor2b_2 _25092_ (.A(_04141_),
    .B_N(_19422_),
    .Y(_01321_));
 sky130_fd_sc_hd__nor2b_2 _25093_ (.A(_04141_),
    .B_N(_19425_),
    .Y(_01323_));
 sky130_fd_sc_hd__nor2b_2 _25094_ (.A(_04141_),
    .B_N(_19427_),
    .Y(_01325_));
 sky130_fd_sc_hd__nor2b_2 _25095_ (.A(_04141_),
    .B_N(_19429_),
    .Y(_01327_));
 sky130_fd_sc_hd__buf_1 _25096_ (.A(_04140_),
    .X(_04142_));
 sky130_fd_sc_hd__nor2b_2 _25097_ (.A(_04142_),
    .B_N(_19440_),
    .Y(_01329_));
 sky130_fd_sc_hd__nor2b_2 _25098_ (.A(_04142_),
    .B_N(_19444_),
    .Y(_01331_));
 sky130_fd_sc_hd__nor2b_2 _25099_ (.A(_04142_),
    .B_N(_19445_),
    .Y(_01333_));
 sky130_fd_sc_hd__nor2b_2 _25100_ (.A(_04142_),
    .B_N(_19454_),
    .Y(_01335_));
 sky130_fd_sc_hd__buf_1 _25101_ (.A(_04140_),
    .X(_04143_));
 sky130_fd_sc_hd__nor2b_2 _25102_ (.A(_04143_),
    .B_N(_19458_),
    .Y(_01337_));
 sky130_fd_sc_hd__nor2b_2 _25103_ (.A(_04143_),
    .B_N(_19462_),
    .Y(_01339_));
 sky130_fd_sc_hd__nor2b_2 _25104_ (.A(_04143_),
    .B_N(_19465_),
    .Y(_01341_));
 sky130_fd_sc_hd__nor2b_2 _25105_ (.A(_04143_),
    .B_N(_19468_),
    .Y(_01343_));
 sky130_fd_sc_hd__buf_1 _25106_ (.A(_04140_),
    .X(_04144_));
 sky130_fd_sc_hd__buf_1 _25107_ (.A(\decoded_imm[20] ),
    .X(_04145_));
 sky130_fd_sc_hd__nor2b_2 _25108_ (.A(_04144_),
    .B_N(_04145_),
    .Y(_01345_));
 sky130_fd_sc_hd__nor2b_2 _25109_ (.A(_04144_),
    .B_N(_19483_),
    .Y(_01347_));
 sky130_fd_sc_hd__buf_1 _25110_ (.A(\decoded_imm[22] ),
    .X(_04146_));
 sky130_fd_sc_hd__nor2b_2 _25111_ (.A(_04144_),
    .B_N(_04146_),
    .Y(_01349_));
 sky130_fd_sc_hd__nor2b_2 _25112_ (.A(_04144_),
    .B_N(_19489_),
    .Y(_01351_));
 sky130_fd_sc_hd__buf_1 _25113_ (.A(_18908_),
    .X(_04147_));
 sky130_fd_sc_hd__nor2b_2 _25114_ (.A(_04147_),
    .B_N(_19491_),
    .Y(_01353_));
 sky130_fd_sc_hd__nor2b_2 _25115_ (.A(_04147_),
    .B_N(_19496_),
    .Y(_01355_));
 sky130_fd_sc_hd__nor2b_2 _25116_ (.A(_04147_),
    .B_N(_19499_),
    .Y(_01357_));
 sky130_fd_sc_hd__nor2b_2 _25117_ (.A(_04147_),
    .B_N(_19501_),
    .Y(_01359_));
 sky130_fd_sc_hd__buf_1 _25118_ (.A(_18908_),
    .X(_04148_));
 sky130_fd_sc_hd__nor2b_2 _25119_ (.A(_04148_),
    .B_N(_19504_),
    .Y(_01361_));
 sky130_fd_sc_hd__nor2b_2 _25120_ (.A(_04148_),
    .B_N(_19508_),
    .Y(_01363_));
 sky130_fd_sc_hd__nor2b_2 _25121_ (.A(_04148_),
    .B_N(_19510_),
    .Y(_01365_));
 sky130_fd_sc_hd__nor2b_2 _25122_ (.A(_04148_),
    .B_N(\decoded_imm[31] ),
    .Y(_01367_));
 sky130_fd_sc_hd__buf_1 _25123_ (.A(_19024_),
    .X(_04149_));
 sky130_fd_sc_hd__nor2b_2 _25124_ (.A(_04149_),
    .B_N(_19382_),
    .Y(_01369_));
 sky130_fd_sc_hd__xor2_2 _25125_ (.A(_18941_),
    .B(_19124_),
    .X(_01371_));
 sky130_fd_sc_hd__nor2b_2 _25126_ (.A(_04149_),
    .B_N(_17594_),
    .Y(_01372_));
 sky130_fd_sc_hd__and2_2 _25127_ (.A(\decoded_imm[0] ),
    .B(pcpi_rs1[0]),
    .X(_04150_));
 sky130_fd_sc_hd__xor2_2 _25128_ (.A(_19114_),
    .B(\decoded_imm[1] ),
    .X(_04151_));
 sky130_fd_sc_hd__xor2_2 _25129_ (.A(_04150_),
    .B(_04151_),
    .X(_01374_));
 sky130_fd_sc_hd__nor2b_2 _25130_ (.A(_04149_),
    .B_N(_17591_),
    .Y(_01375_));
 sky130_fd_sc_hd__xor2_2 _25131_ (.A(_19113_),
    .B(_19400_),
    .X(_04152_));
 sky130_fd_sc_hd__and2_2 _25132_ (.A(_19114_),
    .B(_19397_),
    .X(_04153_));
 sky130_fd_sc_hd__a21o_2 _25133_ (.A1(_04151_),
    .A2(_04150_),
    .B1(_04153_),
    .X(_04154_));
 sky130_fd_sc_hd__xor2_2 _25134_ (.A(_04152_),
    .B(_04154_),
    .X(_01377_));
 sky130_fd_sc_hd__nor2b_2 _25135_ (.A(_04149_),
    .B_N(_17585_),
    .Y(_01378_));
 sky130_fd_sc_hd__nor2_2 _25136_ (.A(_19109_),
    .B(_19404_),
    .Y(_04155_));
 sky130_fd_sc_hd__and2_2 _25137_ (.A(pcpi_rs1[3]),
    .B(\decoded_imm[3] ),
    .X(_04156_));
 sky130_fd_sc_hd__nor2_2 _25138_ (.A(_04155_),
    .B(_04156_),
    .Y(_04157_));
 sky130_fd_sc_hd__o21ai_2 _25139_ (.A1(pcpi_rs1[2]),
    .A2(\decoded_imm[2] ),
    .B1(_04154_),
    .Y(_04158_));
 sky130_fd_sc_hd__nand2_2 _25140_ (.A(_19112_),
    .B(\decoded_imm[2] ),
    .Y(_04159_));
 sky130_fd_sc_hd__nand2_2 _25141_ (.A(_04158_),
    .B(_04159_),
    .Y(_04160_));
 sky130_fd_sc_hd__xor2_2 _25142_ (.A(_04157_),
    .B(_04160_),
    .X(_01380_));
 sky130_fd_sc_hd__buf_1 _25143_ (.A(_19024_),
    .X(_04161_));
 sky130_fd_sc_hd__nor2b_2 _25144_ (.A(_04161_),
    .B_N(_17581_),
    .Y(_01381_));
 sky130_fd_sc_hd__xor2_2 _25145_ (.A(_19108_),
    .B(_19407_),
    .X(_04162_));
 sky130_vsdinv _25146_ (.A(_04155_),
    .Y(_04163_));
 sky130_fd_sc_hd__a21o_2 _25147_ (.A1(_04160_),
    .A2(_04163_),
    .B1(_04156_),
    .X(_04164_));
 sky130_fd_sc_hd__xor2_2 _25148_ (.A(_04162_),
    .B(_04164_),
    .X(_01383_));
 sky130_fd_sc_hd__nor2b_2 _25149_ (.A(_04161_),
    .B_N(_17575_),
    .Y(_01384_));
 sky130_fd_sc_hd__nor2_2 _25150_ (.A(_19104_),
    .B(\decoded_imm[5] ),
    .Y(_04165_));
 sky130_fd_sc_hd__and2_2 _25151_ (.A(pcpi_rs1[5]),
    .B(\decoded_imm[5] ),
    .X(_04166_));
 sky130_fd_sc_hd__nor2_2 _25152_ (.A(_04165_),
    .B(_04166_),
    .Y(_04167_));
 sky130_fd_sc_hd__or2_2 _25153_ (.A(pcpi_rs1[4]),
    .B(\decoded_imm[4] ),
    .X(_04168_));
 sky130_fd_sc_hd__nand2_2 _25154_ (.A(_04164_),
    .B(_04168_),
    .Y(_04169_));
 sky130_fd_sc_hd__nand2_2 _25155_ (.A(_19106_),
    .B(\decoded_imm[4] ),
    .Y(_04170_));
 sky130_fd_sc_hd__nand2_2 _25156_ (.A(_04169_),
    .B(_04170_),
    .Y(_04171_));
 sky130_fd_sc_hd__xor2_2 _25157_ (.A(_04167_),
    .B(_04171_),
    .X(_01386_));
 sky130_fd_sc_hd__nor2b_2 _25158_ (.A(_04161_),
    .B_N(_17571_),
    .Y(_01387_));
 sky130_fd_sc_hd__xor2_2 _25159_ (.A(_19101_),
    .B(\decoded_imm[6] ),
    .X(_04172_));
 sky130_vsdinv _25160_ (.A(_04165_),
    .Y(_04173_));
 sky130_fd_sc_hd__a21o_2 _25161_ (.A1(_04171_),
    .A2(_04173_),
    .B1(_04166_),
    .X(_04174_));
 sky130_fd_sc_hd__xor2_2 _25162_ (.A(_04172_),
    .B(_04174_),
    .X(_01389_));
 sky130_fd_sc_hd__nor2b_2 _25163_ (.A(_04161_),
    .B_N(_17567_),
    .Y(_01390_));
 sky130_fd_sc_hd__xnor2_2 _25164_ (.A(pcpi_rs1[7]),
    .B(\decoded_imm[7] ),
    .Y(_04175_));
 sky130_fd_sc_hd__and2_2 _25165_ (.A(_19103_),
    .B(_19415_),
    .X(_04176_));
 sky130_fd_sc_hd__a21oi_2 _25166_ (.A1(_04174_),
    .A2(_04172_),
    .B1(_04176_),
    .Y(_04177_));
 sky130_fd_sc_hd__xor2_2 _25167_ (.A(_04175_),
    .B(_04177_),
    .X(_01392_));
 sky130_fd_sc_hd__buf_1 _25168_ (.A(_19024_),
    .X(_04178_));
 sky130_fd_sc_hd__nor2b_2 _25169_ (.A(_04178_),
    .B_N(\reg_pc[8] ),
    .Y(_01393_));
 sky130_fd_sc_hd__nor2_2 _25170_ (.A(_19094_),
    .B(\decoded_imm[8] ),
    .Y(_04179_));
 sky130_fd_sc_hd__and2_2 _25171_ (.A(pcpi_rs1[8]),
    .B(\decoded_imm[8] ),
    .X(_04180_));
 sky130_fd_sc_hd__nor2_2 _25172_ (.A(_04179_),
    .B(_04180_),
    .Y(_04181_));
 sky130_fd_sc_hd__and2b_2 _25173_ (.A_N(_04175_),
    .B(_04172_),
    .X(_04182_));
 sky130_fd_sc_hd__o211ai_2 _25174_ (.A1(_19097_),
    .A2(\decoded_imm[7] ),
    .B1(_19101_),
    .C1(\decoded_imm[6] ),
    .Y(_04183_));
 sky130_fd_sc_hd__nand2_2 _25175_ (.A(_19097_),
    .B(\decoded_imm[7] ),
    .Y(_04184_));
 sky130_fd_sc_hd__and2_2 _25176_ (.A(_04183_),
    .B(_04184_),
    .X(_04185_));
 sky130_fd_sc_hd__a21boi_2 _25177_ (.A1(_04174_),
    .A2(_04182_),
    .B1_N(_04185_),
    .Y(_04186_));
 sky130_fd_sc_hd__xnor2_2 _25178_ (.A(_04181_),
    .B(_04186_),
    .Y(_01395_));
 sky130_fd_sc_hd__nor2b_2 _25179_ (.A(_04178_),
    .B_N(_17558_),
    .Y(_01396_));
 sky130_fd_sc_hd__nor2_2 _25180_ (.A(_19091_),
    .B(\decoded_imm[9] ),
    .Y(_04187_));
 sky130_fd_sc_hd__and2_2 _25181_ (.A(pcpi_rs1[9]),
    .B(\decoded_imm[9] ),
    .X(_04188_));
 sky130_fd_sc_hd__nor2_2 _25182_ (.A(_04187_),
    .B(_04188_),
    .Y(_04189_));
 sky130_fd_sc_hd__o21bai_2 _25183_ (.A1(_04179_),
    .A2(_04186_),
    .B1_N(_04180_),
    .Y(_04190_));
 sky130_fd_sc_hd__xor2_2 _25184_ (.A(_04189_),
    .B(_04190_),
    .X(_01398_));
 sky130_fd_sc_hd__nor2b_2 _25185_ (.A(_04178_),
    .B_N(_17553_),
    .Y(_01399_));
 sky130_fd_sc_hd__xor2_2 _25186_ (.A(pcpi_rs1[10]),
    .B(\decoded_imm[10] ),
    .X(_04191_));
 sky130_fd_sc_hd__nand2_2 _25187_ (.A(_04181_),
    .B(_04189_),
    .Y(_04192_));
 sky130_fd_sc_hd__o211ai_2 _25188_ (.A1(_19091_),
    .A2(\decoded_imm[9] ),
    .B1(_19094_),
    .C1(\decoded_imm[8] ),
    .Y(_04193_));
 sky130_fd_sc_hd__or2b_2 _25189_ (.A(_04188_),
    .B_N(_04193_),
    .X(_04194_));
 sky130_fd_sc_hd__o21bai_2 _25190_ (.A1(_04192_),
    .A2(_04186_),
    .B1_N(_04194_),
    .Y(_04195_));
 sky130_fd_sc_hd__xor2_2 _25191_ (.A(_04191_),
    .B(_04195_),
    .X(_01401_));
 sky130_fd_sc_hd__nor2b_2 _25192_ (.A(_04178_),
    .B_N(_17549_),
    .Y(_01402_));
 sky130_fd_sc_hd__xor2_2 _25193_ (.A(pcpi_rs1[11]),
    .B(\decoded_imm[11] ),
    .X(_04196_));
 sky130_fd_sc_hd__nand2_2 _25194_ (.A(_04195_),
    .B(_04191_),
    .Y(_04197_));
 sky130_fd_sc_hd__nand2_2 _25195_ (.A(_19089_),
    .B(\decoded_imm[10] ),
    .Y(_04198_));
 sky130_fd_sc_hd__nand2_2 _25196_ (.A(_04197_),
    .B(_04198_),
    .Y(_04199_));
 sky130_fd_sc_hd__xor2_2 _25197_ (.A(_04196_),
    .B(_04199_),
    .X(_01404_));
 sky130_fd_sc_hd__buf_1 _25198_ (.A(instr_lui),
    .X(_04200_));
 sky130_fd_sc_hd__buf_1 _25199_ (.A(_04200_),
    .X(_04201_));
 sky130_fd_sc_hd__nor2b_2 _25200_ (.A(_04201_),
    .B_N(_17545_),
    .Y(_01405_));
 sky130_fd_sc_hd__xor2_2 _25201_ (.A(pcpi_rs1[12]),
    .B(\decoded_imm[12] ),
    .X(_04202_));
 sky130_fd_sc_hd__nand2_2 _25202_ (.A(_04199_),
    .B(_04196_),
    .Y(_04203_));
 sky130_fd_sc_hd__and2_2 _25203_ (.A(pcpi_rs1[11]),
    .B(\decoded_imm[11] ),
    .X(_04204_));
 sky130_vsdinv _25204_ (.A(_04204_),
    .Y(_04205_));
 sky130_fd_sc_hd__nand2_2 _25205_ (.A(_04203_),
    .B(_04205_),
    .Y(_04206_));
 sky130_fd_sc_hd__xor2_2 _25206_ (.A(_04202_),
    .B(_04206_),
    .X(_01407_));
 sky130_fd_sc_hd__nor2b_2 _25207_ (.A(_04201_),
    .B_N(_17539_),
    .Y(_01408_));
 sky130_fd_sc_hd__xnor2_2 _25208_ (.A(pcpi_rs1[13]),
    .B(\decoded_imm[13] ),
    .Y(_04207_));
 sky130_fd_sc_hd__and2_2 _25209_ (.A(_19084_),
    .B(\decoded_imm[12] ),
    .X(_04208_));
 sky130_fd_sc_hd__a21oi_2 _25210_ (.A1(_04206_),
    .A2(_04202_),
    .B1(_04208_),
    .Y(_04209_));
 sky130_fd_sc_hd__xor2_2 _25211_ (.A(_04207_),
    .B(_04209_),
    .X(_01410_));
 sky130_fd_sc_hd__nor2b_2 _25212_ (.A(_04201_),
    .B_N(_17536_),
    .Y(_01411_));
 sky130_fd_sc_hd__xor2_2 _25213_ (.A(pcpi_rs1[14]),
    .B(\decoded_imm[14] ),
    .X(_04210_));
 sky130_fd_sc_hd__and2_2 _25214_ (.A(pcpi_rs1[13]),
    .B(\decoded_imm[13] ),
    .X(_04211_));
 sky130_fd_sc_hd__o21bai_2 _25215_ (.A1(_04207_),
    .A2(_04209_),
    .B1_N(_04211_),
    .Y(_04212_));
 sky130_fd_sc_hd__xor2_2 _25216_ (.A(_04210_),
    .B(_04212_),
    .X(_01413_));
 sky130_fd_sc_hd__nor2b_2 _25217_ (.A(_04201_),
    .B_N(_17530_),
    .Y(_01414_));
 sky130_fd_sc_hd__xnor2_2 _25218_ (.A(pcpi_rs1[15]),
    .B(\decoded_imm[15] ),
    .Y(_04213_));
 sky130_fd_sc_hd__and2_2 _25219_ (.A(_19080_),
    .B(\decoded_imm[14] ),
    .X(_04214_));
 sky130_fd_sc_hd__a21oi_2 _25220_ (.A1(_04212_),
    .A2(_04210_),
    .B1(_04214_),
    .Y(_04215_));
 sky130_fd_sc_hd__xor2_2 _25221_ (.A(_04213_),
    .B(_04215_),
    .X(_01416_));
 sky130_fd_sc_hd__buf_1 _25222_ (.A(_04200_),
    .X(_04216_));
 sky130_fd_sc_hd__nor2b_2 _25223_ (.A(_04216_),
    .B_N(_17526_),
    .Y(_01417_));
 sky130_fd_sc_hd__xor2_2 _25224_ (.A(pcpi_rs1[16]),
    .B(\decoded_imm[16] ),
    .X(_04217_));
 sky130_fd_sc_hd__and2_2 _25225_ (.A(pcpi_rs1[15]),
    .B(\decoded_imm[15] ),
    .X(_04218_));
 sky130_fd_sc_hd__o21bai_2 _25226_ (.A1(_04213_),
    .A2(_04215_),
    .B1_N(_04218_),
    .Y(_04219_));
 sky130_fd_sc_hd__xor2_2 _25227_ (.A(_04217_),
    .B(_04219_),
    .X(_01419_));
 sky130_fd_sc_hd__nor2b_2 _25228_ (.A(_04216_),
    .B_N(_17524_),
    .Y(_01420_));
 sky130_fd_sc_hd__xnor2_2 _25229_ (.A(pcpi_rs1[17]),
    .B(\decoded_imm[17] ),
    .Y(_04220_));
 sky130_fd_sc_hd__and2_2 _25230_ (.A(_19075_),
    .B(_19458_),
    .X(_04221_));
 sky130_fd_sc_hd__a21oi_2 _25231_ (.A1(_04219_),
    .A2(_04217_),
    .B1(_04221_),
    .Y(_04222_));
 sky130_fd_sc_hd__xor2_2 _25232_ (.A(_04220_),
    .B(_04222_),
    .X(_01422_));
 sky130_fd_sc_hd__nor2b_2 _25233_ (.A(_04216_),
    .B_N(_17516_),
    .Y(_01423_));
 sky130_fd_sc_hd__nor2_2 _25234_ (.A(_19068_),
    .B(_19465_),
    .Y(_04223_));
 sky130_fd_sc_hd__and2_2 _25235_ (.A(pcpi_rs1[18]),
    .B(\decoded_imm[18] ),
    .X(_04224_));
 sky130_fd_sc_hd__nor2_2 _25236_ (.A(_04223_),
    .B(_04224_),
    .Y(_04225_));
 sky130_fd_sc_hd__and2b_2 _25237_ (.A_N(_04220_),
    .B(_04217_),
    .X(_04226_));
 sky130_fd_sc_hd__o211a_2 _25238_ (.A1(_19070_),
    .A2(\decoded_imm[17] ),
    .B1(_19073_),
    .C1(\decoded_imm[16] ),
    .X(_04227_));
 sky130_fd_sc_hd__a21o_2 _25239_ (.A1(_19070_),
    .A2(_19462_),
    .B1(_04227_),
    .X(_04228_));
 sky130_fd_sc_hd__a21oi_2 _25240_ (.A1(_04219_),
    .A2(_04226_),
    .B1(_04228_),
    .Y(_04229_));
 sky130_fd_sc_hd__xnor2_2 _25241_ (.A(_04225_),
    .B(_04229_),
    .Y(_01425_));
 sky130_fd_sc_hd__nor2b_2 _25242_ (.A(_04216_),
    .B_N(_17510_),
    .Y(_01426_));
 sky130_fd_sc_hd__xor2_2 _25243_ (.A(pcpi_rs1[19]),
    .B(\decoded_imm[19] ),
    .X(_04230_));
 sky130_fd_sc_hd__o21bai_2 _25244_ (.A1(_04223_),
    .A2(_04229_),
    .B1_N(_04224_),
    .Y(_04231_));
 sky130_fd_sc_hd__xor2_2 _25245_ (.A(_04230_),
    .B(_04231_),
    .X(_01428_));
 sky130_fd_sc_hd__buf_1 _25246_ (.A(_04200_),
    .X(_04232_));
 sky130_fd_sc_hd__buf_1 _25247_ (.A(\reg_pc[20] ),
    .X(_04233_));
 sky130_fd_sc_hd__nor2b_2 _25248_ (.A(_04232_),
    .B_N(_04233_),
    .Y(_01429_));
 sky130_fd_sc_hd__xnor2_2 _25249_ (.A(pcpi_rs1[20]),
    .B(_04145_),
    .Y(_04234_));
 sky130_fd_sc_hd__and2_2 _25250_ (.A(_19065_),
    .B(_19468_),
    .X(_04235_));
 sky130_fd_sc_hd__a21oi_2 _25251_ (.A1(_04231_),
    .A2(_04230_),
    .B1(_04235_),
    .Y(_04236_));
 sky130_fd_sc_hd__xor2_2 _25252_ (.A(_04234_),
    .B(_04236_),
    .X(_01431_));
 sky130_fd_sc_hd__nor2b_2 _25253_ (.A(_04232_),
    .B_N(_17503_),
    .Y(_01432_));
 sky130_fd_sc_hd__xor2_2 _25254_ (.A(pcpi_rs1[21]),
    .B(\decoded_imm[21] ),
    .X(_04237_));
 sky130_fd_sc_hd__and2_2 _25255_ (.A(_19063_),
    .B(_04145_),
    .X(_04238_));
 sky130_fd_sc_hd__o21bai_2 _25256_ (.A1(_04234_),
    .A2(_04236_),
    .B1_N(_04238_),
    .Y(_04239_));
 sky130_fd_sc_hd__xor2_2 _25257_ (.A(_04237_),
    .B(_04239_),
    .X(_01434_));
 sky130_fd_sc_hd__buf_1 _25258_ (.A(\reg_pc[22] ),
    .X(_04240_));
 sky130_fd_sc_hd__nor2b_2 _25259_ (.A(_04232_),
    .B_N(_04240_),
    .Y(_01435_));
 sky130_fd_sc_hd__xnor2_2 _25260_ (.A(pcpi_rs1[22]),
    .B(_04146_),
    .Y(_04241_));
 sky130_fd_sc_hd__and2_2 _25261_ (.A(_19061_),
    .B(_19483_),
    .X(_04242_));
 sky130_fd_sc_hd__a21oi_2 _25262_ (.A1(_04239_),
    .A2(_04237_),
    .B1(_04242_),
    .Y(_04243_));
 sky130_fd_sc_hd__xor2_2 _25263_ (.A(_04241_),
    .B(_04243_),
    .X(_01437_));
 sky130_fd_sc_hd__nor2b_2 _25264_ (.A(_04232_),
    .B_N(_17492_),
    .Y(_01438_));
 sky130_fd_sc_hd__xor2_2 _25265_ (.A(pcpi_rs1[23]),
    .B(\decoded_imm[23] ),
    .X(_04244_));
 sky130_fd_sc_hd__and2_2 _25266_ (.A(_19059_),
    .B(_04146_),
    .X(_04245_));
 sky130_fd_sc_hd__o21bai_2 _25267_ (.A1(_04241_),
    .A2(_04243_),
    .B1_N(_04245_),
    .Y(_04246_));
 sky130_fd_sc_hd__xor2_2 _25268_ (.A(_04244_),
    .B(_04246_),
    .X(_01440_));
 sky130_fd_sc_hd__buf_1 _25269_ (.A(_04200_),
    .X(_04247_));
 sky130_fd_sc_hd__nor2b_2 _25270_ (.A(_04247_),
    .B_N(_17489_),
    .Y(_01441_));
 sky130_fd_sc_hd__xor2_2 _25271_ (.A(_19703_),
    .B(\decoded_imm[24] ),
    .X(_04248_));
 sky130_fd_sc_hd__and2_2 _25272_ (.A(_19056_),
    .B(_19489_),
    .X(_04249_));
 sky130_fd_sc_hd__a21oi_2 _25273_ (.A1(_04246_),
    .A2(_04244_),
    .B1(_04249_),
    .Y(_04250_));
 sky130_fd_sc_hd__xnor2_2 _25274_ (.A(_04248_),
    .B(_04250_),
    .Y(_01443_));
 sky130_fd_sc_hd__nor2b_2 _25275_ (.A(_04247_),
    .B_N(_17484_),
    .Y(_01444_));
 sky130_fd_sc_hd__buf_1 _25276_ (.A(_19052_),
    .X(_04251_));
 sky130_fd_sc_hd__xor2_2 _25277_ (.A(_04251_),
    .B(_19496_),
    .X(_04252_));
 sky130_fd_sc_hd__and2b_2 _25278_ (.A_N(_04250_),
    .B(_04248_),
    .X(_04253_));
 sky130_fd_sc_hd__a21oi_2 _25279_ (.A1(_19055_),
    .A2(_19491_),
    .B1(_04253_),
    .Y(_04254_));
 sky130_fd_sc_hd__xnor2_2 _25280_ (.A(_04252_),
    .B(_04254_),
    .Y(_01446_));
 sky130_fd_sc_hd__nor2b_2 _25281_ (.A(_04247_),
    .B_N(_17480_),
    .Y(_01447_));
 sky130_fd_sc_hd__xor2_2 _25282_ (.A(_19701_),
    .B(\decoded_imm[26] ),
    .X(_04255_));
 sky130_fd_sc_hd__nand2_2 _25283_ (.A(_04248_),
    .B(_04252_),
    .Y(_04256_));
 sky130_vsdinv _25284_ (.A(_04251_),
    .Y(_04257_));
 sky130_fd_sc_hd__o211ai_2 _25285_ (.A1(_04251_),
    .A2(_19496_),
    .B1(_19054_),
    .C1(_19491_),
    .Y(_04258_));
 sky130_fd_sc_hd__o21ai_2 _25286_ (.A1(_04257_),
    .A2(_19497_),
    .B1(_04258_),
    .Y(_04259_));
 sky130_fd_sc_hd__o21bai_2 _25287_ (.A1(_04256_),
    .A2(_04250_),
    .B1_N(_04259_),
    .Y(_04260_));
 sky130_fd_sc_hd__xor2_2 _25288_ (.A(_04255_),
    .B(_04260_),
    .X(_01449_));
 sky130_fd_sc_hd__nor2b_2 _25289_ (.A(_04247_),
    .B_N(_17476_),
    .Y(_01450_));
 sky130_fd_sc_hd__buf_1 _25290_ (.A(pcpi_rs1[27]),
    .X(_04261_));
 sky130_fd_sc_hd__xnor2_2 _25291_ (.A(_04261_),
    .B(\decoded_imm[27] ),
    .Y(_04262_));
 sky130_fd_sc_hd__and2_2 _25292_ (.A(_19051_),
    .B(_19499_),
    .X(_04263_));
 sky130_fd_sc_hd__a21oi_2 _25293_ (.A1(_04260_),
    .A2(_04255_),
    .B1(_04263_),
    .Y(_04264_));
 sky130_fd_sc_hd__xor2_2 _25294_ (.A(_04262_),
    .B(_04264_),
    .X(_01452_));
 sky130_fd_sc_hd__buf_1 _25295_ (.A(instr_lui),
    .X(_04265_));
 sky130_fd_sc_hd__nor2b_2 _25296_ (.A(_04265_),
    .B_N(_17471_),
    .Y(_01453_));
 sky130_fd_sc_hd__xnor2_2 _25297_ (.A(_19046_),
    .B(_19504_),
    .Y(_04266_));
 sky130_fd_sc_hd__and2b_2 _25298_ (.A_N(_04262_),
    .B(_04255_),
    .X(_04267_));
 sky130_fd_sc_hd__o211ai_2 _25299_ (.A1(_04261_),
    .A2(_19501_),
    .B1(_19701_),
    .C1(_19499_),
    .Y(_04268_));
 sky130_fd_sc_hd__nand2_2 _25300_ (.A(_19047_),
    .B(_19501_),
    .Y(_04269_));
 sky130_fd_sc_hd__and2_2 _25301_ (.A(_04268_),
    .B(_04269_),
    .X(_04270_));
 sky130_fd_sc_hd__a21boi_2 _25302_ (.A1(_04260_),
    .A2(_04267_),
    .B1_N(_04270_),
    .Y(_04271_));
 sky130_fd_sc_hd__xor2_2 _25303_ (.A(_04266_),
    .B(_04271_),
    .X(_01455_));
 sky130_fd_sc_hd__nor2b_2 _25304_ (.A(_04265_),
    .B_N(_17467_),
    .Y(_01456_));
 sky130_fd_sc_hd__xor2_2 _25305_ (.A(_19044_),
    .B(_19508_),
    .X(_04272_));
 sky130_fd_sc_hd__nor2_2 _25306_ (.A(_19045_),
    .B(_19504_),
    .Y(_04273_));
 sky130_fd_sc_hd__and2_2 _25307_ (.A(_19045_),
    .B(\decoded_imm[28] ),
    .X(_04274_));
 sky130_fd_sc_hd__o21bai_2 _25308_ (.A1(_04273_),
    .A2(_04271_),
    .B1_N(_04274_),
    .Y(_04275_));
 sky130_fd_sc_hd__xor2_2 _25309_ (.A(_04272_),
    .B(_04275_),
    .X(_01458_));
 sky130_fd_sc_hd__nor2b_2 _25310_ (.A(_04265_),
    .B_N(_17465_),
    .Y(_01459_));
 sky130_fd_sc_hd__buf_1 _25311_ (.A(_19041_),
    .X(_04276_));
 sky130_fd_sc_hd__xnor2_2 _25312_ (.A(_04276_),
    .B(_19510_),
    .Y(_04277_));
 sky130_vsdinv _25313_ (.A(pcpi_rs1[29]),
    .Y(_04278_));
 sky130_fd_sc_hd__nand2_2 _25314_ (.A(_04278_),
    .B(_19509_),
    .Y(_04279_));
 sky130_fd_sc_hd__and2_2 _25315_ (.A(_19043_),
    .B(_19508_),
    .X(_04280_));
 sky130_fd_sc_hd__a21oi_2 _25316_ (.A1(_04275_),
    .A2(_04279_),
    .B1(_04280_),
    .Y(_04281_));
 sky130_fd_sc_hd__xor2_2 _25317_ (.A(_04277_),
    .B(_04281_),
    .X(_01461_));
 sky130_fd_sc_hd__nor2b_2 _25318_ (.A(_04265_),
    .B_N(\reg_pc[31] ),
    .Y(_01462_));
 sky130_fd_sc_hd__nor2_2 _25319_ (.A(_19042_),
    .B(_19510_),
    .Y(_04282_));
 sky130_fd_sc_hd__and2_2 _25320_ (.A(_04276_),
    .B(\decoded_imm[30] ),
    .X(_04283_));
 sky130_fd_sc_hd__o21bai_2 _25321_ (.A1(_04282_),
    .A2(_04281_),
    .B1_N(_04283_),
    .Y(_04284_));
 sky130_fd_sc_hd__xnor2_2 _25322_ (.A(_16957_),
    .B(\decoded_imm[31] ),
    .Y(_04285_));
 sky130_fd_sc_hd__nand2_2 _25323_ (.A(_04284_),
    .B(_04285_),
    .Y(_04286_));
 sky130_vsdinv _25324_ (.A(_04283_),
    .Y(_04287_));
 sky130_vsdinv _25325_ (.A(_04285_),
    .Y(_04288_));
 sky130_fd_sc_hd__o211ai_2 _25326_ (.A1(_04282_),
    .A2(_04281_),
    .B1(_04287_),
    .C1(_04288_),
    .Y(_04289_));
 sky130_fd_sc_hd__nand2_2 _25327_ (.A(_04286_),
    .B(_04289_),
    .Y(_01464_));
 sky130_fd_sc_hd__and2_2 _25328_ (.A(_04080_),
    .B(_01466_),
    .X(_01467_));
 sky130_fd_sc_hd__buf_1 _25329_ (.A(_16833_),
    .X(_04290_));
 sky130_fd_sc_hd__buf_1 _25330_ (.A(_04290_),
    .X(_04291_));
 sky130_fd_sc_hd__and2_2 _25331_ (.A(_04291_),
    .B(_01469_),
    .X(_01470_));
 sky130_vsdinv _25332_ (.A(\reg_next_pc[4] ),
    .Y(_01471_));
 sky130_fd_sc_hd__buf_1 _25333_ (.A(_17036_),
    .X(_04292_));
 sky130_fd_sc_hd__buf_1 _25334_ (.A(_04292_),
    .X(_04293_));
 sky130_fd_sc_hd__a21oi_2 _25335_ (.A1(_04080_),
    .A2(_01473_),
    .B1(_04293_),
    .Y(_01474_));
 sky130_fd_sc_hd__and2_2 _25336_ (.A(_04291_),
    .B(_01477_),
    .X(_01478_));
 sky130_fd_sc_hd__and2_2 _25337_ (.A(_04291_),
    .B(_01480_),
    .X(_01481_));
 sky130_fd_sc_hd__and2_2 _25338_ (.A(_04291_),
    .B(_01483_),
    .X(_01484_));
 sky130_fd_sc_hd__buf_1 _25339_ (.A(_04290_),
    .X(_04294_));
 sky130_fd_sc_hd__and2_2 _25340_ (.A(_04294_),
    .B(_01486_),
    .X(_01487_));
 sky130_fd_sc_hd__and2_2 _25341_ (.A(_04294_),
    .B(_01489_),
    .X(_01490_));
 sky130_fd_sc_hd__and2_2 _25342_ (.A(_04294_),
    .B(_01492_),
    .X(_01493_));
 sky130_fd_sc_hd__and2_2 _25343_ (.A(_04294_),
    .B(_01495_),
    .X(_01496_));
 sky130_fd_sc_hd__buf_1 _25344_ (.A(_04290_),
    .X(_04295_));
 sky130_fd_sc_hd__and2_2 _25345_ (.A(_04295_),
    .B(_01498_),
    .X(_01499_));
 sky130_fd_sc_hd__and2_2 _25346_ (.A(_04295_),
    .B(_01501_),
    .X(_01502_));
 sky130_fd_sc_hd__and2_2 _25347_ (.A(_04295_),
    .B(_01504_),
    .X(_01505_));
 sky130_fd_sc_hd__and2_2 _25348_ (.A(_04295_),
    .B(_01507_),
    .X(_01508_));
 sky130_fd_sc_hd__buf_1 _25349_ (.A(_04290_),
    .X(_04296_));
 sky130_fd_sc_hd__and2_2 _25350_ (.A(_04296_),
    .B(_01510_),
    .X(_01511_));
 sky130_fd_sc_hd__and2_2 _25351_ (.A(_04296_),
    .B(_01513_),
    .X(_01514_));
 sky130_fd_sc_hd__and2_2 _25352_ (.A(_04296_),
    .B(_01516_),
    .X(_01517_));
 sky130_fd_sc_hd__and2_2 _25353_ (.A(_04296_),
    .B(_01519_),
    .X(_01520_));
 sky130_fd_sc_hd__buf_1 _25354_ (.A(_04079_),
    .X(_04297_));
 sky130_fd_sc_hd__and2_2 _25355_ (.A(_04297_),
    .B(_01522_),
    .X(_01523_));
 sky130_fd_sc_hd__and2_2 _25356_ (.A(_04297_),
    .B(_01525_),
    .X(_01526_));
 sky130_fd_sc_hd__and2_2 _25357_ (.A(_04297_),
    .B(_01528_),
    .X(_01529_));
 sky130_fd_sc_hd__and2_2 _25358_ (.A(_04297_),
    .B(_01531_),
    .X(_01532_));
 sky130_fd_sc_hd__buf_1 _25359_ (.A(_04079_),
    .X(_04298_));
 sky130_fd_sc_hd__and2_2 _25360_ (.A(_04298_),
    .B(_01534_),
    .X(_01535_));
 sky130_fd_sc_hd__and2_2 _25361_ (.A(_04298_),
    .B(_01537_),
    .X(_01538_));
 sky130_fd_sc_hd__and2_2 _25362_ (.A(_04298_),
    .B(_01540_),
    .X(_01541_));
 sky130_fd_sc_hd__and2_2 _25363_ (.A(_04298_),
    .B(_01543_),
    .X(_01544_));
 sky130_fd_sc_hd__buf_1 _25364_ (.A(_04079_),
    .X(_04299_));
 sky130_fd_sc_hd__and2_2 _25365_ (.A(_04299_),
    .B(_01546_),
    .X(_01547_));
 sky130_fd_sc_hd__and2_2 _25366_ (.A(_04299_),
    .B(_01549_),
    .X(_01550_));
 sky130_fd_sc_hd__and2_2 _25367_ (.A(_04299_),
    .B(_01552_),
    .X(_01553_));
 sky130_fd_sc_hd__and2_2 _25368_ (.A(_04299_),
    .B(_01555_),
    .X(_01556_));
 sky130_fd_sc_hd__xor2_2 _25369_ (.A(_02590_),
    .B(_18935_),
    .X(_01557_));
 sky130_fd_sc_hd__and2_2 _25370_ (.A(_02590_),
    .B(_18935_),
    .X(_04300_));
 sky130_fd_sc_hd__xnor2_2 _25371_ (.A(_02560_),
    .B(\decoded_imm_uj[2] ),
    .Y(_04301_));
 sky130_fd_sc_hd__xnor2_2 _25372_ (.A(_04300_),
    .B(_04301_),
    .Y(_01562_));
 sky130_fd_sc_hd__xor2_2 _25373_ (.A(_01561_),
    .B(_02410_),
    .X(_01565_));
 sky130_fd_sc_hd__xor2_2 _25374_ (.A(_17587_),
    .B(_17592_),
    .X(_01567_));
 sky130_fd_sc_hd__xor2_2 _25375_ (.A(_17587_),
    .B(_18934_),
    .X(_04302_));
 sky130_fd_sc_hd__nand3b_2 _25376_ (.A_N(_04301_),
    .B(_02590_),
    .C(\decoded_imm_uj[1] ),
    .Y(_04303_));
 sky130_fd_sc_hd__nand2_2 _25377_ (.A(_02560_),
    .B(\decoded_imm_uj[2] ),
    .Y(_04304_));
 sky130_fd_sc_hd__nand2_2 _25378_ (.A(_04303_),
    .B(_04304_),
    .Y(_04305_));
 sky130_fd_sc_hd__xor2_2 _25379_ (.A(_04302_),
    .B(_04305_),
    .X(_01568_));
 sky130_fd_sc_hd__and2_2 _25380_ (.A(_17586_),
    .B(_17592_),
    .X(_04306_));
 sky130_fd_sc_hd__xor2_2 _25381_ (.A(_02582_),
    .B(_04306_),
    .X(_01571_));
 sky130_fd_sc_hd__xnor2_2 _25382_ (.A(_18932_),
    .B(_17579_),
    .Y(_04307_));
 sky130_fd_sc_hd__o2bb2ai_2 _25383_ (.A1_N(_04304_),
    .A2_N(_04303_),
    .B1(_02571_),
    .B2(\decoded_imm_uj[3] ),
    .Y(_04308_));
 sky130_fd_sc_hd__nand2_2 _25384_ (.A(_17586_),
    .B(_18934_),
    .Y(_04309_));
 sky130_fd_sc_hd__nand2_2 _25385_ (.A(_04308_),
    .B(_04309_),
    .Y(_04310_));
 sky130_fd_sc_hd__xor2_2 _25386_ (.A(_04307_),
    .B(_04310_),
    .X(_01572_));
 sky130_fd_sc_hd__buf_1 _25387_ (.A(_02583_),
    .X(_04311_));
 sky130_fd_sc_hd__and3b_2 _25388_ (.A_N(_17579_),
    .B(_17586_),
    .C(_02560_),
    .X(_04312_));
 sky130_fd_sc_hd__xor2_2 _25389_ (.A(_04311_),
    .B(_04312_),
    .X(_01575_));
 sky130_fd_sc_hd__xor2_2 _25390_ (.A(_04311_),
    .B(\decoded_imm_uj[5] ),
    .X(_04313_));
 sky130_fd_sc_hd__o2bb2ai_2 _25391_ (.A1_N(_04309_),
    .A2_N(_04308_),
    .B1(_18932_),
    .B2(_17583_),
    .Y(_04314_));
 sky130_fd_sc_hd__o21ai_2 _25392_ (.A1(_00367_),
    .A2(_17579_),
    .B1(_04314_),
    .Y(_04315_));
 sky130_fd_sc_hd__xor2_2 _25393_ (.A(_04313_),
    .B(_04315_),
    .X(_01576_));
 sky130_fd_sc_hd__and4_2 _25394_ (.A(_02582_),
    .B(_04311_),
    .C(_17587_),
    .D(_17592_),
    .X(_04316_));
 sky130_fd_sc_hd__xor2_2 _25395_ (.A(_17572_),
    .B(_04316_),
    .X(_01579_));
 sky130_fd_sc_hd__nor2_2 _25396_ (.A(_02584_),
    .B(\decoded_imm_uj[6] ),
    .Y(_04317_));
 sky130_fd_sc_hd__and2_2 _25397_ (.A(_02584_),
    .B(\decoded_imm_uj[6] ),
    .X(_04318_));
 sky130_fd_sc_hd__nor2_2 _25398_ (.A(_04317_),
    .B(_04318_),
    .Y(_04319_));
 sky130_fd_sc_hd__o21ai_2 _25399_ (.A1(_02583_),
    .A2(\decoded_imm_uj[5] ),
    .B1(_04315_),
    .Y(_04320_));
 sky130_fd_sc_hd__o21ai_2 _25400_ (.A1(_17577_),
    .A2(_19411_),
    .B1(_04320_),
    .Y(_04321_));
 sky130_fd_sc_hd__xor2_2 _25401_ (.A(_04319_),
    .B(_04321_),
    .X(_01580_));
 sky130_fd_sc_hd__buf_1 _25402_ (.A(_02585_),
    .X(_04322_));
 sky130_fd_sc_hd__and4_2 _25403_ (.A(_04306_),
    .B(_17572_),
    .C(_02583_),
    .D(_02582_),
    .X(_04323_));
 sky130_fd_sc_hd__xor2_2 _25404_ (.A(_04322_),
    .B(_04323_),
    .X(_01583_));
 sky130_fd_sc_hd__xor2_2 _25405_ (.A(_04322_),
    .B(\decoded_imm_uj[7] ),
    .X(_04324_));
 sky130_vsdinv _25406_ (.A(_04317_),
    .Y(_04325_));
 sky130_fd_sc_hd__a21o_2 _25407_ (.A1(_04321_),
    .A2(_04325_),
    .B1(_04318_),
    .X(_04326_));
 sky130_fd_sc_hd__xor2_2 _25408_ (.A(_04324_),
    .B(_04326_),
    .X(_01584_));
 sky130_fd_sc_hd__and4_2 _25409_ (.A(_04312_),
    .B(_02585_),
    .C(_02584_),
    .D(_04311_),
    .X(_04327_));
 sky130_fd_sc_hd__xor2_2 _25410_ (.A(_17564_),
    .B(_04327_),
    .X(_01587_));
 sky130_fd_sc_hd__xnor2_2 _25411_ (.A(_17564_),
    .B(_18930_),
    .Y(_04328_));
 sky130_fd_sc_hd__nand2_2 _25412_ (.A(_17568_),
    .B(_19417_),
    .Y(_04329_));
 sky130_fd_sc_hd__and2_2 _25413_ (.A(_02585_),
    .B(\decoded_imm_uj[7] ),
    .X(_04330_));
 sky130_fd_sc_hd__a21oi_2 _25414_ (.A1(_04326_),
    .A2(_04329_),
    .B1(_04330_),
    .Y(_04331_));
 sky130_fd_sc_hd__xor2_2 _25415_ (.A(_04328_),
    .B(_04331_),
    .X(_01588_));
 sky130_fd_sc_hd__buf_1 _25416_ (.A(_02587_),
    .X(_04332_));
 sky130_fd_sc_hd__and4_2 _25417_ (.A(_04316_),
    .B(_17564_),
    .C(_04322_),
    .D(_17572_),
    .X(_04333_));
 sky130_fd_sc_hd__xor2_2 _25418_ (.A(_04332_),
    .B(_04333_),
    .X(_01591_));
 sky130_fd_sc_hd__xor2_2 _25419_ (.A(_04332_),
    .B(\decoded_imm_uj[9] ),
    .X(_04334_));
 sky130_fd_sc_hd__nor2_2 _25420_ (.A(_17563_),
    .B(_18930_),
    .Y(_04335_));
 sky130_fd_sc_hd__and2_2 _25421_ (.A(_02586_),
    .B(\decoded_imm_uj[8] ),
    .X(_04336_));
 sky130_fd_sc_hd__o21bai_2 _25422_ (.A1(_04335_),
    .A2(_04331_),
    .B1_N(_04336_),
    .Y(_04337_));
 sky130_fd_sc_hd__xor2_2 _25423_ (.A(_04334_),
    .B(_04337_),
    .X(_01592_));
 sky130_fd_sc_hd__and4_2 _25424_ (.A(_04323_),
    .B(_04332_),
    .C(_17563_),
    .D(_04322_),
    .X(_04338_));
 sky130_fd_sc_hd__xor2_2 _25425_ (.A(_17555_),
    .B(_04338_),
    .X(_01595_));
 sky130_fd_sc_hd__xnor2_2 _25426_ (.A(_17555_),
    .B(_18929_),
    .Y(_04339_));
 sky130_fd_sc_hd__nand2_2 _25427_ (.A(_17560_),
    .B(_19423_),
    .Y(_04340_));
 sky130_fd_sc_hd__and2_2 _25428_ (.A(_02587_),
    .B(\decoded_imm_uj[9] ),
    .X(_04341_));
 sky130_fd_sc_hd__a21oi_2 _25429_ (.A1(_04337_),
    .A2(_04340_),
    .B1(_04341_),
    .Y(_04342_));
 sky130_fd_sc_hd__xor2_2 _25430_ (.A(_04339_),
    .B(_04342_),
    .X(_01596_));
 sky130_fd_sc_hd__and4_2 _25431_ (.A(_04327_),
    .B(_17554_),
    .C(_02587_),
    .D(_17563_),
    .X(_04343_));
 sky130_fd_sc_hd__xor2_2 _25432_ (.A(_17550_),
    .B(_04343_),
    .X(_01599_));
 sky130_fd_sc_hd__xor2_2 _25433_ (.A(_02589_),
    .B(\decoded_imm_uj[11] ),
    .X(_04344_));
 sky130_fd_sc_hd__nor2_2 _25434_ (.A(_17554_),
    .B(_18929_),
    .Y(_04345_));
 sky130_fd_sc_hd__and2_2 _25435_ (.A(_02588_),
    .B(\decoded_imm_uj[10] ),
    .X(_04346_));
 sky130_fd_sc_hd__o21bai_2 _25436_ (.A1(_04345_),
    .A2(_04342_),
    .B1_N(_04346_),
    .Y(_04347_));
 sky130_fd_sc_hd__xor2_2 _25437_ (.A(_04344_),
    .B(_04347_),
    .X(_01600_));
 sky130_fd_sc_hd__and4_2 _25438_ (.A(_04333_),
    .B(_17550_),
    .C(_17555_),
    .D(_04332_),
    .X(_04348_));
 sky130_fd_sc_hd__xor2_2 _25439_ (.A(_17544_),
    .B(_04348_),
    .X(_01603_));
 sky130_fd_sc_hd__xnor2_2 _25440_ (.A(_02561_),
    .B(\decoded_imm_uj[12] ),
    .Y(_04349_));
 sky130_fd_sc_hd__and2_2 _25441_ (.A(_02589_),
    .B(\decoded_imm_uj[11] ),
    .X(_04350_));
 sky130_fd_sc_hd__a21oi_2 _25442_ (.A1(_04347_),
    .A2(_04344_),
    .B1(_04350_),
    .Y(_04351_));
 sky130_fd_sc_hd__xor2_2 _25443_ (.A(_04349_),
    .B(_04351_),
    .X(_01604_));
 sky130_fd_sc_hd__and4_2 _25444_ (.A(_04338_),
    .B(_17544_),
    .C(_02589_),
    .D(_17554_),
    .X(_04352_));
 sky130_fd_sc_hd__xor2_2 _25445_ (.A(_17541_),
    .B(_04352_),
    .X(_01607_));
 sky130_fd_sc_hd__xor2_2 _25446_ (.A(_02562_),
    .B(\decoded_imm_uj[13] ),
    .X(_04353_));
 sky130_fd_sc_hd__and2_2 _25447_ (.A(_02561_),
    .B(\decoded_imm_uj[12] ),
    .X(_04354_));
 sky130_fd_sc_hd__o21bai_2 _25448_ (.A1(_04349_),
    .A2(_04351_),
    .B1_N(_04354_),
    .Y(_04355_));
 sky130_fd_sc_hd__xor2_2 _25449_ (.A(_04353_),
    .B(_04355_),
    .X(_01608_));
 sky130_fd_sc_hd__and4_2 _25450_ (.A(_04343_),
    .B(_02562_),
    .C(_02561_),
    .D(_17550_),
    .X(_04356_));
 sky130_fd_sc_hd__xor2_2 _25451_ (.A(_17534_),
    .B(_04356_),
    .X(_01611_));
 sky130_fd_sc_hd__xnor2_2 _25452_ (.A(_02563_),
    .B(\decoded_imm_uj[14] ),
    .Y(_04357_));
 sky130_fd_sc_hd__and2_2 _25453_ (.A(_02562_),
    .B(\decoded_imm_uj[13] ),
    .X(_04358_));
 sky130_fd_sc_hd__a21oi_2 _25454_ (.A1(_04355_),
    .A2(_04353_),
    .B1(_04358_),
    .Y(_04359_));
 sky130_fd_sc_hd__xor2_2 _25455_ (.A(_04357_),
    .B(_04359_),
    .X(_01612_));
 sky130_fd_sc_hd__and4_2 _25456_ (.A(_04348_),
    .B(_17534_),
    .C(_17541_),
    .D(_17544_),
    .X(_04360_));
 sky130_fd_sc_hd__xor2_2 _25457_ (.A(_17531_),
    .B(_04360_),
    .X(_01615_));
 sky130_fd_sc_hd__xor2_2 _25458_ (.A(_02564_),
    .B(\decoded_imm_uj[15] ),
    .X(_04361_));
 sky130_fd_sc_hd__and2_2 _25459_ (.A(_02563_),
    .B(\decoded_imm_uj[14] ),
    .X(_04362_));
 sky130_fd_sc_hd__o21bai_2 _25460_ (.A1(_04357_),
    .A2(_04359_),
    .B1_N(_04362_),
    .Y(_04363_));
 sky130_fd_sc_hd__xor2_2 _25461_ (.A(_04361_),
    .B(_04363_),
    .X(_01616_));
 sky130_fd_sc_hd__and4_2 _25462_ (.A(_04352_),
    .B(_17531_),
    .C(_02563_),
    .D(_17541_),
    .X(_04364_));
 sky130_fd_sc_hd__xor2_2 _25463_ (.A(_17527_),
    .B(_04364_),
    .X(_01619_));
 sky130_fd_sc_hd__xnor2_2 _25464_ (.A(_02565_),
    .B(\decoded_imm_uj[16] ),
    .Y(_04365_));
 sky130_fd_sc_hd__and2_2 _25465_ (.A(_02564_),
    .B(\decoded_imm_uj[15] ),
    .X(_04366_));
 sky130_fd_sc_hd__a21oi_2 _25466_ (.A1(_04363_),
    .A2(_04361_),
    .B1(_04366_),
    .Y(_04367_));
 sky130_fd_sc_hd__xor2_2 _25467_ (.A(_04365_),
    .B(_04367_),
    .X(_01620_));
 sky130_fd_sc_hd__and4_2 _25468_ (.A(_04356_),
    .B(_02565_),
    .C(_02564_),
    .D(_17534_),
    .X(_04368_));
 sky130_fd_sc_hd__xor2_2 _25469_ (.A(_17520_),
    .B(_04368_),
    .X(_01623_));
 sky130_fd_sc_hd__xor2_2 _25470_ (.A(_02566_),
    .B(\decoded_imm_uj[17] ),
    .X(_04369_));
 sky130_fd_sc_hd__and2_2 _25471_ (.A(_02565_),
    .B(\decoded_imm_uj[16] ),
    .X(_04370_));
 sky130_fd_sc_hd__o21bai_2 _25472_ (.A1(_04365_),
    .A2(_04367_),
    .B1_N(_04370_),
    .Y(_04371_));
 sky130_fd_sc_hd__xor2_2 _25473_ (.A(_04369_),
    .B(_04371_),
    .X(_01624_));
 sky130_fd_sc_hd__and4_2 _25474_ (.A(_04360_),
    .B(_17520_),
    .C(_17527_),
    .D(_17531_),
    .X(_04372_));
 sky130_fd_sc_hd__xor2_2 _25475_ (.A(_17518_),
    .B(_04372_),
    .X(_01627_));
 sky130_fd_sc_hd__xnor2_2 _25476_ (.A(_17518_),
    .B(_18926_),
    .Y(_04373_));
 sky130_fd_sc_hd__and2_2 _25477_ (.A(_02566_),
    .B(\decoded_imm_uj[17] ),
    .X(_04374_));
 sky130_fd_sc_hd__a21oi_2 _25478_ (.A1(_04371_),
    .A2(_04369_),
    .B1(_04374_),
    .Y(_04375_));
 sky130_fd_sc_hd__xor2_2 _25479_ (.A(_04373_),
    .B(_04375_),
    .X(_01628_));
 sky130_fd_sc_hd__and4_2 _25480_ (.A(_04364_),
    .B(_17517_),
    .C(_02566_),
    .D(_17527_),
    .X(_04376_));
 sky130_fd_sc_hd__xor2_2 _25481_ (.A(_17511_),
    .B(_04376_),
    .X(_01631_));
 sky130_fd_sc_hd__xor2_2 _25482_ (.A(_02568_),
    .B(\decoded_imm_uj[19] ),
    .X(_04377_));
 sky130_fd_sc_hd__nor2_2 _25483_ (.A(_17517_),
    .B(_18926_),
    .Y(_04378_));
 sky130_fd_sc_hd__and2_2 _25484_ (.A(_02567_),
    .B(\decoded_imm_uj[18] ),
    .X(_04379_));
 sky130_fd_sc_hd__o21bai_2 _25485_ (.A1(_04378_),
    .A2(_04375_),
    .B1_N(_04379_),
    .Y(_04380_));
 sky130_fd_sc_hd__xor2_2 _25486_ (.A(_04377_),
    .B(_04380_),
    .X(_01632_));
 sky130_fd_sc_hd__and4_2 _25487_ (.A(_04368_),
    .B(_02568_),
    .C(_17517_),
    .D(_17520_),
    .X(_04381_));
 sky130_fd_sc_hd__xor2_2 _25488_ (.A(_17506_),
    .B(_04381_),
    .X(_01635_));
 sky130_fd_sc_hd__xnor2_2 _25489_ (.A(_17506_),
    .B(_18924_),
    .Y(_04382_));
 sky130_fd_sc_hd__and2_2 _25490_ (.A(_02568_),
    .B(\decoded_imm_uj[19] ),
    .X(_04383_));
 sky130_fd_sc_hd__a21oi_2 _25491_ (.A1(_04380_),
    .A2(_04377_),
    .B1(_04383_),
    .Y(_04384_));
 sky130_fd_sc_hd__xor2_2 _25492_ (.A(_04382_),
    .B(_04384_),
    .X(_01636_));
 sky130_fd_sc_hd__and4_2 _25493_ (.A(_04372_),
    .B(_17506_),
    .C(_17511_),
    .D(_17518_),
    .X(_04385_));
 sky130_fd_sc_hd__xor2_2 _25494_ (.A(_17501_),
    .B(_04385_),
    .X(_01639_));
 sky130_fd_sc_hd__xor2_2 _25495_ (.A(_02570_),
    .B(\decoded_imm_uj[20] ),
    .X(_04386_));
 sky130_fd_sc_hd__nor2_2 _25496_ (.A(_17505_),
    .B(\decoded_imm_uj[20] ),
    .Y(_04387_));
 sky130_fd_sc_hd__and2_2 _25497_ (.A(_02569_),
    .B(\decoded_imm_uj[20] ),
    .X(_04388_));
 sky130_fd_sc_hd__o21bai_2 _25498_ (.A1(_04387_),
    .A2(_04384_),
    .B1_N(_04388_),
    .Y(_04389_));
 sky130_fd_sc_hd__xor2_2 _25499_ (.A(_04386_),
    .B(_04389_),
    .X(_01640_));
 sky130_fd_sc_hd__and4_2 _25500_ (.A(_04376_),
    .B(_17500_),
    .C(_17505_),
    .D(_17511_),
    .X(_04390_));
 sky130_fd_sc_hd__xor2_2 _25501_ (.A(_17497_),
    .B(_04390_),
    .X(_01643_));
 sky130_fd_sc_hd__xor2_2 _25502_ (.A(_02572_),
    .B(_18919_),
    .X(_04391_));
 sky130_fd_sc_hd__and2_2 _25503_ (.A(_17501_),
    .B(_19514_),
    .X(_04392_));
 sky130_fd_sc_hd__a21oi_2 _25504_ (.A1(_04389_),
    .A2(_04386_),
    .B1(_04392_),
    .Y(_04393_));
 sky130_fd_sc_hd__xnor2_2 _25505_ (.A(_04391_),
    .B(_04393_),
    .Y(_01644_));
 sky130_fd_sc_hd__and4_2 _25506_ (.A(_04381_),
    .B(_02572_),
    .C(_17500_),
    .D(_17505_),
    .X(_04394_));
 sky130_fd_sc_hd__xor2_2 _25507_ (.A(_17494_),
    .B(_04394_),
    .X(_01647_));
 sky130_fd_sc_hd__nand3_2 _25508_ (.A(_04389_),
    .B(_04386_),
    .C(_04391_),
    .Y(_04395_));
 sky130_fd_sc_hd__o21ai_2 _25509_ (.A1(_02572_),
    .A2(_17500_),
    .B1(_18920_),
    .Y(_04396_));
 sky130_fd_sc_hd__xor2_2 _25510_ (.A(_02573_),
    .B(_18919_),
    .X(_04397_));
 sky130_fd_sc_hd__a21boi_2 _25511_ (.A1(_04395_),
    .A2(_04396_),
    .B1_N(_04397_),
    .Y(_04398_));
 sky130_fd_sc_hd__and3b_2 _25512_ (.A_N(_04397_),
    .B(_04395_),
    .C(_04396_),
    .X(_04399_));
 sky130_fd_sc_hd__nor2_2 _25513_ (.A(_04398_),
    .B(_04399_),
    .Y(_01648_));
 sky130_fd_sc_hd__and4_2 _25514_ (.A(_04385_),
    .B(_17494_),
    .C(_17497_),
    .D(_17501_),
    .X(_04400_));
 sky130_fd_sc_hd__xor2_2 _25515_ (.A(_17490_),
    .B(_04400_),
    .X(_01651_));
 sky130_fd_sc_hd__xor2_2 _25516_ (.A(_02574_),
    .B(_18919_),
    .X(_04401_));
 sky130_fd_sc_hd__a21oi_2 _25517_ (.A1(_17494_),
    .A2(_18924_),
    .B1(_04398_),
    .Y(_04402_));
 sky130_fd_sc_hd__xnor2_2 _25518_ (.A(_04401_),
    .B(_04402_),
    .Y(_01652_));
 sky130_fd_sc_hd__and4_2 _25519_ (.A(_04390_),
    .B(_17490_),
    .C(_17493_),
    .D(_17497_),
    .X(_04403_));
 sky130_fd_sc_hd__xor2_2 _25520_ (.A(_17487_),
    .B(_04403_),
    .X(_01655_));
 sky130_fd_sc_hd__xor2_2 _25521_ (.A(_02575_),
    .B(_18920_),
    .X(_04404_));
 sky130_fd_sc_hd__nand2_2 _25522_ (.A(_04397_),
    .B(_04401_),
    .Y(_04405_));
 sky130_fd_sc_hd__o21ai_2 _25523_ (.A1(_02574_),
    .A2(_17493_),
    .B1(_18920_),
    .Y(_04406_));
 sky130_fd_sc_hd__o211ai_2 _25524_ (.A1(_04405_),
    .A2(_04395_),
    .B1(_04396_),
    .C1(_04406_),
    .Y(_04407_));
 sky130_fd_sc_hd__xor2_2 _25525_ (.A(_04404_),
    .B(_04407_),
    .X(_01656_));
 sky130_fd_sc_hd__and4_2 _25526_ (.A(_04394_),
    .B(_17486_),
    .C(_02574_),
    .D(_17493_),
    .X(_04408_));
 sky130_fd_sc_hd__xor2_2 _25527_ (.A(_17478_),
    .B(_04408_),
    .X(_01659_));
 sky130_fd_sc_hd__xor2_2 _25528_ (.A(_02576_),
    .B(_18921_),
    .X(_04409_));
 sky130_fd_sc_hd__and2_2 _25529_ (.A(_17487_),
    .B(_19514_),
    .X(_04410_));
 sky130_fd_sc_hd__a21oi_2 _25530_ (.A1(_04407_),
    .A2(_04404_),
    .B1(_04410_),
    .Y(_04411_));
 sky130_fd_sc_hd__xnor2_2 _25531_ (.A(_04409_),
    .B(_04411_),
    .Y(_01660_));
 sky130_fd_sc_hd__and4_2 _25532_ (.A(_04400_),
    .B(_17478_),
    .C(_17487_),
    .D(_17490_),
    .X(_04412_));
 sky130_fd_sc_hd__xor2_2 _25533_ (.A(_17475_),
    .B(_04412_),
    .X(_01663_));
 sky130_fd_sc_hd__nand3_2 _25534_ (.A(_04407_),
    .B(_04404_),
    .C(_04409_),
    .Y(_04413_));
 sky130_fd_sc_hd__o21ai_2 _25535_ (.A1(_02576_),
    .A2(_17486_),
    .B1(_18922_),
    .Y(_04414_));
 sky130_fd_sc_hd__xor2_2 _25536_ (.A(_02577_),
    .B(_18921_),
    .X(_04415_));
 sky130_fd_sc_hd__a21boi_2 _25537_ (.A1(_04413_),
    .A2(_04414_),
    .B1_N(_04415_),
    .Y(_04416_));
 sky130_fd_sc_hd__and3b_2 _25538_ (.A_N(_04415_),
    .B(_04413_),
    .C(_04414_),
    .X(_04417_));
 sky130_fd_sc_hd__nor2_2 _25539_ (.A(_04416_),
    .B(_04417_),
    .Y(_01664_));
 sky130_fd_sc_hd__and4_2 _25540_ (.A(_04403_),
    .B(_17475_),
    .C(_02576_),
    .D(_17486_),
    .X(_04418_));
 sky130_fd_sc_hd__xor2_2 _25541_ (.A(_17472_),
    .B(_04418_),
    .X(_01667_));
 sky130_fd_sc_hd__xor2_2 _25542_ (.A(_02578_),
    .B(_18921_),
    .X(_04419_));
 sky130_fd_sc_hd__a21oi_2 _25543_ (.A1(_17475_),
    .A2(_18924_),
    .B1(_04416_),
    .Y(_04420_));
 sky130_fd_sc_hd__xnor2_2 _25544_ (.A(_04419_),
    .B(_04420_),
    .Y(_01668_));
 sky130_fd_sc_hd__and4_2 _25545_ (.A(_04408_),
    .B(_17472_),
    .C(_02577_),
    .D(_17478_),
    .X(_04421_));
 sky130_fd_sc_hd__xor2_2 _25546_ (.A(_17469_),
    .B(_04421_),
    .X(_01671_));
 sky130_fd_sc_hd__xor2_2 _25547_ (.A(_02579_),
    .B(_18922_),
    .X(_04422_));
 sky130_fd_sc_hd__nand2_2 _25548_ (.A(_04415_),
    .B(_04419_),
    .Y(_04423_));
 sky130_fd_sc_hd__o21ai_2 _25549_ (.A1(_02578_),
    .A2(_02577_),
    .B1(_18923_),
    .Y(_04424_));
 sky130_fd_sc_hd__o211ai_2 _25550_ (.A1(_04423_),
    .A2(_04413_),
    .B1(_04414_),
    .C1(_04424_),
    .Y(_04425_));
 sky130_fd_sc_hd__xor2_2 _25551_ (.A(_04422_),
    .B(_04425_),
    .X(_01672_));
 sky130_fd_sc_hd__nand3_2 _25552_ (.A(_04418_),
    .B(_17469_),
    .C(_17472_),
    .Y(_04426_));
 sky130_fd_sc_hd__xor2_2 _25553_ (.A(_17464_),
    .B(_04426_),
    .X(_01675_));
 sky130_fd_sc_hd__buf_1 _25554_ (.A(_18923_),
    .X(_04427_));
 sky130_fd_sc_hd__xnor2_2 _25555_ (.A(_17463_),
    .B(_04427_),
    .Y(_04428_));
 sky130_fd_sc_hd__and2_2 _25556_ (.A(_02579_),
    .B(_04427_),
    .X(_04429_));
 sky130_fd_sc_hd__a21oi_2 _25557_ (.A1(_04425_),
    .A2(_04422_),
    .B1(_04429_),
    .Y(_04430_));
 sky130_fd_sc_hd__xor2_2 _25558_ (.A(_04428_),
    .B(_04430_),
    .X(_01676_));
 sky130_fd_sc_hd__nand3_2 _25559_ (.A(_04421_),
    .B(_17463_),
    .C(_17469_),
    .Y(_04431_));
 sky130_fd_sc_hd__xor2_2 _25560_ (.A(_17460_),
    .B(_04431_),
    .X(_01679_));
 sky130_fd_sc_hd__o211ai_2 _25561_ (.A1(_02580_),
    .A2(_04427_),
    .B1(_04422_),
    .C1(_04425_),
    .Y(_04432_));
 sky130_fd_sc_hd__o21ai_2 _25562_ (.A1(_17463_),
    .A2(_02579_),
    .B1(_04427_),
    .Y(_04433_));
 sky130_fd_sc_hd__xnor2_2 _25563_ (.A(_02581_),
    .B(_19514_),
    .Y(_04434_));
 sky130_fd_sc_hd__a21oi_2 _25564_ (.A1(_04432_),
    .A2(_04433_),
    .B1(_04434_),
    .Y(_04435_));
 sky130_fd_sc_hd__and3_2 _25565_ (.A(_04432_),
    .B(_04433_),
    .C(_04434_),
    .X(_04436_));
 sky130_fd_sc_hd__nor2_2 _25566_ (.A(_04435_),
    .B(_04436_),
    .Y(_01680_));
 sky130_fd_sc_hd__nor2_2 _25567_ (.A(_19667_),
    .B(\mem_wordsize[1] ),
    .Y(_01683_));
 sky130_fd_sc_hd__buf_1 _25568_ (.A(_19667_),
    .X(_04437_));
 sky130_fd_sc_hd__mux2_2 _25569_ (.A0(_04076_),
    .A1(_19117_),
    .S(_04437_),
    .X(_04438_));
 sky130_vsdinv _25570_ (.A(_00304_),
    .Y(_04439_));
 sky130_fd_sc_hd__a21boi_2 _25571_ (.A1(_04438_),
    .A2(_04439_),
    .B1_N(mem_la_write),
    .Y(_01684_));
 sky130_fd_sc_hd__buf_1 _25572_ (.A(_19763_),
    .X(_04440_));
 sky130_fd_sc_hd__nand3_2 _25573_ (.A(_00301_),
    .B(_04440_),
    .C(_01685_),
    .Y(_04441_));
 sky130_vsdinv _25574_ (.A(_04441_),
    .Y(_01686_));
 sky130_vsdinv _25575_ (.A(_19116_),
    .Y(_04442_));
 sky130_fd_sc_hd__nand2_2 _25576_ (.A(_04442_),
    .B(_19775_),
    .Y(_04443_));
 sky130_fd_sc_hd__buf_1 _25577_ (.A(_04443_),
    .X(_04444_));
 sky130_fd_sc_hd__a21boi_2 _25578_ (.A1(_04438_),
    .A2(_04444_),
    .B1_N(mem_la_write),
    .Y(_01687_));
 sky130_fd_sc_hd__nand3_2 _25579_ (.A(_00301_),
    .B(_04440_),
    .C(_01688_),
    .Y(_04445_));
 sky130_vsdinv _25580_ (.A(_04445_),
    .Y(_01689_));
 sky130_fd_sc_hd__buf_1 _25581_ (.A(_19116_),
    .X(_04446_));
 sky130_fd_sc_hd__a21oi_2 _25582_ (.A1(_04446_),
    .A2(_04437_),
    .B1(_01683_),
    .Y(_04447_));
 sky130_fd_sc_hd__o21ai_2 _25583_ (.A1(_04442_),
    .A2(_19543_),
    .B1(_04447_),
    .Y(mem_la_wstrb[2]));
 sky130_fd_sc_hd__and2_2 _25584_ (.A(mem_la_wstrb[2]),
    .B(mem_la_write),
    .X(_01690_));
 sky130_fd_sc_hd__nand3_2 _25585_ (.A(_00301_),
    .B(_04440_),
    .C(_01691_),
    .Y(_04448_));
 sky130_vsdinv _25586_ (.A(_04448_),
    .Y(_01692_));
 sky130_fd_sc_hd__o21ai_2 _25587_ (.A1(_04442_),
    .A2(_19567_),
    .B1(_04447_),
    .Y(mem_la_wstrb[3]));
 sky130_fd_sc_hd__and2_2 _25588_ (.A(mem_la_wstrb[3]),
    .B(_19677_),
    .X(_01693_));
 sky130_fd_sc_hd__nand3_2 _25589_ (.A(_16847_),
    .B(_19763_),
    .C(_01694_),
    .Y(_04449_));
 sky130_vsdinv _25590_ (.A(_04449_),
    .Y(_01695_));
 sky130_fd_sc_hd__nor2_2 _25591_ (.A(_17994_),
    .B(irq[1]),
    .Y(_01696_));
 sky130_vsdinv _25592_ (.A(_01696_),
    .Y(_01697_));
 sky130_fd_sc_hd__o21a_2 _25593_ (.A1(_17994_),
    .A2(irq[1]),
    .B1(_17210_),
    .X(_01698_));
 sky130_fd_sc_hd__buf_1 _25594_ (.A(_17018_),
    .X(_04450_));
 sky130_fd_sc_hd__nand3b_2 _25595_ (.A_N(_02542_),
    .B(_17075_),
    .C(_00297_),
    .Y(_04451_));
 sky130_fd_sc_hd__nor2_2 _25596_ (.A(_04450_),
    .B(_04451_),
    .Y(_01700_));
 sky130_fd_sc_hd__o21a_2 _25597_ (.A1(_19548_),
    .A2(_17210_),
    .B1(_01696_),
    .X(_01701_));
 sky130_fd_sc_hd__and2b_2 _25598_ (.A_N(_01704_),
    .B(_18003_),
    .X(_04452_));
 sky130_fd_sc_hd__a21o_2 _25599_ (.A1(_04451_),
    .A2(_01697_),
    .B1(_04452_),
    .X(_01705_));
 sky130_vsdinv _25600_ (.A(_17029_),
    .Y(_01706_));
 sky130_vsdinv _25601_ (.A(mem_rdata[0]),
    .Y(_01707_));
 sky130_vsdinv _25602_ (.A(mem_rdata[8]),
    .Y(_01812_));
 sky130_fd_sc_hd__buf_1 _25603_ (.A(_19117_),
    .X(_04453_));
 sky130_fd_sc_hd__buf_1 _25604_ (.A(_19543_),
    .X(_04454_));
 sky130_fd_sc_hd__nand3_2 _25605_ (.A(_04453_),
    .B(_04454_),
    .C(mem_rdata[24]),
    .Y(_04455_));
 sky130_fd_sc_hd__nand3b_2 _25606_ (.A_N(_19123_),
    .B(_19118_),
    .C(mem_rdata[16]),
    .Y(_04456_));
 sky130_fd_sc_hd__o211a_2 _25607_ (.A1(_01812_),
    .A2(_04444_),
    .B1(_04455_),
    .C1(_04456_),
    .X(_01708_));
 sky130_vsdinv _25608_ (.A(_04076_),
    .Y(_04457_));
 sky130_fd_sc_hd__buf_1 _25609_ (.A(_04457_),
    .X(_04458_));
 sky130_fd_sc_hd__o2bb2a_2 _25610_ (.A1_N(_19758_),
    .A2_N(_01710_),
    .B1(_01709_),
    .B2(_04458_),
    .X(_01711_));
 sky130_fd_sc_hd__buf_1 _25611_ (.A(instr_rdinstr),
    .X(_04459_));
 sky130_fd_sc_hd__buf_1 _25612_ (.A(_04459_),
    .X(_04460_));
 sky130_fd_sc_hd__and2_2 _25613_ (.A(\count_instr[32] ),
    .B(_18987_),
    .X(_04461_));
 sky130_fd_sc_hd__a221oi_2 _25614_ (.A1(_17814_),
    .A2(_04460_),
    .B1(_18997_),
    .B2(_18058_),
    .C1(_04461_),
    .Y(_01715_));
 sky130_fd_sc_hd__buf_1 _25615_ (.A(instr_maskirq),
    .X(_04462_));
 sky130_fd_sc_hd__buf_1 _25616_ (.A(_04462_),
    .X(_04463_));
 sky130_fd_sc_hd__buf_1 _25617_ (.A(_18952_),
    .X(_04464_));
 sky130_fd_sc_hd__nor3b_2 _25618_ (.A(_17005_),
    .B(_17105_),
    .C_N(_00370_),
    .Y(_04465_));
 sky130_fd_sc_hd__a221oi_2 _25619_ (.A1(_17214_),
    .A2(_04463_),
    .B1(_04464_),
    .B2(_04102_),
    .C1(_04465_),
    .Y(_01718_));
 sky130_fd_sc_hd__and2_2 _25620_ (.A(_18941_),
    .B(\reg_next_pc[0] ),
    .X(_04466_));
 sky130_fd_sc_hd__buf_1 _25621_ (.A(_19678_),
    .X(_04467_));
 sky130_fd_sc_hd__o21ai_2 _25622_ (.A1(_18941_),
    .A2(_19382_),
    .B1(_04467_),
    .Y(_04468_));
 sky130_fd_sc_hd__buf_1 _25623_ (.A(_17021_),
    .X(_04469_));
 sky130_fd_sc_hd__buf_1 _25624_ (.A(_04469_),
    .X(_04470_));
 sky130_fd_sc_hd__a2bb2oi_2 _25625_ (.A1_N(_01719_),
    .A2_N(_04470_),
    .B1(_19774_),
    .B2(_01713_),
    .Y(_04471_));
 sky130_fd_sc_hd__o221ai_2 _25626_ (.A1(_18028_),
    .A2(_01712_),
    .B1(_04466_),
    .B2(_04468_),
    .C1(_04471_),
    .Y(_01720_));
 sky130_vsdinv _25627_ (.A(mem_rdata[1]),
    .Y(_01721_));
 sky130_vsdinv _25628_ (.A(mem_rdata[9]),
    .Y(_01826_));
 sky130_fd_sc_hd__nand3_2 _25629_ (.A(_04453_),
    .B(_04454_),
    .C(mem_rdata[25]),
    .Y(_04472_));
 sky130_fd_sc_hd__nand3b_2 _25630_ (.A_N(_19123_),
    .B(_19118_),
    .C(mem_rdata[17]),
    .Y(_04473_));
 sky130_fd_sc_hd__o211a_2 _25631_ (.A1(_01826_),
    .A2(_04444_),
    .B1(_04472_),
    .C1(_04473_),
    .X(_01722_));
 sky130_fd_sc_hd__o2bb2a_2 _25632_ (.A1_N(_19758_),
    .A2_N(_01724_),
    .B1(_01723_),
    .B2(_04458_),
    .X(_01725_));
 sky130_vsdinv _25633_ (.A(_18267_),
    .Y(_01728_));
 sky130_fd_sc_hd__buf_1 _25634_ (.A(_04459_),
    .X(_04474_));
 sky130_fd_sc_hd__and2_2 _25635_ (.A(\count_instr[33] ),
    .B(_18987_),
    .X(_04475_));
 sky130_fd_sc_hd__a221oi_2 _25636_ (.A1(_17848_),
    .A2(_04474_),
    .B1(_18997_),
    .B2(_18182_),
    .C1(_04475_),
    .Y(_01729_));
 sky130_fd_sc_hd__nand2_2 _25637_ (.A(_17005_),
    .B(_17007_),
    .Y(_04476_));
 sky130_fd_sc_hd__buf_1 _25638_ (.A(_04476_),
    .X(_04477_));
 sky130_fd_sc_hd__buf_1 _25639_ (.A(_04477_),
    .X(_04478_));
 sky130_fd_sc_hd__buf_1 _25640_ (.A(instr_maskirq),
    .X(_04479_));
 sky130_fd_sc_hd__buf_1 _25641_ (.A(_04479_),
    .X(_04480_));
 sky130_fd_sc_hd__and2_2 _25642_ (.A(_17209_),
    .B(_04480_),
    .X(_04481_));
 sky130_fd_sc_hd__a221oi_2 _25643_ (.A1(_18953_),
    .A2(_04103_),
    .B1(\cpuregs_rs1[1] ),
    .B2(_04478_),
    .C1(_04481_),
    .Y(_01731_));
 sky130_fd_sc_hd__buf_1 _25644_ (.A(_16984_),
    .X(_04482_));
 sky130_fd_sc_hd__xor2_2 _25645_ (.A(\reg_pc[1] ),
    .B(_19397_),
    .X(_04483_));
 sky130_fd_sc_hd__nor2_2 _25646_ (.A(_04466_),
    .B(_04483_),
    .Y(_04484_));
 sky130_fd_sc_hd__and2_2 _25647_ (.A(_04483_),
    .B(_04466_),
    .X(_04485_));
 sky130_fd_sc_hd__or2b_2 _25648_ (.A(_01726_),
    .B_N(_17390_),
    .X(_04486_));
 sky130_fd_sc_hd__buf_1 _25649_ (.A(_18540_),
    .X(_04487_));
 sky130_fd_sc_hd__buf_1 _25650_ (.A(_19625_),
    .X(_04488_));
 sky130_fd_sc_hd__a2bb2oi_2 _25651_ (.A1_N(_01732_),
    .A2_N(_04487_),
    .B1(_04488_),
    .B2(_01727_),
    .Y(_04489_));
 sky130_fd_sc_hd__o311ai_2 _25652_ (.A1(_04482_),
    .A2(_04484_),
    .A3(_04485_),
    .B1(_04486_),
    .C1(_04489_),
    .Y(_01733_));
 sky130_vsdinv _25653_ (.A(mem_rdata[2]),
    .Y(_01734_));
 sky130_vsdinv _25654_ (.A(mem_rdata[10]),
    .Y(_01839_));
 sky130_fd_sc_hd__buf_1 _25655_ (.A(_04443_),
    .X(_04490_));
 sky130_fd_sc_hd__buf_1 _25656_ (.A(_04446_),
    .X(_04491_));
 sky130_fd_sc_hd__buf_1 _25657_ (.A(_04491_),
    .X(_04492_));
 sky130_fd_sc_hd__nand3_2 _25658_ (.A(_04492_),
    .B(_04454_),
    .C(mem_rdata[26]),
    .Y(_04493_));
 sky130_fd_sc_hd__buf_1 _25659_ (.A(_04491_),
    .X(_04494_));
 sky130_fd_sc_hd__nand3b_2 _25660_ (.A_N(_19123_),
    .B(_04494_),
    .C(mem_rdata[18]),
    .Y(_04495_));
 sky130_fd_sc_hd__o211a_2 _25661_ (.A1(_01839_),
    .A2(_04490_),
    .B1(_04493_),
    .C1(_04495_),
    .X(_01735_));
 sky130_fd_sc_hd__o2bb2a_2 _25662_ (.A1_N(_19758_),
    .A2_N(_01737_),
    .B1(_01736_),
    .B2(_04458_),
    .X(_01738_));
 sky130_vsdinv _25663_ (.A(_18264_),
    .Y(_01741_));
 sky130_fd_sc_hd__and2_2 _25664_ (.A(_18996_),
    .B(_18099_),
    .X(_04496_));
 sky130_fd_sc_hd__a221oi_2 _25665_ (.A1(\count_instr[34] ),
    .A2(_18988_),
    .B1(_17847_),
    .B2(_18991_),
    .C1(_04496_),
    .Y(_01742_));
 sky130_fd_sc_hd__and2_2 _25666_ (.A(_17990_),
    .B(_04480_),
    .X(_04497_));
 sky130_fd_sc_hd__a221oi_2 _25667_ (.A1(_18953_),
    .A2(_04104_),
    .B1(\cpuregs_rs1[2] ),
    .B2(_04478_),
    .C1(_04497_),
    .Y(_01744_));
 sky130_fd_sc_hd__nor2_2 _25668_ (.A(\reg_pc[2] ),
    .B(_19400_),
    .Y(_04498_));
 sky130_fd_sc_hd__and2_2 _25669_ (.A(\reg_pc[2] ),
    .B(_19400_),
    .X(_04499_));
 sky130_fd_sc_hd__nor2_2 _25670_ (.A(_04498_),
    .B(_04499_),
    .Y(_04500_));
 sky130_fd_sc_hd__and2_2 _25671_ (.A(\reg_pc[1] ),
    .B(_19397_),
    .X(_04501_));
 sky130_fd_sc_hd__a21o_2 _25672_ (.A1(_04483_),
    .A2(_04466_),
    .B1(_04501_),
    .X(_04502_));
 sky130_fd_sc_hd__o21bai_2 _25673_ (.A1(_04500_),
    .A2(_04502_),
    .B1_N(_16984_),
    .Y(_04503_));
 sky130_fd_sc_hd__and2_2 _25674_ (.A(_04502_),
    .B(_04500_),
    .X(_04504_));
 sky130_fd_sc_hd__a2bb2oi_2 _25675_ (.A1_N(_01745_),
    .A2_N(_04470_),
    .B1(_19774_),
    .B2(_01740_),
    .Y(_04505_));
 sky130_fd_sc_hd__o221ai_2 _25676_ (.A1(_18028_),
    .A2(_01739_),
    .B1(_04503_),
    .B2(_04504_),
    .C1(_04505_),
    .Y(_01746_));
 sky130_vsdinv _25677_ (.A(mem_rdata[3]),
    .Y(_01747_));
 sky130_vsdinv _25678_ (.A(mem_rdata[11]),
    .Y(_01852_));
 sky130_fd_sc_hd__nand3_2 _25679_ (.A(_04492_),
    .B(_04454_),
    .C(mem_rdata[27]),
    .Y(_04506_));
 sky130_fd_sc_hd__buf_1 _25680_ (.A(_19775_),
    .X(_04507_));
 sky130_fd_sc_hd__nand3b_2 _25681_ (.A_N(_04507_),
    .B(_04494_),
    .C(mem_rdata[19]),
    .Y(_04508_));
 sky130_fd_sc_hd__o211a_2 _25682_ (.A1(_01852_),
    .A2(_04490_),
    .B1(_04506_),
    .C1(_04508_),
    .X(_01748_));
 sky130_fd_sc_hd__buf_1 _25683_ (.A(_19757_),
    .X(_04509_));
 sky130_fd_sc_hd__o2bb2a_2 _25684_ (.A1_N(_04509_),
    .A2_N(_01750_),
    .B1(_01749_),
    .B2(_04458_),
    .X(_01751_));
 sky130_fd_sc_hd__buf_1 _25685_ (.A(instr_rdinstrh),
    .X(_04510_));
 sky130_fd_sc_hd__buf_1 _25686_ (.A(_04510_),
    .X(_04511_));
 sky130_fd_sc_hd__and2_2 _25687_ (.A(_17727_),
    .B(_04511_),
    .X(_04512_));
 sky130_fd_sc_hd__a221oi_2 _25688_ (.A1(\count_instr[3] ),
    .A2(_04474_),
    .B1(_18997_),
    .B2(_18180_),
    .C1(_04512_),
    .Y(_01755_));
 sky130_fd_sc_hd__buf_1 _25689_ (.A(_17022_),
    .X(_04513_));
 sky130_fd_sc_hd__buf_1 _25690_ (.A(_04513_),
    .X(_04514_));
 sky130_fd_sc_hd__and2_2 _25691_ (.A(_04514_),
    .B(\timer[3] ),
    .X(_04515_));
 sky130_fd_sc_hd__a221oi_2 _25692_ (.A1(_17205_),
    .A2(_04463_),
    .B1(\cpuregs_rs1[3] ),
    .B2(_04478_),
    .C1(_04515_),
    .Y(_01757_));
 sky130_fd_sc_hd__and2_2 _25693_ (.A(\reg_pc[3] ),
    .B(_19404_),
    .X(_04516_));
 sky130_fd_sc_hd__nor2_2 _25694_ (.A(_17584_),
    .B(_19404_),
    .Y(_04517_));
 sky130_vsdinv _25695_ (.A(_04498_),
    .Y(_04518_));
 sky130_fd_sc_hd__a21oi_2 _25696_ (.A1(_04502_),
    .A2(_04518_),
    .B1(_04499_),
    .Y(_04519_));
 sky130_fd_sc_hd__o21a_2 _25697_ (.A1(_04516_),
    .A2(_04517_),
    .B1(_04519_),
    .X(_04520_));
 sky130_fd_sc_hd__o31ai_2 _25698_ (.A1(_04516_),
    .A2(_04517_),
    .A3(_04519_),
    .B1(_04467_),
    .Y(_04521_));
 sky130_fd_sc_hd__buf_1 _25699_ (.A(_19625_),
    .X(_04522_));
 sky130_fd_sc_hd__a2bb2oi_2 _25700_ (.A1_N(_01758_),
    .A2_N(_04470_),
    .B1(_04522_),
    .B2(_01753_),
    .Y(_04523_));
 sky130_fd_sc_hd__o221ai_2 _25701_ (.A1(_18028_),
    .A2(_01752_),
    .B1(_04520_),
    .B2(_04521_),
    .C1(_04523_),
    .Y(_01759_));
 sky130_vsdinv _25702_ (.A(mem_rdata[4]),
    .Y(_01760_));
 sky130_vsdinv _25703_ (.A(mem_rdata[12]),
    .Y(_01865_));
 sky130_fd_sc_hd__buf_1 _25704_ (.A(_19775_),
    .X(_04524_));
 sky130_fd_sc_hd__nand3_2 _25705_ (.A(_04492_),
    .B(_04524_),
    .C(mem_rdata[28]),
    .Y(_04525_));
 sky130_fd_sc_hd__nand3b_2 _25706_ (.A_N(_04507_),
    .B(_04494_),
    .C(mem_rdata[20]),
    .Y(_04526_));
 sky130_fd_sc_hd__o211a_2 _25707_ (.A1(_01865_),
    .A2(_04490_),
    .B1(_04525_),
    .C1(_04526_),
    .X(_01761_));
 sky130_fd_sc_hd__buf_1 _25708_ (.A(_04457_),
    .X(_04527_));
 sky130_fd_sc_hd__o2bb2a_2 _25709_ (.A1_N(_04509_),
    .A2_N(_01763_),
    .B1(_01762_),
    .B2(_04527_),
    .X(_01764_));
 sky130_fd_sc_hd__buf_1 _25710_ (.A(instr_rdcycleh),
    .X(_04528_));
 sky130_fd_sc_hd__buf_1 _25711_ (.A(_04528_),
    .X(_04529_));
 sky130_fd_sc_hd__buf_1 _25712_ (.A(_04529_),
    .X(_04530_));
 sky130_fd_sc_hd__and2_2 _25713_ (.A(\count_instr[36] ),
    .B(_04511_),
    .X(_04531_));
 sky130_fd_sc_hd__a221oi_2 _25714_ (.A1(_17844_),
    .A2(_04474_),
    .B1(_04530_),
    .B2(_18170_),
    .C1(_04531_),
    .Y(_01768_));
 sky130_fd_sc_hd__and2_2 _25715_ (.A(_04514_),
    .B(\timer[4] ),
    .X(_04532_));
 sky130_fd_sc_hd__a221oi_2 _25716_ (.A1(_17202_),
    .A2(_04463_),
    .B1(\cpuregs_rs1[4] ),
    .B2(_04478_),
    .C1(_04532_),
    .Y(_01770_));
 sky130_fd_sc_hd__xor2_2 _25717_ (.A(\reg_pc[4] ),
    .B(\decoded_imm[4] ),
    .X(_04533_));
 sky130_fd_sc_hd__buf_1 _25718_ (.A(_04533_),
    .X(_04534_));
 sky130_fd_sc_hd__o21bai_2 _25719_ (.A1(_04517_),
    .A2(_04519_),
    .B1_N(_04516_),
    .Y(_04535_));
 sky130_fd_sc_hd__buf_1 _25720_ (.A(_04535_),
    .X(_04536_));
 sky130_fd_sc_hd__or2_2 _25721_ (.A(_04534_),
    .B(_04536_),
    .X(_04537_));
 sky130_fd_sc_hd__nand2_2 _25722_ (.A(_04536_),
    .B(_04534_),
    .Y(_04538_));
 sky130_fd_sc_hd__and2b_2 _25723_ (.A_N(_01765_),
    .B(_04073_),
    .X(_04539_));
 sky130_fd_sc_hd__buf_1 _25724_ (.A(_18540_),
    .X(_04540_));
 sky130_fd_sc_hd__o2bb2ai_2 _25725_ (.A1_N(_04450_),
    .A2_N(_01766_),
    .B1(_01771_),
    .B2(_04540_),
    .Y(_04541_));
 sky130_fd_sc_hd__a311o_2 _25726_ (.A1(_04537_),
    .A2(_04538_),
    .A3(_19679_),
    .B1(_04539_),
    .C1(_04541_),
    .X(_01772_));
 sky130_vsdinv _25727_ (.A(mem_rdata[5]),
    .Y(_01773_));
 sky130_vsdinv _25728_ (.A(mem_rdata[13]),
    .Y(_01878_));
 sky130_fd_sc_hd__nand3_2 _25729_ (.A(_04492_),
    .B(_04524_),
    .C(mem_rdata[29]),
    .Y(_04542_));
 sky130_fd_sc_hd__nand3b_2 _25730_ (.A_N(_04507_),
    .B(_04494_),
    .C(mem_rdata[21]),
    .Y(_04543_));
 sky130_fd_sc_hd__o211a_2 _25731_ (.A1(_01878_),
    .A2(_04490_),
    .B1(_04542_),
    .C1(_04543_),
    .X(_01774_));
 sky130_fd_sc_hd__o2bb2a_2 _25732_ (.A1_N(_04509_),
    .A2_N(_01776_),
    .B1(_01775_),
    .B2(_04527_),
    .X(_01777_));
 sky130_vsdinv _25733_ (.A(_18259_),
    .Y(_01780_));
 sky130_fd_sc_hd__buf_1 _25734_ (.A(_04528_),
    .X(_04544_));
 sky130_fd_sc_hd__and2_2 _25735_ (.A(_04544_),
    .B(_18167_),
    .X(_04545_));
 sky130_fd_sc_hd__a221oi_2 _25736_ (.A1(\count_instr[37] ),
    .A2(_18988_),
    .B1(_17840_),
    .B2(_18991_),
    .C1(_04545_),
    .Y(_01781_));
 sky130_fd_sc_hd__buf_1 _25737_ (.A(_04476_),
    .X(_04546_));
 sky130_fd_sc_hd__buf_1 _25738_ (.A(_04546_),
    .X(_04547_));
 sky130_fd_sc_hd__and2_2 _25739_ (.A(_04514_),
    .B(\timer[5] ),
    .X(_04548_));
 sky130_fd_sc_hd__a221oi_2 _25740_ (.A1(_17199_),
    .A2(_04463_),
    .B1(\cpuregs_rs1[5] ),
    .B2(_04547_),
    .C1(_04548_),
    .Y(_01783_));
 sky130_fd_sc_hd__and2_2 _25741_ (.A(_17580_),
    .B(_19407_),
    .X(_04549_));
 sky130_fd_sc_hd__nor2_2 _25742_ (.A(_17574_),
    .B(_19413_),
    .Y(_04550_));
 sky130_fd_sc_hd__and2_2 _25743_ (.A(\reg_pc[5] ),
    .B(\decoded_imm[5] ),
    .X(_04551_));
 sky130_fd_sc_hd__nor2_2 _25744_ (.A(_04550_),
    .B(_04551_),
    .Y(_04552_));
 sky130_fd_sc_hd__a211oi_2 _25745_ (.A1(_04536_),
    .A2(_04534_),
    .B1(_04549_),
    .C1(_04552_),
    .Y(_04553_));
 sky130_fd_sc_hd__and2_2 _25746_ (.A(_04536_),
    .B(_04534_),
    .X(_04554_));
 sky130_fd_sc_hd__o21a_2 _25747_ (.A1(_04549_),
    .A2(_04554_),
    .B1(_04552_),
    .X(_04555_));
 sky130_fd_sc_hd__buf_1 _25748_ (.A(_17389_),
    .X(_04556_));
 sky130_fd_sc_hd__or2b_2 _25749_ (.A(_01778_),
    .B_N(_04556_),
    .X(_04557_));
 sky130_fd_sc_hd__a2bb2oi_2 _25750_ (.A1_N(_01784_),
    .A2_N(_04487_),
    .B1(_04488_),
    .B2(_01779_),
    .Y(_04558_));
 sky130_fd_sc_hd__o311ai_2 _25751_ (.A1(_04482_),
    .A2(_04553_),
    .A3(_04555_),
    .B1(_04557_),
    .C1(_04558_),
    .Y(_01785_));
 sky130_vsdinv _25752_ (.A(mem_rdata[6]),
    .Y(_01786_));
 sky130_vsdinv _25753_ (.A(mem_rdata[14]),
    .Y(_01891_));
 sky130_fd_sc_hd__nand3_2 _25754_ (.A(_04491_),
    .B(_04524_),
    .C(mem_rdata[30]),
    .Y(_04559_));
 sky130_fd_sc_hd__nand3b_2 _25755_ (.A_N(_04507_),
    .B(_04453_),
    .C(mem_rdata[22]),
    .Y(_04560_));
 sky130_fd_sc_hd__o211a_2 _25756_ (.A1(_01891_),
    .A2(_04443_),
    .B1(_04559_),
    .C1(_04560_),
    .X(_01787_));
 sky130_fd_sc_hd__o2bb2a_2 _25757_ (.A1_N(_04509_),
    .A2_N(_01789_),
    .B1(_01788_),
    .B2(_04527_),
    .X(_01790_));
 sky130_vsdinv _25758_ (.A(_18253_),
    .Y(_01793_));
 sky130_fd_sc_hd__and2_2 _25759_ (.A(_17720_),
    .B(_04511_),
    .X(_04561_));
 sky130_fd_sc_hd__a221oi_2 _25760_ (.A1(_17818_),
    .A2(_04474_),
    .B1(_04530_),
    .B2(_18173_),
    .C1(_04561_),
    .Y(_01794_));
 sky130_fd_sc_hd__buf_1 _25761_ (.A(_04479_),
    .X(_04562_));
 sky130_fd_sc_hd__and2_2 _25762_ (.A(_17196_),
    .B(_04562_),
    .X(_04563_));
 sky130_fd_sc_hd__a221oi_2 _25763_ (.A1(_18953_),
    .A2(_04110_),
    .B1(\cpuregs_rs1[6] ),
    .B2(_04547_),
    .C1(_04563_),
    .Y(_01796_));
 sky130_fd_sc_hd__xor2_2 _25764_ (.A(\reg_pc[6] ),
    .B(_19415_),
    .X(_04564_));
 sky130_vsdinv _25765_ (.A(_04564_),
    .Y(_04565_));
 sky130_fd_sc_hd__o211a_2 _25766_ (.A1(_17574_),
    .A2(_19413_),
    .B1(_17580_),
    .C1(_19407_),
    .X(_04566_));
 sky130_fd_sc_hd__a311oi_2 _25767_ (.A1(_04535_),
    .A2(_04533_),
    .A3(_04552_),
    .B1(_04551_),
    .C1(_04566_),
    .Y(_04567_));
 sky130_fd_sc_hd__nor2_2 _25768_ (.A(_04565_),
    .B(_04567_),
    .Y(_04568_));
 sky130_fd_sc_hd__and2_2 _25769_ (.A(_04567_),
    .B(_04565_),
    .X(_04569_));
 sky130_fd_sc_hd__buf_1 _25770_ (.A(_16822_),
    .X(_04570_));
 sky130_fd_sc_hd__buf_1 _25771_ (.A(_17021_),
    .X(_04571_));
 sky130_fd_sc_hd__buf_1 _25772_ (.A(_17018_),
    .X(_04572_));
 sky130_fd_sc_hd__nand2_2 _25773_ (.A(_04572_),
    .B(_01792_),
    .Y(_04573_));
 sky130_fd_sc_hd__o221a_2 _25774_ (.A1(_01791_),
    .A2(_04570_),
    .B1(_04571_),
    .B2(_01797_),
    .C1(_04573_),
    .X(_04574_));
 sky130_fd_sc_hd__o31ai_2 _25775_ (.A1(_19771_),
    .A2(_04568_),
    .A3(_04569_),
    .B1(_04574_),
    .Y(_01798_));
 sky130_vsdinv _25776_ (.A(mem_rdata[7]),
    .Y(_01799_));
 sky130_vsdinv _25777_ (.A(mem_rdata[15]),
    .Y(_01904_));
 sky130_fd_sc_hd__nand3_2 _25778_ (.A(_04491_),
    .B(_04524_),
    .C(mem_rdata[31]),
    .Y(_04575_));
 sky130_fd_sc_hd__nand3b_2 _25779_ (.A_N(_19543_),
    .B(_04453_),
    .C(mem_rdata[23]),
    .Y(_04576_));
 sky130_fd_sc_hd__o211a_2 _25780_ (.A1(_01904_),
    .A2(_04443_),
    .B1(_04575_),
    .C1(_04576_),
    .X(_01800_));
 sky130_fd_sc_hd__buf_1 _25781_ (.A(_19757_),
    .X(_04577_));
 sky130_fd_sc_hd__o2bb2a_2 _25782_ (.A1_N(_04577_),
    .A2_N(_01802_),
    .B1(_01801_),
    .B2(_04527_),
    .X(_01803_));
 sky130_vsdinv _25783_ (.A(_18254_),
    .Y(_01806_));
 sky130_fd_sc_hd__and2_2 _25784_ (.A(_04544_),
    .B(\count_cycle[39] ),
    .X(_04578_));
 sky130_fd_sc_hd__a221oi_2 _25785_ (.A1(\count_instr[39] ),
    .A2(_18988_),
    .B1(_17837_),
    .B2(_18991_),
    .C1(_04578_),
    .Y(_01807_));
 sky130_fd_sc_hd__buf_1 _25786_ (.A(_04462_),
    .X(_04579_));
 sky130_fd_sc_hd__and2_2 _25787_ (.A(_04514_),
    .B(_04111_),
    .X(_04580_));
 sky130_fd_sc_hd__a221oi_2 _25788_ (.A1(\irq_mask[7] ),
    .A2(_04579_),
    .B1(\cpuregs_rs1[7] ),
    .B2(_04547_),
    .C1(_04580_),
    .Y(_01809_));
 sky130_fd_sc_hd__buf_1 _25789_ (.A(_19661_),
    .X(_04581_));
 sky130_vsdinv _25790_ (.A(_01804_),
    .Y(_04582_));
 sky130_fd_sc_hd__a22oi_2 _25791_ (.A1(_04581_),
    .A2(_01805_),
    .B1(_04582_),
    .B2(_17390_),
    .Y(_04583_));
 sky130_fd_sc_hd__and2_2 _25792_ (.A(\reg_pc[6] ),
    .B(\decoded_imm[6] ),
    .X(_04584_));
 sky130_fd_sc_hd__nor2_2 _25793_ (.A(\reg_pc[7] ),
    .B(_19419_),
    .Y(_04585_));
 sky130_fd_sc_hd__and2_2 _25794_ (.A(\reg_pc[7] ),
    .B(_19419_),
    .X(_04586_));
 sky130_fd_sc_hd__nor2_2 _25795_ (.A(_04585_),
    .B(_04586_),
    .Y(_04587_));
 sky130_fd_sc_hd__o21ai_2 _25796_ (.A1(_04584_),
    .A2(_04568_),
    .B1(_04587_),
    .Y(_04588_));
 sky130_fd_sc_hd__buf_1 _25797_ (.A(_19678_),
    .X(_04589_));
 sky130_vsdinv _25798_ (.A(_04584_),
    .Y(_04590_));
 sky130_fd_sc_hd__o221ai_2 _25799_ (.A1(_04586_),
    .A2(_04585_),
    .B1(_04565_),
    .B2(_04567_),
    .C1(_04590_),
    .Y(_04591_));
 sky130_fd_sc_hd__nand3_2 _25800_ (.A(_04588_),
    .B(_04589_),
    .C(_04591_),
    .Y(_04592_));
 sky130_fd_sc_hd__o211ai_2 _25801_ (.A1(_04470_),
    .A2(_01810_),
    .B1(_04583_),
    .C1(_04592_),
    .Y(_01811_));
 sky130_fd_sc_hd__buf_1 _25802_ (.A(_04437_),
    .X(_04593_));
 sky130_fd_sc_hd__buf_1 _25803_ (.A(_04593_),
    .X(_04594_));
 sky130_fd_sc_hd__nand2_2 _25804_ (.A(_04594_),
    .B(_01813_),
    .Y(_01814_));
 sky130_fd_sc_hd__nor2_2 _25805_ (.A(latched_is_lb),
    .B(latched_is_lh),
    .Y(_01816_));
 sky130_vsdinv _25806_ (.A(latched_is_lh),
    .Y(_04595_));
 sky130_fd_sc_hd__buf_1 _25807_ (.A(_04595_),
    .X(_04596_));
 sky130_fd_sc_hd__nand2_2 _25808_ (.A(_04582_),
    .B(latched_is_lb),
    .Y(_04597_));
 sky130_fd_sc_hd__buf_1 _25809_ (.A(_04597_),
    .X(_04598_));
 sky130_fd_sc_hd__o21a_2 _25810_ (.A1(_04596_),
    .A2(_01815_),
    .B1(_04598_),
    .X(_01817_));
 sky130_fd_sc_hd__buf_1 _25811_ (.A(instr_rdinstrh),
    .X(_04599_));
 sky130_fd_sc_hd__buf_1 _25812_ (.A(_04599_),
    .X(_04600_));
 sky130_fd_sc_hd__buf_1 _25813_ (.A(_04459_),
    .X(_04601_));
 sky130_fd_sc_hd__and2_2 _25814_ (.A(\count_instr[8] ),
    .B(_04601_),
    .X(_04602_));
 sky130_fd_sc_hd__a221oi_2 _25815_ (.A1(_17711_),
    .A2(_04600_),
    .B1(_04530_),
    .B2(_18163_),
    .C1(_04602_),
    .Y(_01821_));
 sky130_fd_sc_hd__buf_1 _25816_ (.A(_04513_),
    .X(_04603_));
 sky130_fd_sc_hd__and2_2 _25817_ (.A(_04603_),
    .B(_04113_),
    .X(_04604_));
 sky130_fd_sc_hd__a221oi_2 _25818_ (.A1(_17187_),
    .A2(_04579_),
    .B1(\cpuregs_rs1[8] ),
    .B2(_04547_),
    .C1(_04604_),
    .Y(_01823_));
 sky130_fd_sc_hd__xor2_2 _25819_ (.A(\reg_pc[8] ),
    .B(_19422_),
    .X(_04605_));
 sky130_fd_sc_hd__nand2_2 _25820_ (.A(_04564_),
    .B(_04587_),
    .Y(_04606_));
 sky130_fd_sc_hd__o21ba_2 _25821_ (.A1(_04585_),
    .A2(_04590_),
    .B1_N(_04586_),
    .X(_04607_));
 sky130_fd_sc_hd__o21ai_2 _25822_ (.A1(_04606_),
    .A2(_04567_),
    .B1(_04607_),
    .Y(_04608_));
 sky130_fd_sc_hd__o21a_2 _25823_ (.A1(_04605_),
    .A2(_04608_),
    .B1(_19517_),
    .X(_04609_));
 sky130_fd_sc_hd__nand2_2 _25824_ (.A(_04608_),
    .B(_04605_),
    .Y(_04610_));
 sky130_fd_sc_hd__and2b_2 _25825_ (.A_N(_01818_),
    .B(_04073_),
    .X(_04611_));
 sky130_fd_sc_hd__o2bb2ai_2 _25826_ (.A1_N(_04581_),
    .A2_N(_01819_),
    .B1(_01824_),
    .B2(_04487_),
    .Y(_04612_));
 sky130_fd_sc_hd__a211o_2 _25827_ (.A1(_04609_),
    .A2(_04610_),
    .B1(_04611_),
    .C1(_04612_),
    .X(_01825_));
 sky130_fd_sc_hd__nand2_2 _25828_ (.A(_04594_),
    .B(_01827_),
    .Y(_01828_));
 sky130_fd_sc_hd__o21a_2 _25829_ (.A1(_04596_),
    .A2(_01829_),
    .B1(_04598_),
    .X(_01830_));
 sky130_fd_sc_hd__buf_1 _25830_ (.A(_18990_),
    .X(_04613_));
 sky130_fd_sc_hd__and2_2 _25831_ (.A(_04544_),
    .B(_18164_),
    .X(_04614_));
 sky130_fd_sc_hd__a221oi_2 _25832_ (.A1(_17710_),
    .A2(_04600_),
    .B1(_17812_),
    .B2(_04613_),
    .C1(_04614_),
    .Y(_01834_));
 sky130_fd_sc_hd__buf_1 _25833_ (.A(_18952_),
    .X(_04615_));
 sky130_fd_sc_hd__buf_1 _25834_ (.A(_04546_),
    .X(_04616_));
 sky130_fd_sc_hd__and2_2 _25835_ (.A(_17183_),
    .B(_04562_),
    .X(_04617_));
 sky130_fd_sc_hd__a221oi_2 _25836_ (.A1(_04615_),
    .A2(\timer[9] ),
    .B1(\cpuregs_rs1[9] ),
    .B2(_04616_),
    .C1(_04617_),
    .Y(_01836_));
 sky130_fd_sc_hd__buf_1 _25837_ (.A(_16824_),
    .X(_04618_));
 sky130_fd_sc_hd__buf_1 _25838_ (.A(_04469_),
    .X(_04619_));
 sky130_fd_sc_hd__a2bb2oi_2 _25839_ (.A1_N(_01837_),
    .A2_N(_04619_),
    .B1(_04522_),
    .B2(_01832_),
    .Y(_04620_));
 sky130_fd_sc_hd__and2_2 _25840_ (.A(\reg_pc[8] ),
    .B(_19422_),
    .X(_04621_));
 sky130_vsdinv _25841_ (.A(_04621_),
    .Y(_04622_));
 sky130_fd_sc_hd__nor2_2 _25842_ (.A(_17557_),
    .B(_19425_),
    .Y(_04623_));
 sky130_fd_sc_hd__and2_2 _25843_ (.A(\reg_pc[9] ),
    .B(_19425_),
    .X(_04624_));
 sky130_fd_sc_hd__nor2_2 _25844_ (.A(_04623_),
    .B(_04624_),
    .Y(_04625_));
 sky130_vsdinv _25845_ (.A(_04625_),
    .Y(_04626_));
 sky130_fd_sc_hd__a21o_2 _25846_ (.A1(_04610_),
    .A2(_04622_),
    .B1(_04626_),
    .X(_04627_));
 sky130_fd_sc_hd__nand3_2 _25847_ (.A(_04610_),
    .B(_04622_),
    .C(_04626_),
    .Y(_04628_));
 sky130_fd_sc_hd__nand3_2 _25848_ (.A(_04627_),
    .B(_04589_),
    .C(_04628_),
    .Y(_04629_));
 sky130_fd_sc_hd__o211ai_2 _25849_ (.A1(_04618_),
    .A2(_01831_),
    .B1(_04620_),
    .C1(_04629_),
    .Y(_01838_));
 sky130_fd_sc_hd__nand2_2 _25850_ (.A(_04594_),
    .B(_01840_),
    .Y(_01841_));
 sky130_fd_sc_hd__o21a_2 _25851_ (.A1(_04596_),
    .A2(_01842_),
    .B1(_04598_),
    .X(_01843_));
 sky130_fd_sc_hd__buf_1 _25852_ (.A(_04459_),
    .X(_04630_));
 sky130_fd_sc_hd__and2_2 _25853_ (.A(\count_instr[42] ),
    .B(_04511_),
    .X(_04631_));
 sky130_fd_sc_hd__a221oi_2 _25854_ (.A1(_17823_),
    .A2(_04630_),
    .B1(_04530_),
    .B2(_18149_),
    .C1(_04631_),
    .Y(_01847_));
 sky130_fd_sc_hd__and2_2 _25855_ (.A(_04603_),
    .B(\timer[10] ),
    .X(_04632_));
 sky130_fd_sc_hd__a221oi_2 _25856_ (.A1(_17180_),
    .A2(_04579_),
    .B1(\cpuregs_rs1[10] ),
    .B2(_04616_),
    .C1(_04632_),
    .Y(_01849_));
 sky130_fd_sc_hd__buf_1 _25857_ (.A(_16985_),
    .X(_04633_));
 sky130_fd_sc_hd__and2_2 _25858_ (.A(\reg_pc[10] ),
    .B(_19427_),
    .X(_04634_));
 sky130_fd_sc_hd__nor2_2 _25859_ (.A(_17552_),
    .B(_19427_),
    .Y(_04635_));
 sky130_fd_sc_hd__o21bai_2 _25860_ (.A1(_04623_),
    .A2(_04622_),
    .B1_N(_04624_),
    .Y(_04636_));
 sky130_fd_sc_hd__a31oi_2 _25861_ (.A1(_04608_),
    .A2(_04605_),
    .A3(_04625_),
    .B1(_04636_),
    .Y(_04637_));
 sky130_fd_sc_hd__o21a_2 _25862_ (.A1(_04634_),
    .A2(_04635_),
    .B1(_04637_),
    .X(_04638_));
 sky130_fd_sc_hd__nor3_2 _25863_ (.A(_04634_),
    .B(_04635_),
    .C(_04637_),
    .Y(_04639_));
 sky130_fd_sc_hd__nand2_2 _25864_ (.A(_04572_),
    .B(_01845_),
    .Y(_04640_));
 sky130_fd_sc_hd__o221a_2 _25865_ (.A1(_01844_),
    .A2(_04570_),
    .B1(_04571_),
    .B2(_01850_),
    .C1(_04640_),
    .X(_04641_));
 sky130_fd_sc_hd__o31ai_2 _25866_ (.A1(_04633_),
    .A2(_04638_),
    .A3(_04639_),
    .B1(_04641_),
    .Y(_01851_));
 sky130_fd_sc_hd__nand2_2 _25867_ (.A(_04594_),
    .B(_01853_),
    .Y(_01854_));
 sky130_fd_sc_hd__o21a_2 _25868_ (.A1(_04596_),
    .A2(_01855_),
    .B1(_04598_),
    .X(_01856_));
 sky130_fd_sc_hd__buf_1 _25869_ (.A(_18996_),
    .X(_04642_));
 sky130_fd_sc_hd__buf_1 _25870_ (.A(instr_rdinstr),
    .X(_04643_));
 sky130_fd_sc_hd__and2_2 _25871_ (.A(_17826_),
    .B(_04643_),
    .X(_04644_));
 sky130_fd_sc_hd__a221oi_2 _25872_ (.A1(_17686_),
    .A2(_04600_),
    .B1(_04642_),
    .B2(_18146_),
    .C1(_04644_),
    .Y(_01860_));
 sky130_fd_sc_hd__and2_2 _25873_ (.A(_04603_),
    .B(_04117_),
    .X(_04645_));
 sky130_fd_sc_hd__a221oi_2 _25874_ (.A1(\irq_mask[11] ),
    .A2(_04579_),
    .B1(\cpuregs_rs1[11] ),
    .B2(_04616_),
    .C1(_04645_),
    .Y(_01862_));
 sky130_fd_sc_hd__and2_2 _25875_ (.A(\reg_pc[11] ),
    .B(_19429_),
    .X(_04646_));
 sky130_vsdinv _25876_ (.A(_04646_),
    .Y(_04647_));
 sky130_fd_sc_hd__or2_2 _25877_ (.A(\reg_pc[11] ),
    .B(_19429_),
    .X(_04648_));
 sky130_fd_sc_hd__o21bai_2 _25878_ (.A1(_04635_),
    .A2(_04637_),
    .B1_N(_04634_),
    .Y(_04649_));
 sky130_fd_sc_hd__a21o_2 _25879_ (.A1(_04647_),
    .A2(_04648_),
    .B1(_04649_),
    .X(_04650_));
 sky130_fd_sc_hd__nand3_2 _25880_ (.A(_04649_),
    .B(_04647_),
    .C(_04648_),
    .Y(_04651_));
 sky130_fd_sc_hd__and2b_2 _25881_ (.A_N(_01857_),
    .B(_04073_),
    .X(_04652_));
 sky130_fd_sc_hd__o2bb2ai_2 _25882_ (.A1_N(_04450_),
    .A2_N(_01858_),
    .B1(_01863_),
    .B2(_04540_),
    .Y(_04653_));
 sky130_fd_sc_hd__a311o_2 _25883_ (.A1(_04650_),
    .A2(_04651_),
    .A3(_19679_),
    .B1(_04652_),
    .C1(_04653_),
    .X(_01864_));
 sky130_fd_sc_hd__buf_1 _25884_ (.A(_04593_),
    .X(_04654_));
 sky130_fd_sc_hd__nand2_2 _25885_ (.A(_04654_),
    .B(_01866_),
    .Y(_01867_));
 sky130_fd_sc_hd__buf_1 _25886_ (.A(_04595_),
    .X(_04655_));
 sky130_fd_sc_hd__buf_1 _25887_ (.A(_04597_),
    .X(_04656_));
 sky130_fd_sc_hd__o21a_2 _25888_ (.A1(_04655_),
    .A2(_01868_),
    .B1(_04656_),
    .X(_01869_));
 sky130_fd_sc_hd__and2_2 _25889_ (.A(_04544_),
    .B(_18150_),
    .X(_04657_));
 sky130_fd_sc_hd__a221oi_2 _25890_ (.A1(_17702_),
    .A2(_04600_),
    .B1(\count_instr[12] ),
    .B2(_04613_),
    .C1(_04657_),
    .Y(_01873_));
 sky130_fd_sc_hd__and2_2 _25891_ (.A(_17176_),
    .B(_04562_),
    .X(_04658_));
 sky130_fd_sc_hd__a221oi_2 _25892_ (.A1(_04615_),
    .A2(\timer[12] ),
    .B1(\cpuregs_rs1[12] ),
    .B2(_04616_),
    .C1(_04658_),
    .Y(_01875_));
 sky130_fd_sc_hd__nor2_2 _25893_ (.A(_17545_),
    .B(_19440_),
    .Y(_04659_));
 sky130_fd_sc_hd__and2_2 _25894_ (.A(\reg_pc[12] ),
    .B(_19440_),
    .X(_04660_));
 sky130_fd_sc_hd__nor2_2 _25895_ (.A(_04659_),
    .B(_04660_),
    .Y(_04661_));
 sky130_fd_sc_hd__a211oi_2 _25896_ (.A1(_04649_),
    .A2(_04648_),
    .B1(_04646_),
    .C1(_04661_),
    .Y(_04662_));
 sky130_fd_sc_hd__a21boi_2 _25897_ (.A1(_04651_),
    .A2(_04647_),
    .B1_N(_04661_),
    .Y(_04663_));
 sky130_fd_sc_hd__nand2_2 _25898_ (.A(_04572_),
    .B(_01871_),
    .Y(_04664_));
 sky130_fd_sc_hd__o221a_2 _25899_ (.A1(_01870_),
    .A2(_04570_),
    .B1(_04571_),
    .B2(_01876_),
    .C1(_04664_),
    .X(_04665_));
 sky130_fd_sc_hd__o31ai_2 _25900_ (.A1(_04633_),
    .A2(_04662_),
    .A3(_04663_),
    .B1(_04665_),
    .Y(_01877_));
 sky130_fd_sc_hd__nand2_2 _25901_ (.A(_04654_),
    .B(_01879_),
    .Y(_01880_));
 sky130_fd_sc_hd__o21a_2 _25902_ (.A1(_04655_),
    .A2(_01881_),
    .B1(_04656_),
    .X(_01882_));
 sky130_vsdinv _25903_ (.A(_18237_),
    .Y(_01885_));
 sky130_fd_sc_hd__buf_1 _25904_ (.A(_04599_),
    .X(_04666_));
 sky130_fd_sc_hd__and2_2 _25905_ (.A(_17797_),
    .B(_04643_),
    .X(_04667_));
 sky130_fd_sc_hd__a221oi_2 _25906_ (.A1(_17701_),
    .A2(_04666_),
    .B1(_04642_),
    .B2(_18157_),
    .C1(_04667_),
    .Y(_01886_));
 sky130_fd_sc_hd__buf_1 _25907_ (.A(_04462_),
    .X(_04668_));
 sky130_fd_sc_hd__buf_1 _25908_ (.A(_04546_),
    .X(_04669_));
 sky130_fd_sc_hd__and2_2 _25909_ (.A(_04603_),
    .B(\timer[13] ),
    .X(_04670_));
 sky130_fd_sc_hd__a221oi_2 _25910_ (.A1(_17170_),
    .A2(_04668_),
    .B1(\cpuregs_rs1[13] ),
    .B2(_04669_),
    .C1(_04670_),
    .Y(_01888_));
 sky130_fd_sc_hd__and2_2 _25911_ (.A(\reg_pc[13] ),
    .B(_19444_),
    .X(_04671_));
 sky130_vsdinv _25912_ (.A(_04671_),
    .Y(_04672_));
 sky130_fd_sc_hd__or2_2 _25913_ (.A(\reg_pc[13] ),
    .B(_19444_),
    .X(_04673_));
 sky130_fd_sc_hd__a21oi_2 _25914_ (.A1(_04649_),
    .A2(_04648_),
    .B1(_04646_),
    .Y(_04674_));
 sky130_fd_sc_hd__o21bai_2 _25915_ (.A1(_04659_),
    .A2(_04674_),
    .B1_N(_04660_),
    .Y(_04675_));
 sky130_fd_sc_hd__a21o_2 _25916_ (.A1(_04672_),
    .A2(_04673_),
    .B1(_04675_),
    .X(_04676_));
 sky130_fd_sc_hd__nand3_2 _25917_ (.A(_04675_),
    .B(_04672_),
    .C(_04673_),
    .Y(_04677_));
 sky130_fd_sc_hd__buf_1 _25918_ (.A(_19759_),
    .X(_04678_));
 sky130_fd_sc_hd__and2b_2 _25919_ (.A_N(_01883_),
    .B(_04678_),
    .X(_04679_));
 sky130_fd_sc_hd__buf_1 _25920_ (.A(_18540_),
    .X(_04680_));
 sky130_fd_sc_hd__o2bb2ai_2 _25921_ (.A1_N(_04450_),
    .A2_N(_01884_),
    .B1(_01889_),
    .B2(_04680_),
    .Y(_04681_));
 sky130_fd_sc_hd__a311o_2 _25922_ (.A1(_04676_),
    .A2(_04677_),
    .A3(_19679_),
    .B1(_04679_),
    .C1(_04681_),
    .X(_01890_));
 sky130_fd_sc_hd__nand2_2 _25923_ (.A(_04654_),
    .B(_01892_),
    .Y(_01893_));
 sky130_fd_sc_hd__o21a_2 _25924_ (.A1(_04655_),
    .A2(_01894_),
    .B1(_04656_),
    .X(_01895_));
 sky130_fd_sc_hd__buf_1 _25925_ (.A(_04510_),
    .X(_04682_));
 sky130_fd_sc_hd__and2_2 _25926_ (.A(\count_instr[46] ),
    .B(_04682_),
    .X(_04683_));
 sky130_fd_sc_hd__a221oi_2 _25927_ (.A1(_17805_),
    .A2(_04630_),
    .B1(_04642_),
    .B2(_18152_),
    .C1(_04683_),
    .Y(_01899_));
 sky130_fd_sc_hd__and2_2 _25928_ (.A(_17166_),
    .B(_04562_),
    .X(_04684_));
 sky130_fd_sc_hd__a221oi_2 _25929_ (.A1(_04615_),
    .A2(\timer[14] ),
    .B1(\cpuregs_rs1[14] ),
    .B2(_04669_),
    .C1(_04684_),
    .Y(_01901_));
 sky130_fd_sc_hd__nor2_2 _25930_ (.A(\reg_pc[14] ),
    .B(_19445_),
    .Y(_04685_));
 sky130_fd_sc_hd__and2_2 _25931_ (.A(\reg_pc[14] ),
    .B(_19445_),
    .X(_04686_));
 sky130_fd_sc_hd__nor2_2 _25932_ (.A(_04685_),
    .B(_04686_),
    .Y(_04687_));
 sky130_fd_sc_hd__a211oi_2 _25933_ (.A1(_04675_),
    .A2(_04673_),
    .B1(_04671_),
    .C1(_04687_),
    .Y(_04688_));
 sky130_fd_sc_hd__a21boi_2 _25934_ (.A1(_04677_),
    .A2(_04672_),
    .B1_N(_04687_),
    .Y(_04689_));
 sky130_fd_sc_hd__nand2_2 _25935_ (.A(_04572_),
    .B(_01897_),
    .Y(_04690_));
 sky130_fd_sc_hd__o221a_2 _25936_ (.A1(_01896_),
    .A2(_04570_),
    .B1(_04571_),
    .B2(_01902_),
    .C1(_04690_),
    .X(_04691_));
 sky130_fd_sc_hd__o31ai_2 _25937_ (.A1(_04633_),
    .A2(_04688_),
    .A3(_04689_),
    .B1(_04691_),
    .Y(_01903_));
 sky130_fd_sc_hd__nand2_2 _25938_ (.A(_04654_),
    .B(_01905_),
    .Y(_01906_));
 sky130_fd_sc_hd__o21a_2 _25939_ (.A1(_04655_),
    .A2(_01907_),
    .B1(_04656_),
    .X(_01908_));
 sky130_vsdinv _25940_ (.A(\count_cycle[15] ),
    .Y(_01911_));
 sky130_fd_sc_hd__and2_2 _25941_ (.A(\count_instr[15] ),
    .B(_04643_),
    .X(_04692_));
 sky130_fd_sc_hd__a221oi_2 _25942_ (.A1(\count_instr[47] ),
    .A2(_04666_),
    .B1(_04642_),
    .B2(\count_cycle[47] ),
    .C1(_04692_),
    .Y(_01912_));
 sky130_fd_sc_hd__buf_1 _25943_ (.A(_04479_),
    .X(_04693_));
 sky130_fd_sc_hd__and2_2 _25944_ (.A(_17931_),
    .B(_04693_),
    .X(_04694_));
 sky130_fd_sc_hd__a221oi_2 _25945_ (.A1(_04615_),
    .A2(_04121_),
    .B1(\cpuregs_rs1[15] ),
    .B2(_04669_),
    .C1(_04694_),
    .Y(_01914_));
 sky130_fd_sc_hd__and2_2 _25946_ (.A(_17529_),
    .B(_19454_),
    .X(_04695_));
 sky130_vsdinv _25947_ (.A(_04695_),
    .Y(_04696_));
 sky130_fd_sc_hd__or2_2 _25948_ (.A(\reg_pc[15] ),
    .B(_19454_),
    .X(_04697_));
 sky130_fd_sc_hd__a21oi_2 _25949_ (.A1(_04675_),
    .A2(_04673_),
    .B1(_04671_),
    .Y(_04698_));
 sky130_fd_sc_hd__o21bai_2 _25950_ (.A1(_04685_),
    .A2(_04698_),
    .B1_N(_04686_),
    .Y(_04699_));
 sky130_fd_sc_hd__a21o_2 _25951_ (.A1(_04696_),
    .A2(_04697_),
    .B1(_04699_),
    .X(_04700_));
 sky130_fd_sc_hd__nand3_2 _25952_ (.A(_04699_),
    .B(_04696_),
    .C(_04697_),
    .Y(_04701_));
 sky130_fd_sc_hd__buf_1 _25953_ (.A(_19517_),
    .X(_04702_));
 sky130_fd_sc_hd__and2b_2 _25954_ (.A_N(_01909_),
    .B(_04678_),
    .X(_04703_));
 sky130_fd_sc_hd__buf_1 _25955_ (.A(_17018_),
    .X(_04704_));
 sky130_fd_sc_hd__o2bb2ai_2 _25956_ (.A1_N(_04704_),
    .A2_N(_01910_),
    .B1(_01915_),
    .B2(_04680_),
    .Y(_04705_));
 sky130_fd_sc_hd__a311o_2 _25957_ (.A1(_04700_),
    .A2(_04701_),
    .A3(_04702_),
    .B1(_04703_),
    .C1(_04705_),
    .X(_01916_));
 sky130_fd_sc_hd__buf_1 _25958_ (.A(_19568_),
    .X(_04706_));
 sky130_fd_sc_hd__buf_1 _25959_ (.A(_04706_),
    .X(_04707_));
 sky130_fd_sc_hd__buf_1 _25960_ (.A(_04457_),
    .X(_04708_));
 sky130_fd_sc_hd__buf_1 _25961_ (.A(_04708_),
    .X(_04709_));
 sky130_fd_sc_hd__nand3_2 _25962_ (.A(_04707_),
    .B(_04709_),
    .C(mem_rdata[16]),
    .Y(_01917_));
 sky130_vsdinv _25963_ (.A(_18234_),
    .Y(_01920_));
 sky130_fd_sc_hd__buf_1 _25964_ (.A(_04528_),
    .X(_04710_));
 sky130_fd_sc_hd__and2_2 _25965_ (.A(_04710_),
    .B(_18142_),
    .X(_04711_));
 sky130_fd_sc_hd__a221oi_2 _25966_ (.A1(_17681_),
    .A2(_04666_),
    .B1(_17795_),
    .B2(_04613_),
    .C1(_04711_),
    .Y(_01921_));
 sky130_fd_sc_hd__buf_1 _25967_ (.A(_04513_),
    .X(_04712_));
 sky130_fd_sc_hd__and2_2 _25968_ (.A(_04712_),
    .B(\timer[16] ),
    .X(_04713_));
 sky130_fd_sc_hd__a221oi_2 _25969_ (.A1(_17162_),
    .A2(_04668_),
    .B1(\cpuregs_rs1[16] ),
    .B2(_04669_),
    .C1(_04713_),
    .Y(_01923_));
 sky130_fd_sc_hd__xor2_2 _25970_ (.A(\reg_pc[16] ),
    .B(_19458_),
    .X(_04714_));
 sky130_fd_sc_hd__a21bo_2 _25971_ (.A1(_04701_),
    .A2(_04696_),
    .B1_N(_04714_),
    .X(_04715_));
 sky130_fd_sc_hd__nand3b_2 _25972_ (.A_N(_04714_),
    .B(_04701_),
    .C(_04696_),
    .Y(_04716_));
 sky130_fd_sc_hd__nand2_2 _25973_ (.A(_18003_),
    .B(_01919_),
    .Y(_04717_));
 sky130_fd_sc_hd__o221ai_2 _25974_ (.A1(_01918_),
    .A2(_17384_),
    .B1(_01924_),
    .B2(_18541_),
    .C1(_04717_),
    .Y(_04718_));
 sky130_fd_sc_hd__a31o_2 _25975_ (.A1(_04715_),
    .A2(_19766_),
    .A3(_04716_),
    .B1(_04718_),
    .X(_01925_));
 sky130_fd_sc_hd__nand3_2 _25976_ (.A(_04707_),
    .B(_04709_),
    .C(mem_rdata[17]),
    .Y(_01926_));
 sky130_vsdinv _25977_ (.A(_18232_),
    .Y(_01929_));
 sky130_fd_sc_hd__buf_1 _25978_ (.A(_18996_),
    .X(_04719_));
 sky130_fd_sc_hd__and2_2 _25979_ (.A(\count_instr[49] ),
    .B(_04682_),
    .X(_04720_));
 sky130_fd_sc_hd__a221oi_2 _25980_ (.A1(_17792_),
    .A2(_04630_),
    .B1(_04719_),
    .B2(_18138_),
    .C1(_04720_),
    .Y(_01930_));
 sky130_fd_sc_hd__buf_1 _25981_ (.A(_04546_),
    .X(_04721_));
 sky130_fd_sc_hd__and2_2 _25982_ (.A(_04712_),
    .B(\timer[17] ),
    .X(_04722_));
 sky130_fd_sc_hd__a221oi_2 _25983_ (.A1(_17159_),
    .A2(_04668_),
    .B1(\cpuregs_rs1[17] ),
    .B2(_04721_),
    .C1(_04722_),
    .Y(_01932_));
 sky130_fd_sc_hd__a2bb2oi_2 _25984_ (.A1_N(_01933_),
    .A2_N(_04619_),
    .B1(_04522_),
    .B2(_01928_),
    .Y(_04723_));
 sky130_fd_sc_hd__and2_2 _25985_ (.A(\reg_pc[16] ),
    .B(\decoded_imm[16] ),
    .X(_04724_));
 sky130_vsdinv _25986_ (.A(_04724_),
    .Y(_04725_));
 sky130_fd_sc_hd__nor2_2 _25987_ (.A(\reg_pc[17] ),
    .B(_19462_),
    .Y(_04726_));
 sky130_fd_sc_hd__and2_2 _25988_ (.A(\reg_pc[17] ),
    .B(\decoded_imm[17] ),
    .X(_04727_));
 sky130_fd_sc_hd__nor2_2 _25989_ (.A(_04726_),
    .B(_04727_),
    .Y(_04728_));
 sky130_fd_sc_hd__a21bo_2 _25990_ (.A1(_04715_),
    .A2(_04725_),
    .B1_N(_04728_),
    .X(_04729_));
 sky130_fd_sc_hd__nand3b_2 _25991_ (.A_N(_04728_),
    .B(_04715_),
    .C(_04725_),
    .Y(_04730_));
 sky130_fd_sc_hd__nand3_2 _25992_ (.A(_04729_),
    .B(_04589_),
    .C(_04730_),
    .Y(_04731_));
 sky130_fd_sc_hd__o211ai_2 _25993_ (.A1(_04618_),
    .A2(_01927_),
    .B1(_04723_),
    .C1(_04731_),
    .Y(_01934_));
 sky130_fd_sc_hd__nand3_2 _25994_ (.A(_04707_),
    .B(_04709_),
    .C(mem_rdata[18]),
    .Y(_01935_));
 sky130_fd_sc_hd__and2_2 _25995_ (.A(_17675_),
    .B(_04682_),
    .X(_04732_));
 sky130_fd_sc_hd__a221oi_2 _25996_ (.A1(_17789_),
    .A2(_04630_),
    .B1(_04719_),
    .B2(_18139_),
    .C1(_04732_),
    .Y(_01939_));
 sky130_fd_sc_hd__buf_1 _25997_ (.A(_18952_),
    .X(_04733_));
 sky130_fd_sc_hd__and2_2 _25998_ (.A(_17157_),
    .B(_04693_),
    .X(_04734_));
 sky130_fd_sc_hd__a221oi_2 _25999_ (.A1(_04733_),
    .A2(\timer[18] ),
    .B1(\cpuregs_rs1[18] ),
    .B2(_04721_),
    .C1(_04734_),
    .Y(_01941_));
 sky130_fd_sc_hd__and2_2 _26000_ (.A(\reg_pc[18] ),
    .B(_19465_),
    .X(_04735_));
 sky130_vsdinv _26001_ (.A(_04735_),
    .Y(_04736_));
 sky130_fd_sc_hd__or2_2 _26002_ (.A(\reg_pc[18] ),
    .B(\decoded_imm[18] ),
    .X(_04737_));
 sky130_fd_sc_hd__nand2_2 _26003_ (.A(_04714_),
    .B(_04728_),
    .Y(_04738_));
 sky130_fd_sc_hd__a21oi_2 _26004_ (.A1(_04699_),
    .A2(_04697_),
    .B1(_04695_),
    .Y(_04739_));
 sky130_fd_sc_hd__o21bai_2 _26005_ (.A1(_04726_),
    .A2(_04725_),
    .B1_N(_04727_),
    .Y(_04740_));
 sky130_fd_sc_hd__o21bai_2 _26006_ (.A1(_04738_),
    .A2(_04739_),
    .B1_N(_04740_),
    .Y(_04741_));
 sky130_fd_sc_hd__a21o_2 _26007_ (.A1(_04736_),
    .A2(_04737_),
    .B1(_04741_),
    .X(_04742_));
 sky130_fd_sc_hd__nand3_2 _26008_ (.A(_04741_),
    .B(_04736_),
    .C(_04737_),
    .Y(_04743_));
 sky130_fd_sc_hd__and2b_2 _26009_ (.A_N(_01936_),
    .B(_04678_),
    .X(_04744_));
 sky130_fd_sc_hd__o2bb2ai_2 _26010_ (.A1_N(_04704_),
    .A2_N(_01937_),
    .B1(_01942_),
    .B2(_04680_),
    .Y(_04745_));
 sky130_fd_sc_hd__a311o_2 _26011_ (.A1(_04742_),
    .A2(_04743_),
    .A3(_04702_),
    .B1(_04744_),
    .C1(_04745_),
    .X(_01943_));
 sky130_fd_sc_hd__nand3_2 _26012_ (.A(_04707_),
    .B(_04709_),
    .C(mem_rdata[19]),
    .Y(_01944_));
 sky130_fd_sc_hd__and2_2 _26013_ (.A(_04710_),
    .B(_18136_),
    .X(_04746_));
 sky130_fd_sc_hd__a221oi_2 _26014_ (.A1(_17677_),
    .A2(_04666_),
    .B1(_17787_),
    .B2(_04613_),
    .C1(_04746_),
    .Y(_01948_));
 sky130_fd_sc_hd__and2_2 _26015_ (.A(_04712_),
    .B(\timer[19] ),
    .X(_04747_));
 sky130_fd_sc_hd__a221oi_2 _26016_ (.A1(_17154_),
    .A2(_04668_),
    .B1(\cpuregs_rs1[19] ),
    .B2(_04721_),
    .C1(_04747_),
    .Y(_01950_));
 sky130_fd_sc_hd__nor2_2 _26017_ (.A(_17509_),
    .B(_19468_),
    .Y(_04748_));
 sky130_fd_sc_hd__and2_2 _26018_ (.A(\reg_pc[19] ),
    .B(\decoded_imm[19] ),
    .X(_04749_));
 sky130_fd_sc_hd__nor2_2 _26019_ (.A(_04748_),
    .B(_04749_),
    .Y(_04750_));
 sky130_fd_sc_hd__a211oi_2 _26020_ (.A1(_04741_),
    .A2(_04737_),
    .B1(_04735_),
    .C1(_04750_),
    .Y(_04751_));
 sky130_fd_sc_hd__a21boi_2 _26021_ (.A1(_04743_),
    .A2(_04736_),
    .B1_N(_04750_),
    .Y(_04752_));
 sky130_fd_sc_hd__or2b_2 _26022_ (.A(_01945_),
    .B_N(_04556_),
    .X(_04753_));
 sky130_fd_sc_hd__a2bb2oi_2 _26023_ (.A1_N(_01951_),
    .A2_N(_04487_),
    .B1(_04488_),
    .B2(_01946_),
    .Y(_04754_));
 sky130_fd_sc_hd__o311ai_2 _26024_ (.A1(_04482_),
    .A2(_04751_),
    .A3(_04752_),
    .B1(_04753_),
    .C1(_04754_),
    .Y(_01952_));
 sky130_fd_sc_hd__buf_1 _26025_ (.A(_04706_),
    .X(_04755_));
 sky130_fd_sc_hd__buf_1 _26026_ (.A(_04708_),
    .X(_04756_));
 sky130_fd_sc_hd__nand3_2 _26027_ (.A(_04755_),
    .B(_04756_),
    .C(mem_rdata[20]),
    .Y(_01953_));
 sky130_fd_sc_hd__buf_1 _26028_ (.A(_04510_),
    .X(_04757_));
 sky130_fd_sc_hd__and2_2 _26029_ (.A(_17783_),
    .B(_04643_),
    .X(_04758_));
 sky130_fd_sc_hd__a221oi_2 _26030_ (.A1(_17671_),
    .A2(_04757_),
    .B1(_04719_),
    .B2(_18124_),
    .C1(_04758_),
    .Y(_01957_));
 sky130_fd_sc_hd__and2_2 _26031_ (.A(_17151_),
    .B(_04693_),
    .X(_04759_));
 sky130_fd_sc_hd__a221oi_2 _26032_ (.A1(_04733_),
    .A2(\timer[20] ),
    .B1(\cpuregs_rs1[20] ),
    .B2(_04721_),
    .C1(_04759_),
    .Y(_01959_));
 sky130_fd_sc_hd__a2bb2oi_2 _26033_ (.A1_N(_01960_),
    .A2_N(_04619_),
    .B1(_04522_),
    .B2(_01955_),
    .Y(_04760_));
 sky130_fd_sc_hd__and2_2 _26034_ (.A(\reg_pc[20] ),
    .B(_04145_),
    .X(_04761_));
 sky130_vsdinv _26035_ (.A(_04761_),
    .Y(_04762_));
 sky130_fd_sc_hd__nand2_2 _26036_ (.A(_17507_),
    .B(_19478_),
    .Y(_04763_));
 sky130_fd_sc_hd__a21oi_2 _26037_ (.A1(_04741_),
    .A2(_04737_),
    .B1(_04735_),
    .Y(_04764_));
 sky130_fd_sc_hd__o21bai_2 _26038_ (.A1(_04748_),
    .A2(_04764_),
    .B1_N(_04749_),
    .Y(_04765_));
 sky130_fd_sc_hd__a21o_2 _26039_ (.A1(_04762_),
    .A2(_04763_),
    .B1(_04765_),
    .X(_04766_));
 sky130_fd_sc_hd__buf_1 _26040_ (.A(_19678_),
    .X(_04767_));
 sky130_fd_sc_hd__nand3_2 _26041_ (.A(_04765_),
    .B(_04762_),
    .C(_04763_),
    .Y(_04768_));
 sky130_fd_sc_hd__nand3_2 _26042_ (.A(_04766_),
    .B(_04767_),
    .C(_04768_),
    .Y(_04769_));
 sky130_fd_sc_hd__o211ai_2 _26043_ (.A1(_04618_),
    .A2(_01954_),
    .B1(_04760_),
    .C1(_04769_),
    .Y(_01961_));
 sky130_fd_sc_hd__nand3_2 _26044_ (.A(_04755_),
    .B(_04756_),
    .C(mem_rdata[21]),
    .Y(_01962_));
 sky130_vsdinv _26045_ (.A(_18221_),
    .Y(_01965_));
 sky130_fd_sc_hd__buf_1 _26046_ (.A(_18990_),
    .X(_04770_));
 sky130_fd_sc_hd__and2_2 _26047_ (.A(_04710_),
    .B(_18126_),
    .X(_04771_));
 sky130_fd_sc_hd__a221oi_2 _26048_ (.A1(\count_instr[53] ),
    .A2(_04757_),
    .B1(\count_instr[21] ),
    .B2(_04770_),
    .C1(_04771_),
    .Y(_01966_));
 sky130_fd_sc_hd__buf_1 _26049_ (.A(_04462_),
    .X(_04772_));
 sky130_fd_sc_hd__buf_1 _26050_ (.A(_04476_),
    .X(_04773_));
 sky130_fd_sc_hd__and2_2 _26051_ (.A(_04712_),
    .B(\timer[21] ),
    .X(_04774_));
 sky130_fd_sc_hd__a221oi_2 _26052_ (.A1(_17146_),
    .A2(_04772_),
    .B1(\cpuregs_rs1[21] ),
    .B2(_04773_),
    .C1(_04774_),
    .Y(_01968_));
 sky130_fd_sc_hd__buf_1 _26053_ (.A(_19625_),
    .X(_04775_));
 sky130_fd_sc_hd__a2bb2oi_2 _26054_ (.A1_N(_01969_),
    .A2_N(_04619_),
    .B1(_04775_),
    .B2(_01964_),
    .Y(_04776_));
 sky130_fd_sc_hd__nor2_2 _26055_ (.A(\reg_pc[21] ),
    .B(_19483_),
    .Y(_04777_));
 sky130_fd_sc_hd__and2_2 _26056_ (.A(\reg_pc[21] ),
    .B(\decoded_imm[21] ),
    .X(_04778_));
 sky130_fd_sc_hd__nor2_2 _26057_ (.A(_04777_),
    .B(_04778_),
    .Y(_04779_));
 sky130_fd_sc_hd__a21bo_2 _26058_ (.A1(_04768_),
    .A2(_04762_),
    .B1_N(_04779_),
    .X(_04780_));
 sky130_fd_sc_hd__nand3b_2 _26059_ (.A_N(_04779_),
    .B(_04768_),
    .C(_04762_),
    .Y(_04781_));
 sky130_fd_sc_hd__nand3_2 _26060_ (.A(_04780_),
    .B(_04767_),
    .C(_04781_),
    .Y(_04782_));
 sky130_fd_sc_hd__o211ai_2 _26061_ (.A1(_04618_),
    .A2(_01963_),
    .B1(_04776_),
    .C1(_04782_),
    .Y(_01970_));
 sky130_fd_sc_hd__nand3_2 _26062_ (.A(_04755_),
    .B(_04756_),
    .C(mem_rdata[22]),
    .Y(_01971_));
 sky130_vsdinv _26063_ (.A(_18217_),
    .Y(_01974_));
 sky130_fd_sc_hd__and2_2 _26064_ (.A(_04710_),
    .B(_18129_),
    .X(_04783_));
 sky130_fd_sc_hd__a221oi_2 _26065_ (.A1(_17666_),
    .A2(_04757_),
    .B1(\count_instr[22] ),
    .B2(_04770_),
    .C1(_04783_),
    .Y(_01975_));
 sky130_fd_sc_hd__buf_1 _26066_ (.A(_17022_),
    .X(_04784_));
 sky130_fd_sc_hd__and2_2 _26067_ (.A(_04784_),
    .B(\timer[22] ),
    .X(_04785_));
 sky130_fd_sc_hd__a221oi_2 _26068_ (.A1(_17143_),
    .A2(_04772_),
    .B1(\cpuregs_rs1[22] ),
    .B2(_04773_),
    .C1(_04785_),
    .Y(_01977_));
 sky130_fd_sc_hd__buf_1 _26069_ (.A(_17384_),
    .X(_04786_));
 sky130_fd_sc_hd__buf_1 _26070_ (.A(_04469_),
    .X(_04787_));
 sky130_fd_sc_hd__a2bb2oi_2 _26071_ (.A1_N(_01978_),
    .A2_N(_04787_),
    .B1(_04775_),
    .B2(_01973_),
    .Y(_04788_));
 sky130_fd_sc_hd__and2_2 _26072_ (.A(\reg_pc[22] ),
    .B(_04146_),
    .X(_04789_));
 sky130_vsdinv _26073_ (.A(_04789_),
    .Y(_04790_));
 sky130_fd_sc_hd__nand2_2 _26074_ (.A(_17498_),
    .B(_19487_),
    .Y(_04791_));
 sky130_fd_sc_hd__a21oi_2 _26075_ (.A1(_04765_),
    .A2(_04763_),
    .B1(_04761_),
    .Y(_04792_));
 sky130_fd_sc_hd__o21bai_2 _26076_ (.A1(_04777_),
    .A2(_04792_),
    .B1_N(_04778_),
    .Y(_04793_));
 sky130_fd_sc_hd__a21o_2 _26077_ (.A1(_04790_),
    .A2(_04791_),
    .B1(_04793_),
    .X(_04794_));
 sky130_fd_sc_hd__nand3_2 _26078_ (.A(_04793_),
    .B(_04790_),
    .C(_04791_),
    .Y(_04795_));
 sky130_fd_sc_hd__nand3_2 _26079_ (.A(_04794_),
    .B(_04767_),
    .C(_04795_),
    .Y(_04796_));
 sky130_fd_sc_hd__o211ai_2 _26080_ (.A1(_04786_),
    .A2(_01972_),
    .B1(_04788_),
    .C1(_04796_),
    .Y(_01979_));
 sky130_fd_sc_hd__nand3_2 _26081_ (.A(_04755_),
    .B(_04756_),
    .C(mem_rdata[23]),
    .Y(_01980_));
 sky130_vsdinv _26082_ (.A(\count_cycle[23] ),
    .Y(_01983_));
 sky130_fd_sc_hd__and2_2 _26083_ (.A(\count_instr[55] ),
    .B(_04682_),
    .X(_04797_));
 sky130_fd_sc_hd__a221oi_2 _26084_ (.A1(\count_instr[23] ),
    .A2(_04601_),
    .B1(_04719_),
    .B2(\count_cycle[55] ),
    .C1(_04797_),
    .Y(_01984_));
 sky130_fd_sc_hd__and2_2 _26085_ (.A(_17896_),
    .B(_04693_),
    .X(_04798_));
 sky130_fd_sc_hd__a221oi_2 _26086_ (.A1(_04733_),
    .A2(_04132_),
    .B1(\cpuregs_rs1[23] ),
    .B2(_04773_),
    .C1(_04798_),
    .Y(_01986_));
 sky130_fd_sc_hd__a2bb2oi_2 _26087_ (.A1_N(_01987_),
    .A2_N(_04787_),
    .B1(_04775_),
    .B2(_01982_),
    .Y(_04799_));
 sky130_fd_sc_hd__nor2_2 _26088_ (.A(\reg_pc[23] ),
    .B(_19489_),
    .Y(_04800_));
 sky130_fd_sc_hd__and2_2 _26089_ (.A(\reg_pc[23] ),
    .B(\decoded_imm[23] ),
    .X(_04801_));
 sky130_fd_sc_hd__nor2_2 _26090_ (.A(_04800_),
    .B(_04801_),
    .Y(_04802_));
 sky130_fd_sc_hd__a21bo_2 _26091_ (.A1(_04795_),
    .A2(_04790_),
    .B1_N(_04802_),
    .X(_04803_));
 sky130_fd_sc_hd__nand3b_2 _26092_ (.A_N(_04802_),
    .B(_04795_),
    .C(_04790_),
    .Y(_04804_));
 sky130_fd_sc_hd__nand3_2 _26093_ (.A(_04803_),
    .B(_04767_),
    .C(_04804_),
    .Y(_04805_));
 sky130_fd_sc_hd__o211ai_2 _26094_ (.A1(_04786_),
    .A2(_01981_),
    .B1(_04799_),
    .C1(_04805_),
    .Y(_01988_));
 sky130_fd_sc_hd__buf_1 _26095_ (.A(_04706_),
    .X(_04806_));
 sky130_fd_sc_hd__buf_1 _26096_ (.A(_04708_),
    .X(_04807_));
 sky130_fd_sc_hd__nand3_2 _26097_ (.A(_04806_),
    .B(_04807_),
    .C(mem_rdata[24]),
    .Y(_01989_));
 sky130_vsdinv _26098_ (.A(_18210_),
    .Y(_01992_));
 sky130_fd_sc_hd__buf_1 _26099_ (.A(instr_rdcycleh),
    .X(_04808_));
 sky130_fd_sc_hd__and2_2 _26100_ (.A(_04808_),
    .B(_18070_),
    .X(_04809_));
 sky130_fd_sc_hd__a221oi_2 _26101_ (.A1(_17659_),
    .A2(_04757_),
    .B1(\count_instr[24] ),
    .B2(_04770_),
    .C1(_04809_),
    .Y(_01993_));
 sky130_fd_sc_hd__buf_1 _26102_ (.A(_04479_),
    .X(_04810_));
 sky130_fd_sc_hd__and2_2 _26103_ (.A(_17134_),
    .B(_04810_),
    .X(_04811_));
 sky130_fd_sc_hd__a221oi_2 _26104_ (.A1(_04733_),
    .A2(\timer[24] ),
    .B1(\cpuregs_rs1[24] ),
    .B2(_04773_),
    .C1(_04811_),
    .Y(_01995_));
 sky130_fd_sc_hd__xor2_2 _26105_ (.A(_17489_),
    .B(\decoded_imm[24] ),
    .X(_04812_));
 sky130_fd_sc_hd__or3b_2 _26106_ (.A(_04801_),
    .B(_04812_),
    .C_N(_04803_),
    .X(_04813_));
 sky130_fd_sc_hd__a21oi_2 _26107_ (.A1(_04793_),
    .A2(_04791_),
    .B1(_04789_),
    .Y(_04814_));
 sky130_fd_sc_hd__o21bai_2 _26108_ (.A1(_04800_),
    .A2(_04814_),
    .B1_N(_04801_),
    .Y(_04815_));
 sky130_fd_sc_hd__nand2_2 _26109_ (.A(_04815_),
    .B(_04812_),
    .Y(_04816_));
 sky130_fd_sc_hd__and2b_2 _26110_ (.A_N(_01990_),
    .B(_04678_),
    .X(_04817_));
 sky130_fd_sc_hd__o2bb2ai_2 _26111_ (.A1_N(_04704_),
    .A2_N(_01991_),
    .B1(_01996_),
    .B2(_04680_),
    .Y(_04818_));
 sky130_fd_sc_hd__a311o_2 _26112_ (.A1(_04813_),
    .A2(_04816_),
    .A3(_04702_),
    .B1(_04817_),
    .C1(_04818_),
    .X(_01997_));
 sky130_fd_sc_hd__nand3_2 _26113_ (.A(_04806_),
    .B(_04807_),
    .C(mem_rdata[25]),
    .Y(_01998_));
 sky130_vsdinv _26114_ (.A(_18211_),
    .Y(_02001_));
 sky130_fd_sc_hd__buf_1 _26115_ (.A(_04510_),
    .X(_04819_));
 sky130_fd_sc_hd__and2_2 _26116_ (.A(_04808_),
    .B(_18091_),
    .X(_04820_));
 sky130_fd_sc_hd__a221oi_2 _26117_ (.A1(\count_instr[57] ),
    .A2(_04819_),
    .B1(_17772_),
    .B2(_04770_),
    .C1(_04820_),
    .Y(_02002_));
 sky130_fd_sc_hd__buf_1 _26118_ (.A(_04476_),
    .X(_04821_));
 sky130_fd_sc_hd__and2_2 _26119_ (.A(_04784_),
    .B(\timer[25] ),
    .X(_04822_));
 sky130_fd_sc_hd__a221oi_2 _26120_ (.A1(_17129_),
    .A2(_04772_),
    .B1(\cpuregs_rs1[25] ),
    .B2(_04821_),
    .C1(_04822_),
    .Y(_02004_));
 sky130_fd_sc_hd__and2_2 _26121_ (.A(\reg_pc[24] ),
    .B(\decoded_imm[24] ),
    .X(_04823_));
 sky130_fd_sc_hd__nor2_2 _26122_ (.A(_17483_),
    .B(\decoded_imm[25] ),
    .Y(_04824_));
 sky130_fd_sc_hd__and2_2 _26123_ (.A(\reg_pc[25] ),
    .B(\decoded_imm[25] ),
    .X(_04825_));
 sky130_fd_sc_hd__nor2_2 _26124_ (.A(_04824_),
    .B(_04825_),
    .Y(_04826_));
 sky130_fd_sc_hd__a211oi_2 _26125_ (.A1(_04815_),
    .A2(_04812_),
    .B1(_04823_),
    .C1(_04826_),
    .Y(_04827_));
 sky130_vsdinv _26126_ (.A(_04823_),
    .Y(_04828_));
 sky130_fd_sc_hd__a21boi_2 _26127_ (.A1(_04816_),
    .A2(_04828_),
    .B1_N(_04826_),
    .Y(_04829_));
 sky130_fd_sc_hd__or2b_2 _26128_ (.A(_01999_),
    .B_N(_04556_),
    .X(_04830_));
 sky130_fd_sc_hd__a2bb2oi_2 _26129_ (.A1_N(_02005_),
    .A2_N(_04540_),
    .B1(_04581_),
    .B2(_02000_),
    .Y(_04831_));
 sky130_fd_sc_hd__o311ai_2 _26130_ (.A1(_04482_),
    .A2(_04827_),
    .A3(_04829_),
    .B1(_04830_),
    .C1(_04831_),
    .Y(_02006_));
 sky130_fd_sc_hd__nand3_2 _26131_ (.A(_04806_),
    .B(_04807_),
    .C(mem_rdata[26]),
    .Y(_02007_));
 sky130_vsdinv _26132_ (.A(_18208_),
    .Y(_02010_));
 sky130_fd_sc_hd__and2_2 _26133_ (.A(_04808_),
    .B(_18117_),
    .X(_04832_));
 sky130_fd_sc_hd__a221oi_2 _26134_ (.A1(\count_instr[58] ),
    .A2(_04819_),
    .B1(_17767_),
    .B2(_04460_),
    .C1(_04832_),
    .Y(_02011_));
 sky130_fd_sc_hd__and2_2 _26135_ (.A(_17126_),
    .B(_04810_),
    .X(_04833_));
 sky130_fd_sc_hd__a221oi_2 _26136_ (.A1(_04464_),
    .A2(\timer[26] ),
    .B1(\cpuregs_rs1[26] ),
    .B2(_04821_),
    .C1(_04833_),
    .Y(_02013_));
 sky130_fd_sc_hd__and2_2 _26137_ (.A(_04812_),
    .B(_04826_),
    .X(_04834_));
 sky130_fd_sc_hd__xor2_2 _26138_ (.A(\reg_pc[26] ),
    .B(\decoded_imm[26] ),
    .X(_04835_));
 sky130_fd_sc_hd__o21bai_2 _26139_ (.A1(_04824_),
    .A2(_04828_),
    .B1_N(_04825_),
    .Y(_04836_));
 sky130_fd_sc_hd__a211oi_2 _26140_ (.A1(_04815_),
    .A2(_04834_),
    .B1(_04835_),
    .C1(_04836_),
    .Y(_04837_));
 sky130_vsdinv _26141_ (.A(_04835_),
    .Y(_04838_));
 sky130_fd_sc_hd__a21oi_2 _26142_ (.A1(_04815_),
    .A2(_04834_),
    .B1(_04836_),
    .Y(_04839_));
 sky130_fd_sc_hd__nor2_2 _26143_ (.A(_04838_),
    .B(_04839_),
    .Y(_04840_));
 sky130_fd_sc_hd__nand2_2 _26144_ (.A(_19661_),
    .B(_02009_),
    .Y(_04841_));
 sky130_fd_sc_hd__o221a_2 _26145_ (.A1(_02008_),
    .A2(_16823_),
    .B1(_04469_),
    .B2(_02014_),
    .C1(_04841_),
    .X(_04842_));
 sky130_fd_sc_hd__o31ai_2 _26146_ (.A1(_04633_),
    .A2(_04837_),
    .A3(_04840_),
    .B1(_04842_),
    .Y(_02015_));
 sky130_fd_sc_hd__nand3_2 _26147_ (.A(_04806_),
    .B(_04807_),
    .C(mem_rdata[27]),
    .Y(_02016_));
 sky130_vsdinv _26148_ (.A(_18205_),
    .Y(_02019_));
 sky130_fd_sc_hd__and2_2 _26149_ (.A(_04808_),
    .B(_18073_),
    .X(_04843_));
 sky130_fd_sc_hd__a221oi_2 _26150_ (.A1(_17648_),
    .A2(_04819_),
    .B1(_17763_),
    .B2(_04460_),
    .C1(_04843_),
    .Y(_02020_));
 sky130_fd_sc_hd__and2_2 _26151_ (.A(_04784_),
    .B(\timer[27] ),
    .X(_04844_));
 sky130_fd_sc_hd__a221oi_2 _26152_ (.A1(\irq_mask[27] ),
    .A2(_04772_),
    .B1(\cpuregs_rs1[27] ),
    .B2(_04821_),
    .C1(_04844_),
    .Y(_02022_));
 sky130_fd_sc_hd__and2_2 _26153_ (.A(\reg_pc[26] ),
    .B(\decoded_imm[26] ),
    .X(_04845_));
 sky130_fd_sc_hd__nor2_2 _26154_ (.A(\reg_pc[27] ),
    .B(\decoded_imm[27] ),
    .Y(_04846_));
 sky130_fd_sc_hd__and2_2 _26155_ (.A(\reg_pc[27] ),
    .B(\decoded_imm[27] ),
    .X(_04847_));
 sky130_fd_sc_hd__nor2_2 _26156_ (.A(_04846_),
    .B(_04847_),
    .Y(_04848_));
 sky130_fd_sc_hd__o21ai_2 _26157_ (.A1(_04845_),
    .A2(_04840_),
    .B1(_04848_),
    .Y(_04849_));
 sky130_vsdinv _26158_ (.A(_04845_),
    .Y(_04850_));
 sky130_fd_sc_hd__o221ai_2 _26159_ (.A1(_04847_),
    .A2(_04846_),
    .B1(_04838_),
    .B2(_04839_),
    .C1(_04850_),
    .Y(_04851_));
 sky130_fd_sc_hd__and2b_2 _26160_ (.A_N(_02017_),
    .B(_17389_),
    .X(_04852_));
 sky130_fd_sc_hd__o2bb2ai_2 _26161_ (.A1_N(_04704_),
    .A2_N(_02018_),
    .B1(_02023_),
    .B2(_18541_),
    .Y(_04853_));
 sky130_fd_sc_hd__a311o_2 _26162_ (.A1(_04849_),
    .A2(_04851_),
    .A3(_04702_),
    .B1(_04852_),
    .C1(_04853_),
    .X(_02024_));
 sky130_fd_sc_hd__buf_1 _26163_ (.A(_04706_),
    .X(_04854_));
 sky130_fd_sc_hd__buf_1 _26164_ (.A(_04708_),
    .X(_04855_));
 sky130_fd_sc_hd__nand3_2 _26165_ (.A(_04854_),
    .B(_04855_),
    .C(mem_rdata[28]),
    .Y(_02025_));
 sky130_vsdinv _26166_ (.A(_18202_),
    .Y(_02028_));
 sky130_fd_sc_hd__and2_2 _26167_ (.A(_04528_),
    .B(_18093_),
    .X(_04856_));
 sky130_fd_sc_hd__a221oi_2 _26168_ (.A1(_17650_),
    .A2(_04819_),
    .B1(_17760_),
    .B2(_04460_),
    .C1(_04856_),
    .Y(_02029_));
 sky130_fd_sc_hd__and2_2 _26169_ (.A(_04784_),
    .B(\timer[28] ),
    .X(_04857_));
 sky130_fd_sc_hd__a221oi_2 _26170_ (.A1(_17116_),
    .A2(_04480_),
    .B1(\cpuregs_rs1[28] ),
    .B2(_04821_),
    .C1(_04857_),
    .Y(_02031_));
 sky130_fd_sc_hd__and2_2 _26171_ (.A(\reg_pc[28] ),
    .B(\decoded_imm[28] ),
    .X(_04858_));
 sky130_fd_sc_hd__nor2_2 _26172_ (.A(\reg_pc[28] ),
    .B(\decoded_imm[28] ),
    .Y(_04859_));
 sky130_fd_sc_hd__nand2_2 _26173_ (.A(_04835_),
    .B(_04848_),
    .Y(_04860_));
 sky130_fd_sc_hd__o21ba_2 _26174_ (.A1(_04846_),
    .A2(_04850_),
    .B1_N(_04847_),
    .X(_04861_));
 sky130_fd_sc_hd__o221a_2 _26175_ (.A1(_04858_),
    .A2(_04859_),
    .B1(_04860_),
    .B2(_04839_),
    .C1(_04861_),
    .X(_04862_));
 sky130_fd_sc_hd__o21ai_2 _26176_ (.A1(_04860_),
    .A2(_04839_),
    .B1(_04861_),
    .Y(_04863_));
 sky130_fd_sc_hd__nor3b_2 _26177_ (.A(_04858_),
    .B(_04859_),
    .C_N(_04863_),
    .Y(_04864_));
 sky130_fd_sc_hd__or2b_2 _26178_ (.A(_02026_),
    .B_N(_04556_),
    .X(_04865_));
 sky130_fd_sc_hd__a2bb2oi_2 _26179_ (.A1_N(_02032_),
    .A2_N(_04540_),
    .B1(_04581_),
    .B2(_02027_),
    .Y(_04866_));
 sky130_fd_sc_hd__o311ai_2 _26180_ (.A1(_16985_),
    .A2(_04862_),
    .A3(_04864_),
    .B1(_04865_),
    .C1(_04866_),
    .Y(_02033_));
 sky130_fd_sc_hd__nand3_2 _26181_ (.A(_04854_),
    .B(_04855_),
    .C(mem_rdata[29]),
    .Y(_02034_));
 sky130_vsdinv _26182_ (.A(_18203_),
    .Y(_02037_));
 sky130_fd_sc_hd__and2_2 _26183_ (.A(_17644_),
    .B(_04599_),
    .X(_04867_));
 sky130_fd_sc_hd__a221oi_2 _26184_ (.A1(_17757_),
    .A2(_04601_),
    .B1(_04529_),
    .B2(_18075_),
    .C1(_04867_),
    .Y(_02038_));
 sky130_fd_sc_hd__and2_2 _26185_ (.A(_17113_),
    .B(_04810_),
    .X(_04868_));
 sky130_fd_sc_hd__a221oi_2 _26186_ (.A1(_04464_),
    .A2(\timer[29] ),
    .B1(\cpuregs_rs1[29] ),
    .B2(_04477_),
    .C1(_04868_),
    .Y(_02040_));
 sky130_fd_sc_hd__a2bb2oi_2 _26187_ (.A1_N(_02041_),
    .A2_N(_04787_),
    .B1(_04775_),
    .B2(_02036_),
    .Y(_04869_));
 sky130_fd_sc_hd__and2_2 _26188_ (.A(\reg_pc[29] ),
    .B(\decoded_imm[29] ),
    .X(_04870_));
 sky130_fd_sc_hd__nor2_2 _26189_ (.A(\reg_pc[29] ),
    .B(\decoded_imm[29] ),
    .Y(_04871_));
 sky130_vsdinv _26190_ (.A(_04859_),
    .Y(_04872_));
 sky130_fd_sc_hd__a21oi_2 _26191_ (.A1(_04863_),
    .A2(_04872_),
    .B1(_04858_),
    .Y(_04873_));
 sky130_fd_sc_hd__nor3_2 _26192_ (.A(_04870_),
    .B(_04871_),
    .C(_04873_),
    .Y(_04874_));
 sky130_fd_sc_hd__o21ai_2 _26193_ (.A1(_04870_),
    .A2(_04871_),
    .B1(_04873_),
    .Y(_04875_));
 sky130_fd_sc_hd__nand3b_2 _26194_ (.A_N(_04874_),
    .B(_04467_),
    .C(_04875_),
    .Y(_04876_));
 sky130_fd_sc_hd__o211ai_2 _26195_ (.A1(_04786_),
    .A2(_02035_),
    .B1(_04869_),
    .C1(_04876_),
    .Y(_02042_));
 sky130_fd_sc_hd__nand3_2 _26196_ (.A(_04854_),
    .B(_04855_),
    .C(mem_rdata[30]),
    .Y(_02043_));
 sky130_fd_sc_hd__and2_2 _26197_ (.A(_17755_),
    .B(_18990_),
    .X(_04877_));
 sky130_fd_sc_hd__a221oi_2 _26198_ (.A1(\count_instr[62] ),
    .A2(_18987_),
    .B1(_04529_),
    .B2(\count_cycle[62] ),
    .C1(_04877_),
    .Y(_02047_));
 sky130_fd_sc_hd__and2_2 _26199_ (.A(_04513_),
    .B(\timer[30] ),
    .X(_04878_));
 sky130_fd_sc_hd__a221oi_2 _26200_ (.A1(_17108_),
    .A2(_04480_),
    .B1(\cpuregs_rs1[30] ),
    .B2(_04477_),
    .C1(_04878_),
    .Y(_02049_));
 sky130_fd_sc_hd__a2bb2oi_2 _26201_ (.A1_N(_02050_),
    .A2_N(_04787_),
    .B1(_04488_),
    .B2(_02045_),
    .Y(_04879_));
 sky130_fd_sc_hd__xor2_2 _26202_ (.A(\reg_pc[30] ),
    .B(\decoded_imm[30] ),
    .X(_04880_));
 sky130_fd_sc_hd__o21bai_2 _26203_ (.A1(_04871_),
    .A2(_04873_),
    .B1_N(_04870_),
    .Y(_04881_));
 sky130_fd_sc_hd__nor2_2 _26204_ (.A(_04880_),
    .B(_04881_),
    .Y(_04882_));
 sky130_fd_sc_hd__nand2_2 _26205_ (.A(_04881_),
    .B(_04880_),
    .Y(_04883_));
 sky130_fd_sc_hd__nand3b_2 _26206_ (.A_N(_04882_),
    .B(_04467_),
    .C(_04883_),
    .Y(_04884_));
 sky130_fd_sc_hd__o211ai_2 _26207_ (.A1(_04786_),
    .A2(_02044_),
    .B1(_04879_),
    .C1(_04884_),
    .Y(_02051_));
 sky130_fd_sc_hd__nand3_2 _26208_ (.A(_04854_),
    .B(_04855_),
    .C(mem_rdata[31]),
    .Y(_02052_));
 sky130_vsdinv _26209_ (.A(\count_cycle[31] ),
    .Y(_02055_));
 sky130_fd_sc_hd__and2_2 _26210_ (.A(\count_instr[63] ),
    .B(_04599_),
    .X(_04885_));
 sky130_fd_sc_hd__a221oi_2 _26211_ (.A1(\count_instr[31] ),
    .A2(_04601_),
    .B1(_04529_),
    .B2(\count_cycle[63] ),
    .C1(_04885_),
    .Y(_02056_));
 sky130_fd_sc_hd__and2_2 _26212_ (.A(_17088_),
    .B(_04810_),
    .X(_04886_));
 sky130_fd_sc_hd__a221oi_2 _26213_ (.A1(_04464_),
    .A2(\timer[31] ),
    .B1(\cpuregs_rs1[31] ),
    .B2(_04477_),
    .C1(_04886_),
    .Y(_02058_));
 sky130_fd_sc_hd__and2_2 _26214_ (.A(\reg_pc[30] ),
    .B(\decoded_imm[30] ),
    .X(_04887_));
 sky130_vsdinv _26215_ (.A(_04887_),
    .Y(_04888_));
 sky130_fd_sc_hd__xnor2_2 _26216_ (.A(\reg_pc[31] ),
    .B(\decoded_imm[31] ),
    .Y(_04889_));
 sky130_fd_sc_hd__a21oi_2 _26217_ (.A1(_04883_),
    .A2(_04888_),
    .B1(_04889_),
    .Y(_04890_));
 sky130_fd_sc_hd__nand3_2 _26218_ (.A(_04883_),
    .B(_04888_),
    .C(_04889_),
    .Y(_04891_));
 sky130_fd_sc_hd__nand2_2 _26219_ (.A(_04891_),
    .B(_04589_),
    .Y(_04892_));
 sky130_fd_sc_hd__nand2_2 _26220_ (.A(_18003_),
    .B(_02054_),
    .Y(_04893_));
 sky130_fd_sc_hd__o221ai_2 _26221_ (.A1(_02053_),
    .A2(_17384_),
    .B1(_02059_),
    .B2(_18541_),
    .C1(_04893_),
    .Y(_04894_));
 sky130_fd_sc_hd__o21bai_2 _26222_ (.A1(_04890_),
    .A2(_04892_),
    .B1_N(_04894_),
    .Y(_02060_));
 sky130_fd_sc_hd__nand3b_2 _26223_ (.A_N(\decoded_rd[4] ),
    .B(_17051_),
    .C(_18022_),
    .Y(_02061_));
 sky130_fd_sc_hd__o21bai_2 _26224_ (.A1(_02064_),
    .A2(_19771_),
    .B1_N(_19773_),
    .Y(_02065_));
 sky130_fd_sc_hd__o2111a_2 _26225_ (.A1(_18014_),
    .A2(_18019_),
    .B1(_18022_),
    .C1(_00309_),
    .D1(_17051_),
    .X(_02066_));
 sky130_vsdinv _26226_ (.A(_17029_),
    .Y(_02067_));
 sky130_fd_sc_hd__and2_2 _26227_ (.A(_16981_),
    .B(_00343_),
    .X(_04895_));
 sky130_fd_sc_hd__o21ai_2 _26228_ (.A1(_19771_),
    .A2(_04895_),
    .B1(_19037_),
    .Y(_02068_));
 sky130_fd_sc_hd__buf_1 _26229_ (.A(_17034_),
    .X(_04896_));
 sky130_fd_sc_hd__and2b_2 _26230_ (.A_N(latched_branch),
    .B(_16987_),
    .X(_04897_));
 sky130_fd_sc_hd__buf_1 _26231_ (.A(_04897_),
    .X(_04898_));
 sky130_fd_sc_hd__buf_1 _26232_ (.A(_04898_),
    .X(_04899_));
 sky130_fd_sc_hd__nor3_2 _26233_ (.A(_04896_),
    .B(_04293_),
    .C(_04899_),
    .Y(_02069_));
 sky130_fd_sc_hd__buf_1 _26234_ (.A(_04898_),
    .X(_04900_));
 sky130_fd_sc_hd__and2_2 _26235_ (.A(_04292_),
    .B(_19382_),
    .X(_04901_));
 sky130_fd_sc_hd__a221o_2 _26236_ (.A1(_16888_),
    .A2(_04896_),
    .B1(_04900_),
    .B2(_02070_),
    .C1(_04901_),
    .X(_02071_));
 sky130_fd_sc_hd__and2_2 _26237_ (.A(_04292_),
    .B(\reg_next_pc[1] ),
    .X(_04902_));
 sky130_fd_sc_hd__a221o_2 _26238_ (.A1(_16890_),
    .A2(_04896_),
    .B1(_04900_),
    .B2(_01465_),
    .C1(_04902_),
    .X(_02072_));
 sky130_vsdinv _26239_ (.A(_17591_),
    .Y(_02073_));
 sky130_fd_sc_hd__buf_1 _26240_ (.A(_04897_),
    .X(_04903_));
 sky130_fd_sc_hd__buf_1 _26241_ (.A(_17033_),
    .X(_04904_));
 sky130_fd_sc_hd__nand3b_2 _26242_ (.A_N(_17989_),
    .B(_04904_),
    .C(_17991_),
    .Y(_04905_));
 sky130_vsdinv _26243_ (.A(_04905_),
    .Y(_04906_));
 sky130_fd_sc_hd__a221o_2 _26244_ (.A1(_04293_),
    .A2(\reg_next_pc[2] ),
    .B1(_00293_),
    .B2(_04903_),
    .C1(_04906_),
    .X(_02074_));
 sky130_fd_sc_hd__xor2_2 _26245_ (.A(_17585_),
    .B(_17591_),
    .X(_02075_));
 sky130_fd_sc_hd__buf_1 _26246_ (.A(\irq_state[0] ),
    .X(_04907_));
 sky130_fd_sc_hd__buf_1 _26247_ (.A(_04907_),
    .X(_04908_));
 sky130_fd_sc_hd__and2_2 _26248_ (.A(_04908_),
    .B(\reg_next_pc[3] ),
    .X(_04909_));
 sky130_fd_sc_hd__a221o_2 _26249_ (.A1(_16889_),
    .A2(_04896_),
    .B1(_04900_),
    .B2(_01468_),
    .C1(_04909_),
    .X(_02076_));
 sky130_fd_sc_hd__nand2_2 _26250_ (.A(_17585_),
    .B(_17590_),
    .Y(_04910_));
 sky130_fd_sc_hd__xnor2_2 _26251_ (.A(_17581_),
    .B(_04910_),
    .Y(_02077_));
 sky130_fd_sc_hd__buf_1 _26252_ (.A(_04904_),
    .X(_04911_));
 sky130_fd_sc_hd__and2_2 _26253_ (.A(_04908_),
    .B(\reg_next_pc[4] ),
    .X(_04912_));
 sky130_fd_sc_hd__a221o_2 _26254_ (.A1(_16898_),
    .A2(_04911_),
    .B1(_04900_),
    .B2(_01472_),
    .C1(_04912_),
    .X(_02078_));
 sky130_fd_sc_hd__nand3_2 _26255_ (.A(_17581_),
    .B(_17584_),
    .C(_17590_),
    .Y(_04913_));
 sky130_fd_sc_hd__xnor2_2 _26256_ (.A(_17575_),
    .B(_04913_),
    .Y(_02079_));
 sky130_fd_sc_hd__buf_1 _26257_ (.A(_04898_),
    .X(_04914_));
 sky130_fd_sc_hd__and2_2 _26258_ (.A(_04908_),
    .B(\reg_next_pc[5] ),
    .X(_04915_));
 sky130_fd_sc_hd__a221o_2 _26259_ (.A1(_16900_),
    .A2(_04911_),
    .B1(_04914_),
    .B2(_01476_),
    .C1(_04915_),
    .X(_02080_));
 sky130_fd_sc_hd__and4_2 _26260_ (.A(_17574_),
    .B(_17580_),
    .C(_17584_),
    .D(_17590_),
    .X(_04916_));
 sky130_fd_sc_hd__xor2_2 _26261_ (.A(_17571_),
    .B(_04916_),
    .X(_02081_));
 sky130_fd_sc_hd__and2_2 _26262_ (.A(_04908_),
    .B(\reg_next_pc[6] ),
    .X(_04917_));
 sky130_fd_sc_hd__a221o_2 _26263_ (.A1(_16899_),
    .A2(_04911_),
    .B1(_04914_),
    .B2(_01479_),
    .C1(_04917_),
    .X(_02082_));
 sky130_fd_sc_hd__nand3b_2 _26264_ (.A_N(_04913_),
    .B(_17571_),
    .C(_17575_),
    .Y(_04918_));
 sky130_fd_sc_hd__xnor2_2 _26265_ (.A(_17567_),
    .B(_04918_),
    .Y(_02083_));
 sky130_fd_sc_hd__a32o_2 _26266_ (.A1(_16897_),
    .A2(_17035_),
    .A3(_17968_),
    .B1(_19772_),
    .B2(\reg_next_pc[7] ),
    .X(_04919_));
 sky130_fd_sc_hd__a21o_2 _26267_ (.A1(_01482_),
    .A2(_04899_),
    .B1(_04919_),
    .X(_02084_));
 sky130_fd_sc_hd__nand3_2 _26268_ (.A(_04916_),
    .B(_17567_),
    .C(\reg_pc[6] ),
    .Y(_04920_));
 sky130_fd_sc_hd__xor2_2 _26269_ (.A(_17565_),
    .B(_04920_),
    .X(_02085_));
 sky130_fd_sc_hd__buf_1 _26270_ (.A(_04907_),
    .X(_04921_));
 sky130_fd_sc_hd__and2_2 _26271_ (.A(_04921_),
    .B(\reg_next_pc[8] ),
    .X(_04922_));
 sky130_fd_sc_hd__a221o_2 _26272_ (.A1(_16883_),
    .A2(_04911_),
    .B1(_04914_),
    .B2(_01485_),
    .C1(_04922_),
    .X(_02086_));
 sky130_fd_sc_hd__nor2_2 _26273_ (.A(_17565_),
    .B(_04920_),
    .Y(_04923_));
 sky130_fd_sc_hd__xor2_2 _26274_ (.A(_17558_),
    .B(_04923_),
    .X(_02087_));
 sky130_fd_sc_hd__buf_1 _26275_ (.A(_17033_),
    .X(_04924_));
 sky130_fd_sc_hd__buf_1 _26276_ (.A(_04924_),
    .X(_04925_));
 sky130_fd_sc_hd__and2_2 _26277_ (.A(_04921_),
    .B(\reg_next_pc[9] ),
    .X(_04926_));
 sky130_fd_sc_hd__a221o_2 _26278_ (.A1(_16885_),
    .A2(_04925_),
    .B1(_04914_),
    .B2(_01488_),
    .C1(_04926_),
    .X(_02088_));
 sky130_fd_sc_hd__nor3b_2 _26279_ (.A(_17565_),
    .B(_04920_),
    .C_N(_17557_),
    .Y(_04927_));
 sky130_fd_sc_hd__xor2_2 _26280_ (.A(_17553_),
    .B(_04927_),
    .X(_02089_));
 sky130_fd_sc_hd__buf_1 _26281_ (.A(_04897_),
    .X(_04928_));
 sky130_fd_sc_hd__buf_1 _26282_ (.A(_04928_),
    .X(_04929_));
 sky130_fd_sc_hd__and2_2 _26283_ (.A(_04921_),
    .B(\reg_next_pc[10] ),
    .X(_04930_));
 sky130_fd_sc_hd__a221o_2 _26284_ (.A1(_16884_),
    .A2(_04925_),
    .B1(_04929_),
    .B2(_01491_),
    .C1(_04930_),
    .X(_02090_));
 sky130_fd_sc_hd__nand3_2 _26285_ (.A(_04923_),
    .B(_17553_),
    .C(_17558_),
    .Y(_04931_));
 sky130_fd_sc_hd__xnor2_2 _26286_ (.A(_17549_),
    .B(_04931_),
    .Y(_02091_));
 sky130_fd_sc_hd__a32o_2 _26287_ (.A1(_16882_),
    .A2(_17035_),
    .A3(_17951_),
    .B1(_19772_),
    .B2(\reg_next_pc[11] ),
    .X(_04932_));
 sky130_fd_sc_hd__a21o_2 _26288_ (.A1(_01494_),
    .A2(_04899_),
    .B1(_04932_),
    .X(_02092_));
 sky130_fd_sc_hd__nand3_2 _26289_ (.A(_04927_),
    .B(\reg_pc[11] ),
    .C(_17552_),
    .Y(_04933_));
 sky130_fd_sc_hd__xor2_2 _26290_ (.A(_17546_),
    .B(_04933_),
    .X(_02093_));
 sky130_fd_sc_hd__and2_2 _26291_ (.A(_04921_),
    .B(\reg_next_pc[12] ),
    .X(_04934_));
 sky130_fd_sc_hd__a221o_2 _26292_ (.A1(_16920_),
    .A2(_04925_),
    .B1(_04929_),
    .B2(_01497_),
    .C1(_04934_),
    .X(_02094_));
 sky130_fd_sc_hd__nor2_2 _26293_ (.A(_17546_),
    .B(_04933_),
    .Y(_04935_));
 sky130_fd_sc_hd__xor2_2 _26294_ (.A(_17539_),
    .B(_04935_),
    .X(_02095_));
 sky130_fd_sc_hd__buf_1 _26295_ (.A(_04907_),
    .X(_04936_));
 sky130_fd_sc_hd__and2_2 _26296_ (.A(_04936_),
    .B(\reg_next_pc[13] ),
    .X(_04937_));
 sky130_fd_sc_hd__a221o_2 _26297_ (.A1(_16922_),
    .A2(_04925_),
    .B1(_04929_),
    .B2(_01500_),
    .C1(_04937_),
    .X(_02096_));
 sky130_fd_sc_hd__nor3b_2 _26298_ (.A(_17546_),
    .B(_04933_),
    .C_N(_17538_),
    .Y(_04938_));
 sky130_fd_sc_hd__xor2_2 _26299_ (.A(_17536_),
    .B(_04938_),
    .X(_02097_));
 sky130_fd_sc_hd__buf_1 _26300_ (.A(_04924_),
    .X(_04939_));
 sky130_fd_sc_hd__and2_2 _26301_ (.A(_04936_),
    .B(\reg_next_pc[14] ),
    .X(_04940_));
 sky130_fd_sc_hd__a221o_2 _26302_ (.A1(_16921_),
    .A2(_04939_),
    .B1(_04929_),
    .B2(_01503_),
    .C1(_04940_),
    .X(_02098_));
 sky130_fd_sc_hd__nand3_2 _26303_ (.A(_04935_),
    .B(_17536_),
    .C(_17539_),
    .Y(_04941_));
 sky130_fd_sc_hd__xnor2_2 _26304_ (.A(_17530_),
    .B(_04941_),
    .Y(_02099_));
 sky130_fd_sc_hd__nand3b_2 _26305_ (.A_N(_17931_),
    .B(_04904_),
    .C(_17933_),
    .Y(_04942_));
 sky130_vsdinv _26306_ (.A(_04942_),
    .Y(_04943_));
 sky130_fd_sc_hd__a221o_2 _26307_ (.A1(_04293_),
    .A2(\reg_next_pc[15] ),
    .B1(_01506_),
    .B2(_04903_),
    .C1(_04943_),
    .X(_02100_));
 sky130_vsdinv _26308_ (.A(_17526_),
    .Y(_04944_));
 sky130_fd_sc_hd__nand3_2 _26309_ (.A(_04938_),
    .B(_17529_),
    .C(_17535_),
    .Y(_04945_));
 sky130_fd_sc_hd__xor2_2 _26310_ (.A(_04944_),
    .B(_04945_),
    .X(_02101_));
 sky130_fd_sc_hd__buf_1 _26311_ (.A(_04928_),
    .X(_04946_));
 sky130_fd_sc_hd__and2_2 _26312_ (.A(_04936_),
    .B(\reg_next_pc[16] ),
    .X(_04947_));
 sky130_fd_sc_hd__a221o_2 _26313_ (.A1(_16903_),
    .A2(_04939_),
    .B1(_04946_),
    .B2(_01509_),
    .C1(_04947_),
    .X(_02102_));
 sky130_fd_sc_hd__nor2_2 _26314_ (.A(_04944_),
    .B(_04945_),
    .Y(_04948_));
 sky130_fd_sc_hd__xor2_2 _26315_ (.A(_17524_),
    .B(_04948_),
    .X(_02103_));
 sky130_fd_sc_hd__and2_2 _26316_ (.A(_04936_),
    .B(\reg_next_pc[17] ),
    .X(_04949_));
 sky130_fd_sc_hd__a221o_2 _26317_ (.A1(_16906_),
    .A2(_04939_),
    .B1(_04946_),
    .B2(_01512_),
    .C1(_04949_),
    .X(_02104_));
 sky130_fd_sc_hd__and4_2 _26318_ (.A(_04923_),
    .B(_17549_),
    .C(_17552_),
    .D(_17557_),
    .X(_04950_));
 sky130_fd_sc_hd__and4_2 _26319_ (.A(_04950_),
    .B(_17535_),
    .C(_17538_),
    .D(_17545_),
    .X(_04951_));
 sky130_fd_sc_hd__and4_2 _26320_ (.A(_04951_),
    .B(_17523_),
    .C(_17526_),
    .D(_17530_),
    .X(_04952_));
 sky130_fd_sc_hd__xor2_2 _26321_ (.A(_17516_),
    .B(_04952_),
    .X(_02105_));
 sky130_fd_sc_hd__buf_1 _26322_ (.A(_04907_),
    .X(_04953_));
 sky130_fd_sc_hd__and2_2 _26323_ (.A(_04953_),
    .B(\reg_next_pc[18] ),
    .X(_04954_));
 sky130_fd_sc_hd__a221o_2 _26324_ (.A1(_16904_),
    .A2(_04939_),
    .B1(_04946_),
    .B2(_01515_),
    .C1(_04954_),
    .X(_02106_));
 sky130_fd_sc_hd__nand3_2 _26325_ (.A(_04948_),
    .B(_17516_),
    .C(_17524_),
    .Y(_04955_));
 sky130_fd_sc_hd__xnor2_2 _26326_ (.A(_17510_),
    .B(_04955_),
    .Y(_02107_));
 sky130_fd_sc_hd__buf_1 _26327_ (.A(_04924_),
    .X(_04956_));
 sky130_fd_sc_hd__and2_2 _26328_ (.A(_04953_),
    .B(\reg_next_pc[19] ),
    .X(_04957_));
 sky130_fd_sc_hd__a221o_2 _26329_ (.A1(_16905_),
    .A2(_04956_),
    .B1(_04946_),
    .B2(_01518_),
    .C1(_04957_),
    .X(_02108_));
 sky130_fd_sc_hd__and4_2 _26330_ (.A(_04948_),
    .B(_17509_),
    .C(_17515_),
    .D(_17523_),
    .X(_04958_));
 sky130_fd_sc_hd__xor2_2 _26331_ (.A(_04233_),
    .B(_04958_),
    .X(_02109_));
 sky130_fd_sc_hd__buf_1 _26332_ (.A(_04928_),
    .X(_04959_));
 sky130_fd_sc_hd__and2_2 _26333_ (.A(_04953_),
    .B(\reg_next_pc[20] ),
    .X(_04960_));
 sky130_fd_sc_hd__a221o_2 _26334_ (.A1(_16893_),
    .A2(_04956_),
    .B1(_04959_),
    .B2(_01521_),
    .C1(_04960_),
    .X(_02110_));
 sky130_fd_sc_hd__and4_2 _26335_ (.A(_04952_),
    .B(_04233_),
    .C(_17510_),
    .D(_17515_),
    .X(_04961_));
 sky130_fd_sc_hd__xor2_2 _26336_ (.A(_17503_),
    .B(_04961_),
    .X(_02111_));
 sky130_fd_sc_hd__and2_2 _26337_ (.A(_04953_),
    .B(\reg_next_pc[21] ),
    .X(_04962_));
 sky130_fd_sc_hd__a221o_2 _26338_ (.A1(_16895_),
    .A2(_04956_),
    .B1(_04959_),
    .B2(_01524_),
    .C1(_04962_),
    .X(_02112_));
 sky130_fd_sc_hd__and4_2 _26339_ (.A(_04935_),
    .B(_17529_),
    .C(_17535_),
    .D(_17538_),
    .X(_04963_));
 sky130_fd_sc_hd__and4_2 _26340_ (.A(_04963_),
    .B(_17515_),
    .C(_17523_),
    .D(\reg_pc[16] ),
    .X(_04964_));
 sky130_fd_sc_hd__and4_2 _26341_ (.A(_04964_),
    .B(\reg_pc[21] ),
    .C(\reg_pc[20] ),
    .D(_17509_),
    .X(_04965_));
 sky130_fd_sc_hd__xor2_2 _26342_ (.A(_04240_),
    .B(_04965_),
    .X(_02113_));
 sky130_fd_sc_hd__buf_1 _26343_ (.A(_17036_),
    .X(_04966_));
 sky130_fd_sc_hd__and2_2 _26344_ (.A(_04966_),
    .B(\reg_next_pc[22] ),
    .X(_04967_));
 sky130_fd_sc_hd__a221o_2 _26345_ (.A1(_16894_),
    .A2(_04956_),
    .B1(_04959_),
    .B2(_01527_),
    .C1(_04967_),
    .X(_02114_));
 sky130_fd_sc_hd__and4_2 _26346_ (.A(_04958_),
    .B(_04240_),
    .C(_17503_),
    .D(_04233_),
    .X(_04968_));
 sky130_fd_sc_hd__xor2_2 _26347_ (.A(_17492_),
    .B(_04968_),
    .X(_02115_));
 sky130_fd_sc_hd__nand3b_2 _26348_ (.A_N(_17896_),
    .B(_04904_),
    .C(_17899_),
    .Y(_04969_));
 sky130_vsdinv _26349_ (.A(_04969_),
    .Y(_04970_));
 sky130_fd_sc_hd__a221o_2 _26350_ (.A1(_17038_),
    .A2(\reg_next_pc[23] ),
    .B1(_01530_),
    .B2(_04898_),
    .C1(_04970_),
    .X(_02116_));
 sky130_vsdinv _26351_ (.A(_17489_),
    .Y(_04971_));
 sky130_fd_sc_hd__nand3_2 _26352_ (.A(_04965_),
    .B(_17492_),
    .C(_04240_),
    .Y(_04972_));
 sky130_fd_sc_hd__xor2_2 _26353_ (.A(_04971_),
    .B(_04972_),
    .X(_02117_));
 sky130_fd_sc_hd__buf_1 _26354_ (.A(_04924_),
    .X(_04973_));
 sky130_fd_sc_hd__and2_2 _26355_ (.A(_04966_),
    .B(\reg_next_pc[24] ),
    .X(_04974_));
 sky130_fd_sc_hd__a221o_2 _26356_ (.A1(_16915_),
    .A2(_04973_),
    .B1(_04959_),
    .B2(_01533_),
    .C1(_04974_),
    .X(_02118_));
 sky130_fd_sc_hd__nor2_2 _26357_ (.A(_04971_),
    .B(_04972_),
    .Y(_04975_));
 sky130_fd_sc_hd__xor2_2 _26358_ (.A(_17484_),
    .B(_04975_),
    .X(_02119_));
 sky130_fd_sc_hd__buf_1 _26359_ (.A(_04928_),
    .X(_04976_));
 sky130_fd_sc_hd__and2_2 _26360_ (.A(_04966_),
    .B(\reg_next_pc[25] ),
    .X(_04977_));
 sky130_fd_sc_hd__a221o_2 _26361_ (.A1(_16917_),
    .A2(_04973_),
    .B1(_04976_),
    .B2(_01536_),
    .C1(_04977_),
    .X(_02120_));
 sky130_fd_sc_hd__nor3b_2 _26362_ (.A(_04971_),
    .B(_04972_),
    .C_N(_17484_),
    .Y(_04978_));
 sky130_fd_sc_hd__xor2_2 _26363_ (.A(_17480_),
    .B(_04978_),
    .X(_02121_));
 sky130_fd_sc_hd__and2_2 _26364_ (.A(_04966_),
    .B(\reg_next_pc[26] ),
    .X(_04979_));
 sky130_fd_sc_hd__a221o_2 _26365_ (.A1(_16916_),
    .A2(_04973_),
    .B1(_04976_),
    .B2(_01539_),
    .C1(_04979_),
    .X(_02122_));
 sky130_fd_sc_hd__nand3_2 _26366_ (.A(_04975_),
    .B(\reg_pc[26] ),
    .C(_17483_),
    .Y(_04980_));
 sky130_fd_sc_hd__xnor2_2 _26367_ (.A(_17476_),
    .B(_04980_),
    .Y(_02123_));
 sky130_fd_sc_hd__a32o_2 _26368_ (.A1(_16914_),
    .A2(_17035_),
    .A3(_17881_),
    .B1(_19772_),
    .B2(\reg_next_pc[27] ),
    .X(_04981_));
 sky130_fd_sc_hd__a21o_2 _26369_ (.A1(_01542_),
    .A2(_04899_),
    .B1(_04981_),
    .X(_02124_));
 sky130_fd_sc_hd__and4_2 _26370_ (.A(_04975_),
    .B(\reg_pc[27] ),
    .C(_17480_),
    .D(_17483_),
    .X(_04982_));
 sky130_fd_sc_hd__xor2_2 _26371_ (.A(_17471_),
    .B(_04982_),
    .X(_02125_));
 sky130_fd_sc_hd__buf_1 _26372_ (.A(_17036_),
    .X(_04983_));
 sky130_fd_sc_hd__and2_2 _26373_ (.A(_04983_),
    .B(\reg_next_pc[28] ),
    .X(_04984_));
 sky130_fd_sc_hd__a221o_2 _26374_ (.A1(_16908_),
    .A2(_04973_),
    .B1(_04976_),
    .B2(_01545_),
    .C1(_04984_),
    .X(_02126_));
 sky130_vsdinv _26375_ (.A(\reg_pc[28] ),
    .Y(_04985_));
 sky130_fd_sc_hd__nor3b_2 _26376_ (.A(_04985_),
    .B(_04980_),
    .C_N(_17476_),
    .Y(_04986_));
 sky130_fd_sc_hd__xor2_2 _26377_ (.A(_17467_),
    .B(_04986_),
    .X(_02127_));
 sky130_fd_sc_hd__and2_2 _26378_ (.A(_04983_),
    .B(\reg_next_pc[29] ),
    .X(_04987_));
 sky130_fd_sc_hd__a221o_2 _26379_ (.A1(_16911_),
    .A2(_17046_),
    .B1(_04976_),
    .B2(_01548_),
    .C1(_04987_),
    .X(_02128_));
 sky130_fd_sc_hd__nand3_2 _26380_ (.A(_04982_),
    .B(\reg_pc[29] ),
    .C(_17471_),
    .Y(_04988_));
 sky130_fd_sc_hd__xnor2_2 _26381_ (.A(_17465_),
    .B(_04988_),
    .Y(_02129_));
 sky130_fd_sc_hd__and2_2 _26382_ (.A(_04983_),
    .B(\reg_next_pc[30] ),
    .X(_04989_));
 sky130_fd_sc_hd__a221o_2 _26383_ (.A1(_16909_),
    .A2(_17046_),
    .B1(_04903_),
    .B2(_01551_),
    .C1(_04989_),
    .X(_02130_));
 sky130_fd_sc_hd__nand3_2 _26384_ (.A(_04986_),
    .B(_17465_),
    .C(_17467_),
    .Y(_04990_));
 sky130_fd_sc_hd__xnor2_2 _26385_ (.A(\reg_pc[31] ),
    .B(_04990_),
    .Y(_02131_));
 sky130_fd_sc_hd__and2_2 _26386_ (.A(_04983_),
    .B(\reg_next_pc[31] ),
    .X(_04991_));
 sky130_fd_sc_hd__a221o_2 _26387_ (.A1(_16910_),
    .A2(_17046_),
    .B1(_04903_),
    .B2(_01554_),
    .C1(_04991_),
    .X(_02132_));
 sky130_fd_sc_hd__nor2_2 _26388_ (.A(instr_or),
    .B(instr_ori),
    .Y(_04992_));
 sky130_vsdinv _26389_ (.A(_04992_),
    .Y(_04993_));
 sky130_fd_sc_hd__buf_1 _26390_ (.A(_04993_),
    .X(_04994_));
 sky130_fd_sc_hd__buf_1 _26391_ (.A(_04994_),
    .X(_04995_));
 sky130_fd_sc_hd__nor3b_2 _26392_ (.A(is_compare),
    .B(_04995_),
    .C_N(_16993_),
    .Y(_04996_));
 sky130_fd_sc_hd__nor2_2 _26393_ (.A(_17303_),
    .B(_17347_),
    .Y(_04997_));
 sky130_fd_sc_hd__buf_1 _26394_ (.A(_04997_),
    .X(_04998_));
 sky130_fd_sc_hd__buf_1 _26395_ (.A(_04998_),
    .X(_04999_));
 sky130_fd_sc_hd__buf_1 _26396_ (.A(instr_and),
    .X(_05000_));
 sky130_fd_sc_hd__buf_1 _26397_ (.A(instr_andi),
    .X(_05001_));
 sky130_fd_sc_hd__nor2_2 _26398_ (.A(_05000_),
    .B(_05001_),
    .Y(_05002_));
 sky130_fd_sc_hd__buf_1 _26399_ (.A(_05002_),
    .X(_05003_));
 sky130_fd_sc_hd__nor2_2 _26400_ (.A(instr_sll),
    .B(instr_slli),
    .Y(_05004_));
 sky130_fd_sc_hd__and4_2 _26401_ (.A(_04996_),
    .B(_04999_),
    .C(_05003_),
    .D(_05004_),
    .X(_02133_));
 sky130_fd_sc_hd__buf_1 _26402_ (.A(_16994_),
    .X(_05005_));
 sky130_fd_sc_hd__buf_1 _26403_ (.A(_05005_),
    .X(_05006_));
 sky130_vsdinv _26404_ (.A(_04997_),
    .Y(_05007_));
 sky130_fd_sc_hd__buf_1 _26405_ (.A(_05007_),
    .X(_05008_));
 sky130_vsdinv _26406_ (.A(_05004_),
    .Y(_05009_));
 sky130_fd_sc_hd__buf_1 _26407_ (.A(_05009_),
    .X(_05010_));
 sky130_fd_sc_hd__buf_1 _26408_ (.A(_05010_),
    .X(_05011_));
 sky130_fd_sc_hd__o211a_2 _26409_ (.A1(_05000_),
    .A2(_05001_),
    .B1(_18453_),
    .C1(_19122_),
    .X(_05012_));
 sky130_fd_sc_hd__nor2_2 _26410_ (.A(_18453_),
    .B(_19122_),
    .Y(_05013_));
 sky130_fd_sc_hd__o2bb2ai_2 _26411_ (.A1_N(_17072_),
    .A2_N(is_compare),
    .B1(_04992_),
    .B2(_05013_),
    .Y(_05014_));
 sky130_fd_sc_hd__a211o_2 _26412_ (.A1(\alu_shl[0] ),
    .A2(_05011_),
    .B1(_05012_),
    .C1(_05014_),
    .X(_05015_));
 sky130_fd_sc_hd__a221o_2 _26413_ (.A1(\alu_shr[0] ),
    .A2(_05006_),
    .B1(_02591_),
    .B2(_05008_),
    .C1(_05015_),
    .X(_02134_));
 sky130_fd_sc_hd__buf_1 _26414_ (.A(_05007_),
    .X(_05016_));
 sky130_fd_sc_hd__buf_1 _26415_ (.A(_05016_),
    .X(_05017_));
 sky130_fd_sc_hd__buf_1 _26416_ (.A(_05005_),
    .X(_05018_));
 sky130_fd_sc_hd__buf_1 _26417_ (.A(_17275_),
    .X(_05019_));
 sky130_fd_sc_hd__buf_1 _26418_ (.A(_17339_),
    .X(_05020_));
 sky130_fd_sc_hd__o22a_2 _26419_ (.A1(_05019_),
    .A2(_05020_),
    .B1(_18449_),
    .B2(_04446_),
    .X(_05021_));
 sky130_fd_sc_hd__buf_1 _26420_ (.A(_17269_),
    .X(_05022_));
 sky130_fd_sc_hd__buf_1 _26421_ (.A(_17334_),
    .X(_05023_));
 sky130_fd_sc_hd__o211a_2 _26422_ (.A1(_05022_),
    .A2(_05023_),
    .B1(_18450_),
    .C1(_04446_),
    .X(_05024_));
 sky130_fd_sc_hd__a211o_2 _26423_ (.A1(\alu_shl[1] ),
    .A2(_05011_),
    .B1(_05021_),
    .C1(_05024_),
    .X(_05025_));
 sky130_fd_sc_hd__a221o_2 _26424_ (.A1(_19741_),
    .A2(_05017_),
    .B1(_05018_),
    .B2(\alu_shr[1] ),
    .C1(_05025_),
    .X(_02135_));
 sky130_fd_sc_hd__buf_1 _26425_ (.A(_16994_),
    .X(_05026_));
 sky130_fd_sc_hd__buf_1 _26426_ (.A(_05026_),
    .X(_05027_));
 sky130_fd_sc_hd__o211a_2 _26427_ (.A1(_17303_),
    .A2(_17347_),
    .B1(_19730_),
    .C1(_19729_),
    .X(_05028_));
 sky130_fd_sc_hd__buf_1 _26428_ (.A(_05009_),
    .X(_05029_));
 sky130_fd_sc_hd__buf_1 _26429_ (.A(_05002_),
    .X(_05030_));
 sky130_fd_sc_hd__nor2_2 _26430_ (.A(_19730_),
    .B(_05030_),
    .Y(_05031_));
 sky130_fd_sc_hd__a221o_2 _26431_ (.A1(_05029_),
    .A2(\alu_shl[2] ),
    .B1(_04995_),
    .B2(_19729_),
    .C1(_05031_),
    .X(_05032_));
 sky130_fd_sc_hd__a211o_2 _26432_ (.A1(\alu_shr[2] ),
    .A2(_05027_),
    .B1(_05028_),
    .C1(_05032_),
    .X(_02136_));
 sky130_fd_sc_hd__nor2_2 _26433_ (.A(_04999_),
    .B(_19727_),
    .Y(_05033_));
 sky130_fd_sc_hd__or2_2 _26434_ (.A(_18444_),
    .B(_19110_),
    .X(_05034_));
 sky130_fd_sc_hd__o211a_2 _26435_ (.A1(_17270_),
    .A2(_17335_),
    .B1(_18444_),
    .C1(_19110_),
    .X(_05035_));
 sky130_fd_sc_hd__a221o_2 _26436_ (.A1(_05029_),
    .A2(\alu_shl[3] ),
    .B1(_04995_),
    .B2(_05034_),
    .C1(_05035_),
    .X(_05036_));
 sky130_fd_sc_hd__a211o_2 _26437_ (.A1(\alu_shr[3] ),
    .A2(_05027_),
    .B1(_05033_),
    .C1(_05036_),
    .X(_02137_));
 sky130_fd_sc_hd__nor3_2 _26438_ (.A(_19733_),
    .B(_04999_),
    .C(_19734_),
    .Y(_05037_));
 sky130_fd_sc_hd__buf_1 _26439_ (.A(_05010_),
    .X(_05038_));
 sky130_vsdinv _26440_ (.A(_19733_),
    .Y(_05039_));
 sky130_fd_sc_hd__buf_1 _26441_ (.A(_04993_),
    .X(_05040_));
 sky130_fd_sc_hd__o211a_2 _26442_ (.A1(_17270_),
    .A2(_17335_),
    .B1(_18441_),
    .C1(_19107_),
    .X(_05041_));
 sky130_fd_sc_hd__a221o_2 _26443_ (.A1(_05038_),
    .A2(\alu_shl[4] ),
    .B1(_05039_),
    .B2(_05040_),
    .C1(_05041_),
    .X(_05042_));
 sky130_fd_sc_hd__a211o_2 _26444_ (.A1(\alu_shr[4] ),
    .A2(_05027_),
    .B1(_05037_),
    .C1(_05042_),
    .X(_02138_));
 sky130_fd_sc_hd__buf_1 _26445_ (.A(_04998_),
    .X(_05043_));
 sky130_fd_sc_hd__nor3_2 _26446_ (.A(_19735_),
    .B(_05043_),
    .C(_19736_),
    .Y(_05044_));
 sky130_vsdinv _26447_ (.A(_19735_),
    .Y(_05045_));
 sky130_fd_sc_hd__buf_1 _26448_ (.A(_05000_),
    .X(_05046_));
 sky130_fd_sc_hd__buf_1 _26449_ (.A(_05001_),
    .X(_05047_));
 sky130_fd_sc_hd__o211a_2 _26450_ (.A1(_05046_),
    .A2(_05047_),
    .B1(_18439_),
    .C1(_19105_),
    .X(_05048_));
 sky130_fd_sc_hd__a221o_2 _26451_ (.A1(_05038_),
    .A2(\alu_shl[5] ),
    .B1(_05045_),
    .B2(_05040_),
    .C1(_05048_),
    .X(_05049_));
 sky130_fd_sc_hd__a211o_2 _26452_ (.A1(\alu_shr[5] ),
    .A2(_05027_),
    .B1(_05044_),
    .C1(_05049_),
    .X(_02139_));
 sky130_fd_sc_hd__xor2_2 _26453_ (.A(_18435_),
    .B(_19102_),
    .X(_05050_));
 sky130_fd_sc_hd__buf_1 _26454_ (.A(_05009_),
    .X(_05051_));
 sky130_fd_sc_hd__buf_1 _26455_ (.A(_04993_),
    .X(_05052_));
 sky130_fd_sc_hd__nor2_2 _26456_ (.A(_19740_),
    .B(_05030_),
    .Y(_05053_));
 sky130_fd_sc_hd__a221o_2 _26457_ (.A1(_05051_),
    .A2(\alu_shl[6] ),
    .B1(_05052_),
    .B2(_19739_),
    .C1(_05053_),
    .X(_05054_));
 sky130_fd_sc_hd__a221o_2 _26458_ (.A1(\alu_shr[6] ),
    .A2(_05006_),
    .B1(_05050_),
    .B2(_05008_),
    .C1(_05054_),
    .X(_02140_));
 sky130_fd_sc_hd__buf_1 _26459_ (.A(_05026_),
    .X(_05055_));
 sky130_fd_sc_hd__o22a_2 _26460_ (.A1(_05019_),
    .A2(_05020_),
    .B1(_18432_),
    .B2(_19099_),
    .X(_05056_));
 sky130_fd_sc_hd__buf_1 _26461_ (.A(_17269_),
    .X(_05057_));
 sky130_fd_sc_hd__buf_1 _26462_ (.A(_17334_),
    .X(_05058_));
 sky130_fd_sc_hd__o211a_2 _26463_ (.A1(_05057_),
    .A2(_05058_),
    .B1(_18433_),
    .C1(_19099_),
    .X(_05059_));
 sky130_fd_sc_hd__a211o_2 _26464_ (.A1(\alu_shl[7] ),
    .A2(_05011_),
    .B1(_05056_),
    .C1(_05059_),
    .X(_05060_));
 sky130_fd_sc_hd__a221o_2 _26465_ (.A1(_19742_),
    .A2(_05017_),
    .B1(_05055_),
    .B2(\alu_shr[7] ),
    .C1(_05060_),
    .X(_02141_));
 sky130_fd_sc_hd__buf_1 _26466_ (.A(_05026_),
    .X(_05061_));
 sky130_fd_sc_hd__nor3_2 _26467_ (.A(_19745_),
    .B(_05043_),
    .C(_19746_),
    .Y(_05062_));
 sky130_vsdinv _26468_ (.A(_19745_),
    .Y(_05063_));
 sky130_fd_sc_hd__o211a_2 _26469_ (.A1(_05046_),
    .A2(_05047_),
    .B1(_18430_),
    .C1(_19096_),
    .X(_05064_));
 sky130_fd_sc_hd__a221o_2 _26470_ (.A1(_05038_),
    .A2(\alu_shl[8] ),
    .B1(_05063_),
    .B2(_05040_),
    .C1(_05064_),
    .X(_05065_));
 sky130_fd_sc_hd__a211o_2 _26471_ (.A1(\alu_shr[8] ),
    .A2(_05061_),
    .B1(_05062_),
    .C1(_05065_),
    .X(_02142_));
 sky130_fd_sc_hd__nor2_2 _26472_ (.A(_04999_),
    .B(_19747_),
    .Y(_05066_));
 sky130_fd_sc_hd__or2_2 _26473_ (.A(_18427_),
    .B(_19093_),
    .X(_05067_));
 sky130_fd_sc_hd__o211a_2 _26474_ (.A1(_05046_),
    .A2(_05047_),
    .B1(_18427_),
    .C1(_19093_),
    .X(_05068_));
 sky130_fd_sc_hd__a221o_2 _26475_ (.A1(_05038_),
    .A2(\alu_shl[9] ),
    .B1(_04995_),
    .B2(_05067_),
    .C1(_05068_),
    .X(_05069_));
 sky130_fd_sc_hd__a211o_2 _26476_ (.A1(\alu_shr[9] ),
    .A2(_05061_),
    .B1(_05066_),
    .C1(_05069_),
    .X(_02143_));
 sky130_fd_sc_hd__or2_2 _26477_ (.A(_18425_),
    .B(_19090_),
    .X(_05070_));
 sky130_fd_sc_hd__nand2_2 _26478_ (.A(_18425_),
    .B(_19090_),
    .Y(_05071_));
 sky130_fd_sc_hd__nor2_2 _26479_ (.A(_05071_),
    .B(_05030_),
    .Y(_05072_));
 sky130_fd_sc_hd__a221o_2 _26480_ (.A1(_05051_),
    .A2(\alu_shl[10] ),
    .B1(_05052_),
    .B2(_05070_),
    .C1(_05072_),
    .X(_05073_));
 sky130_fd_sc_hd__a221o_2 _26481_ (.A1(_19752_),
    .A2(_05017_),
    .B1(_05055_),
    .B2(\alu_shr[10] ),
    .C1(_05073_),
    .X(_02144_));
 sky130_vsdinv _26482_ (.A(_19748_),
    .Y(_05074_));
 sky130_fd_sc_hd__o211a_2 _26483_ (.A1(_05000_),
    .A2(_05001_),
    .B1(_18423_),
    .C1(_19087_),
    .X(_05075_));
 sky130_fd_sc_hd__a221o_2 _26484_ (.A1(_05051_),
    .A2(\alu_shl[11] ),
    .B1(_05074_),
    .B2(_04994_),
    .C1(_05075_),
    .X(_05076_));
 sky130_fd_sc_hd__a221o_2 _26485_ (.A1(_19750_),
    .A2(_05017_),
    .B1(_05055_),
    .B2(\alu_shr[11] ),
    .C1(_05076_),
    .X(_02145_));
 sky130_fd_sc_hd__buf_1 _26486_ (.A(_05016_),
    .X(_05077_));
 sky130_fd_sc_hd__o22a_2 _26487_ (.A1(_05019_),
    .A2(_05020_),
    .B1(pcpi_rs2[12]),
    .B2(_19085_),
    .X(_05078_));
 sky130_fd_sc_hd__o211a_2 _26488_ (.A1(_05057_),
    .A2(_05058_),
    .B1(_18421_),
    .C1(_19085_),
    .X(_05079_));
 sky130_fd_sc_hd__a211o_2 _26489_ (.A1(\alu_shl[12] ),
    .A2(_05011_),
    .B1(_05078_),
    .C1(_05079_),
    .X(_05080_));
 sky130_fd_sc_hd__a221o_2 _26490_ (.A1(_19723_),
    .A2(_05077_),
    .B1(_05055_),
    .B2(\alu_shr[12] ),
    .C1(_05080_),
    .X(_02146_));
 sky130_fd_sc_hd__buf_1 _26491_ (.A(_05026_),
    .X(_05081_));
 sky130_fd_sc_hd__inv_2 _26492_ (.A(_18419_),
    .Y(_02354_));
 sky130_vsdinv _26493_ (.A(_19083_),
    .Y(_05082_));
 sky130_fd_sc_hd__o21ai_2 _26494_ (.A1(_17316_),
    .A2(_19009_),
    .B1(\alu_shl[13] ),
    .Y(_05083_));
 sky130_fd_sc_hd__o22ai_2 _26495_ (.A1(_17276_),
    .A2(_17340_),
    .B1(_18420_),
    .B2(_19083_),
    .Y(_05084_));
 sky130_fd_sc_hd__o311ai_2 _26496_ (.A1(_02354_),
    .A2(_05082_),
    .A3(_05003_),
    .B1(_05083_),
    .C1(_05084_),
    .Y(_05085_));
 sky130_fd_sc_hd__a221o_2 _26497_ (.A1(_19724_),
    .A2(_05077_),
    .B1(_05081_),
    .B2(\alu_shr[13] ),
    .C1(_05085_),
    .X(_02147_));
 sky130_fd_sc_hd__nor2_2 _26498_ (.A(_18417_),
    .B(_19081_),
    .Y(_05086_));
 sky130_fd_sc_hd__o21ai_2 _26499_ (.A1(_17316_),
    .A2(_19009_),
    .B1(\alu_shl[14] ),
    .Y(_05087_));
 sky130_fd_sc_hd__o211ai_2 _26500_ (.A1(_17270_),
    .A2(_17335_),
    .B1(_18417_),
    .C1(_19081_),
    .Y(_05088_));
 sky130_fd_sc_hd__o211ai_2 _26501_ (.A1(_05086_),
    .A2(_04992_),
    .B1(_05087_),
    .C1(_05088_),
    .Y(_05089_));
 sky130_fd_sc_hd__a221o_2 _26502_ (.A1(_19725_),
    .A2(_05077_),
    .B1(_05081_),
    .B2(\alu_shr[14] ),
    .C1(_05089_),
    .X(_02148_));
 sky130_fd_sc_hd__buf_1 _26503_ (.A(_05010_),
    .X(_05090_));
 sky130_fd_sc_hd__o22a_2 _26504_ (.A1(_05019_),
    .A2(_05020_),
    .B1(_18415_),
    .B2(_19077_),
    .X(_05091_));
 sky130_fd_sc_hd__o211a_2 _26505_ (.A1(_05057_),
    .A2(_05058_),
    .B1(_18415_),
    .C1(_19077_),
    .X(_05092_));
 sky130_fd_sc_hd__a211o_2 _26506_ (.A1(\alu_shl[15] ),
    .A2(_05090_),
    .B1(_05091_),
    .C1(_05092_),
    .X(_05093_));
 sky130_fd_sc_hd__a221o_2 _26507_ (.A1(_19722_),
    .A2(_05077_),
    .B1(_05081_),
    .B2(\alu_shr[15] ),
    .C1(_05093_),
    .X(_02149_));
 sky130_fd_sc_hd__buf_1 _26508_ (.A(_05016_),
    .X(_05094_));
 sky130_fd_sc_hd__buf_1 _26509_ (.A(_17275_),
    .X(_05095_));
 sky130_fd_sc_hd__buf_1 _26510_ (.A(_17339_),
    .X(_05096_));
 sky130_fd_sc_hd__o22a_2 _26511_ (.A1(_05095_),
    .A2(_05096_),
    .B1(_18412_),
    .B2(_19074_),
    .X(_05097_));
 sky130_fd_sc_hd__o211a_2 _26512_ (.A1(_05057_),
    .A2(_05058_),
    .B1(_18412_),
    .C1(_19074_),
    .X(_05098_));
 sky130_fd_sc_hd__a211o_2 _26513_ (.A1(\alu_shl[16] ),
    .A2(_05090_),
    .B1(_05097_),
    .C1(_05098_),
    .X(_05099_));
 sky130_fd_sc_hd__a221o_2 _26514_ (.A1(_19696_),
    .A2(_05094_),
    .B1(_05081_),
    .B2(\alu_shr[16] ),
    .C1(_05099_),
    .X(_02150_));
 sky130_fd_sc_hd__buf_1 _26515_ (.A(_05005_),
    .X(_05100_));
 sky130_fd_sc_hd__inv_2 _26516_ (.A(_18410_),
    .Y(_02366_));
 sky130_vsdinv _26517_ (.A(_19072_),
    .Y(_05101_));
 sky130_fd_sc_hd__o21ai_2 _26518_ (.A1(_17316_),
    .A2(_19009_),
    .B1(\alu_shl[17] ),
    .Y(_05102_));
 sky130_fd_sc_hd__o22ai_2 _26519_ (.A1(_17276_),
    .A2(_17340_),
    .B1(_18411_),
    .B2(_19072_),
    .Y(_05103_));
 sky130_fd_sc_hd__o311ai_2 _26520_ (.A1(_02366_),
    .A2(_05101_),
    .A3(_05003_),
    .B1(_05102_),
    .C1(_05103_),
    .Y(_05104_));
 sky130_fd_sc_hd__a221o_2 _26521_ (.A1(_19697_),
    .A2(_05094_),
    .B1(_05100_),
    .B2(\alu_shr[17] ),
    .C1(_05104_),
    .X(_02151_));
 sky130_fd_sc_hd__buf_1 _26522_ (.A(_05009_),
    .X(_05105_));
 sky130_fd_sc_hd__or2_2 _26523_ (.A(_18408_),
    .B(_19069_),
    .X(_05106_));
 sky130_fd_sc_hd__nand2_2 _26524_ (.A(_18408_),
    .B(_19069_),
    .Y(_05107_));
 sky130_fd_sc_hd__buf_1 _26525_ (.A(_05002_),
    .X(_05108_));
 sky130_fd_sc_hd__nor2_2 _26526_ (.A(_05107_),
    .B(_05108_),
    .Y(_05109_));
 sky130_fd_sc_hd__a221o_2 _26527_ (.A1(_05105_),
    .A2(\alu_shl[18] ),
    .B1(_05052_),
    .B2(_05106_),
    .C1(_05109_),
    .X(_05110_));
 sky130_fd_sc_hd__a221o_2 _26528_ (.A1(_19698_),
    .A2(_05094_),
    .B1(_05100_),
    .B2(\alu_shr[18] ),
    .C1(_05110_),
    .X(_02152_));
 sky130_fd_sc_hd__o22a_2 _26529_ (.A1(_05095_),
    .A2(_05096_),
    .B1(_18406_),
    .B2(_19066_),
    .X(_05111_));
 sky130_fd_sc_hd__buf_1 _26530_ (.A(_17269_),
    .X(_05112_));
 sky130_fd_sc_hd__buf_1 _26531_ (.A(_17334_),
    .X(_05113_));
 sky130_fd_sc_hd__o211a_2 _26532_ (.A1(_05112_),
    .A2(_05113_),
    .B1(_18407_),
    .C1(_19066_),
    .X(_05114_));
 sky130_fd_sc_hd__a211o_2 _26533_ (.A1(\alu_shl[19] ),
    .A2(_05090_),
    .B1(_05111_),
    .C1(_05114_),
    .X(_05115_));
 sky130_fd_sc_hd__a221o_2 _26534_ (.A1(_19695_),
    .A2(_05094_),
    .B1(_05100_),
    .B2(\alu_shr[19] ),
    .C1(_05115_),
    .X(_02153_));
 sky130_fd_sc_hd__buf_1 _26535_ (.A(_05007_),
    .X(_05116_));
 sky130_fd_sc_hd__o22a_2 _26536_ (.A1(_05095_),
    .A2(_05096_),
    .B1(_18404_),
    .B2(_19064_),
    .X(_05117_));
 sky130_fd_sc_hd__o211a_2 _26537_ (.A1(_05112_),
    .A2(_05113_),
    .B1(_18404_),
    .C1(_19064_),
    .X(_05118_));
 sky130_fd_sc_hd__a211o_2 _26538_ (.A1(\alu_shl[20] ),
    .A2(_05090_),
    .B1(_05117_),
    .C1(_05118_),
    .X(_05119_));
 sky130_fd_sc_hd__a221o_2 _26539_ (.A1(_19691_),
    .A2(_05116_),
    .B1(_05100_),
    .B2(\alu_shr[20] ),
    .C1(_05119_),
    .X(_02154_));
 sky130_fd_sc_hd__buf_1 _26540_ (.A(_05005_),
    .X(_05120_));
 sky130_fd_sc_hd__inv_2 _26541_ (.A(_18402_),
    .Y(_02378_));
 sky130_vsdinv _26542_ (.A(_19062_),
    .Y(_05121_));
 sky130_fd_sc_hd__o21ai_2 _26543_ (.A1(instr_sll),
    .A2(instr_slli),
    .B1(\alu_shl[21] ),
    .Y(_05122_));
 sky130_fd_sc_hd__o22ai_2 _26544_ (.A1(_17276_),
    .A2(_17340_),
    .B1(_18403_),
    .B2(_19062_),
    .Y(_05123_));
 sky130_fd_sc_hd__o311ai_2 _26545_ (.A1(_02378_),
    .A2(_05121_),
    .A3(_05003_),
    .B1(_05122_),
    .C1(_05123_),
    .Y(_05124_));
 sky130_fd_sc_hd__a221o_2 _26546_ (.A1(_19692_),
    .A2(_05116_),
    .B1(_05120_),
    .B2(\alu_shr[21] ),
    .C1(_05124_),
    .X(_02155_));
 sky130_fd_sc_hd__or2_2 _26547_ (.A(_18400_),
    .B(_19060_),
    .X(_05125_));
 sky130_fd_sc_hd__nand2_2 _26548_ (.A(_18400_),
    .B(_19060_),
    .Y(_05126_));
 sky130_fd_sc_hd__nor2_2 _26549_ (.A(_05126_),
    .B(_05108_),
    .Y(_05127_));
 sky130_fd_sc_hd__a221o_2 _26550_ (.A1(_05105_),
    .A2(\alu_shl[22] ),
    .B1(_05052_),
    .B2(_05125_),
    .C1(_05127_),
    .X(_05128_));
 sky130_fd_sc_hd__a221o_2 _26551_ (.A1(_19693_),
    .A2(_05116_),
    .B1(_05120_),
    .B2(\alu_shr[22] ),
    .C1(_05128_),
    .X(_02156_));
 sky130_fd_sc_hd__o22a_2 _26552_ (.A1(_05095_),
    .A2(_05096_),
    .B1(_18398_),
    .B2(_19057_),
    .X(_05129_));
 sky130_fd_sc_hd__o211a_2 _26553_ (.A1(_05112_),
    .A2(_05113_),
    .B1(_18399_),
    .C1(_19057_),
    .X(_05130_));
 sky130_fd_sc_hd__a211o_2 _26554_ (.A1(\alu_shl[23] ),
    .A2(_05029_),
    .B1(_05129_),
    .C1(_05130_),
    .X(_05131_));
 sky130_fd_sc_hd__a221o_2 _26555_ (.A1(_19690_),
    .A2(_05116_),
    .B1(_05120_),
    .B2(\alu_shr[23] ),
    .C1(_05131_),
    .X(_02157_));
 sky130_fd_sc_hd__nor3_2 _26556_ (.A(_19704_),
    .B(_05043_),
    .C(_19705_),
    .Y(_05132_));
 sky130_fd_sc_hd__buf_1 _26557_ (.A(_05010_),
    .X(_05133_));
 sky130_vsdinv _26558_ (.A(_19704_),
    .Y(_05134_));
 sky130_fd_sc_hd__buf_1 _26559_ (.A(_04993_),
    .X(_05135_));
 sky130_fd_sc_hd__o211a_2 _26560_ (.A1(_05046_),
    .A2(_05047_),
    .B1(_18396_),
    .C1(_19054_),
    .X(_05136_));
 sky130_fd_sc_hd__a221o_2 _26561_ (.A1(_05133_),
    .A2(\alu_shl[24] ),
    .B1(_05134_),
    .B2(_05135_),
    .C1(_05136_),
    .X(_05137_));
 sky130_fd_sc_hd__a211o_2 _26562_ (.A1(\alu_shr[24] ),
    .A2(_05061_),
    .B1(_05132_),
    .C1(_05137_),
    .X(_02158_));
 sky130_fd_sc_hd__nor3_2 _26563_ (.A(_19706_),
    .B(_05043_),
    .C(_19707_),
    .Y(_05138_));
 sky130_vsdinv _26564_ (.A(_19706_),
    .Y(_05139_));
 sky130_fd_sc_hd__o211a_2 _26565_ (.A1(_05022_),
    .A2(_05023_),
    .B1(_18394_),
    .C1(_19053_),
    .X(_05140_));
 sky130_fd_sc_hd__a221o_2 _26566_ (.A1(_05133_),
    .A2(\alu_shl[25] ),
    .B1(_05139_),
    .B2(_05135_),
    .C1(_05140_),
    .X(_05141_));
 sky130_fd_sc_hd__a211o_2 _26567_ (.A1(\alu_shr[25] ),
    .A2(_05061_),
    .B1(_05138_),
    .C1(_05141_),
    .X(_02159_));
 sky130_fd_sc_hd__o22a_2 _26568_ (.A1(_17275_),
    .A2(_17339_),
    .B1(_18392_),
    .B2(_19050_),
    .X(_05142_));
 sky130_fd_sc_hd__o211a_2 _26569_ (.A1(_05112_),
    .A2(_05113_),
    .B1(_18392_),
    .C1(_19050_),
    .X(_05143_));
 sky130_fd_sc_hd__a211o_2 _26570_ (.A1(\alu_shl[26] ),
    .A2(_05029_),
    .B1(_05142_),
    .C1(_05143_),
    .X(_05144_));
 sky130_fd_sc_hd__a221o_2 _26571_ (.A1(_19702_),
    .A2(_05008_),
    .B1(_05120_),
    .B2(\alu_shr[26] ),
    .C1(_05144_),
    .X(_02160_));
 sky130_fd_sc_hd__or2_2 _26572_ (.A(pcpi_rs2[27]),
    .B(_19048_),
    .X(_05145_));
 sky130_fd_sc_hd__nand2_2 _26573_ (.A(_18391_),
    .B(_19048_),
    .Y(_05146_));
 sky130_fd_sc_hd__nor2_2 _26574_ (.A(_05146_),
    .B(_05108_),
    .Y(_05147_));
 sky130_fd_sc_hd__a221o_2 _26575_ (.A1(_05105_),
    .A2(\alu_shl[27] ),
    .B1(_04994_),
    .B2(_05145_),
    .C1(_05147_),
    .X(_05148_));
 sky130_fd_sc_hd__a221o_2 _26576_ (.A1(_19700_),
    .A2(_05008_),
    .B1(_05006_),
    .B2(\alu_shr[27] ),
    .C1(_05148_),
    .X(_02161_));
 sky130_fd_sc_hd__o211a_2 _26577_ (.A1(_17303_),
    .A2(_17347_),
    .B1(_19717_),
    .C1(_19716_),
    .X(_05149_));
 sky130_fd_sc_hd__nor2_2 _26578_ (.A(_19717_),
    .B(_05030_),
    .Y(_05150_));
 sky130_fd_sc_hd__a221o_2 _26579_ (.A1(_05133_),
    .A2(\alu_shl[28] ),
    .B1(_05040_),
    .B2(_19716_),
    .C1(_05150_),
    .X(_05151_));
 sky130_fd_sc_hd__a211o_2 _26580_ (.A1(\alu_shr[28] ),
    .A2(_05018_),
    .B1(_05149_),
    .C1(_05151_),
    .X(_02162_));
 sky130_fd_sc_hd__nor3_2 _26581_ (.A(_19714_),
    .B(_04998_),
    .C(_19713_),
    .Y(_05152_));
 sky130_vsdinv _26582_ (.A(_19714_),
    .Y(_05153_));
 sky130_fd_sc_hd__o211a_2 _26583_ (.A1(_05022_),
    .A2(_05023_),
    .B1(_18386_),
    .C1(_19044_),
    .X(_05154_));
 sky130_fd_sc_hd__a221o_2 _26584_ (.A1(_05133_),
    .A2(\alu_shl[29] ),
    .B1(_05153_),
    .B2(_05135_),
    .C1(_05154_),
    .X(_05155_));
 sky130_fd_sc_hd__a211o_2 _26585_ (.A1(\alu_shr[29] ),
    .A2(_05018_),
    .B1(_05152_),
    .C1(_05155_),
    .X(_02163_));
 sky130_fd_sc_hd__nor3_2 _26586_ (.A(_19709_),
    .B(_04998_),
    .C(_19710_),
    .Y(_05156_));
 sky130_vsdinv _26587_ (.A(_19709_),
    .Y(_05157_));
 sky130_fd_sc_hd__o211a_2 _26588_ (.A1(_05022_),
    .A2(_05023_),
    .B1(_18385_),
    .C1(_04276_),
    .X(_05158_));
 sky130_fd_sc_hd__a221o_2 _26589_ (.A1(_05051_),
    .A2(\alu_shl[30] ),
    .B1(_05157_),
    .B2(_05135_),
    .C1(_05158_),
    .X(_05159_));
 sky130_fd_sc_hd__a211o_2 _26590_ (.A1(\alu_shr[30] ),
    .A2(_05018_),
    .B1(_05156_),
    .C1(_05159_),
    .X(_02164_));
 sky130_fd_sc_hd__or2_2 _26591_ (.A(pcpi_rs1[31]),
    .B(_16977_),
    .X(_05160_));
 sky130_fd_sc_hd__nand2_2 _26592_ (.A(_16957_),
    .B(_16977_),
    .Y(_05161_));
 sky130_fd_sc_hd__nor2_2 _26593_ (.A(_05161_),
    .B(_05108_),
    .Y(_05162_));
 sky130_fd_sc_hd__a221o_2 _26594_ (.A1(_05105_),
    .A2(\alu_shl[31] ),
    .B1(_04994_),
    .B2(_05160_),
    .C1(_05162_),
    .X(_05163_));
 sky130_fd_sc_hd__a221o_2 _26595_ (.A1(\alu_shr[31] ),
    .A2(_05006_),
    .B1(_19711_),
    .B2(_05016_),
    .C1(_05163_),
    .X(_02165_));
 sky130_fd_sc_hd__and3_2 _26596_ (.A(_00289_),
    .B(_16858_),
    .C(_04440_),
    .X(_02166_));
 sky130_fd_sc_hd__nand2_2 _26597_ (.A(_04438_),
    .B(_04439_),
    .Y(mem_la_wstrb[0]));
 sky130_fd_sc_hd__nand2_2 _26598_ (.A(_04438_),
    .B(_04444_),
    .Y(mem_la_wstrb[1]));
 sky130_fd_sc_hd__buf_1 _26599_ (.A(_19757_),
    .X(_05164_));
 sky130_fd_sc_hd__a22o_2 _26600_ (.A1(_18430_),
    .A2(_05164_),
    .B1(_18455_),
    .B2(_04078_),
    .X(_02167_));
 sky130_fd_sc_hd__a22o_2 _26601_ (.A1(_18428_),
    .A2(_05164_),
    .B1(_18527_),
    .B2(_04078_),
    .X(_02168_));
 sky130_fd_sc_hd__a22o_2 _26602_ (.A1(_18426_),
    .A2(_05164_),
    .B1(_18526_),
    .B2(_04078_),
    .X(_02169_));
 sky130_fd_sc_hd__buf_1 _26603_ (.A(_04437_),
    .X(_05165_));
 sky130_fd_sc_hd__buf_1 _26604_ (.A(_04076_),
    .X(_05166_));
 sky130_fd_sc_hd__a22o_2 _26605_ (.A1(_18424_),
    .A2(_05165_),
    .B1(_19535_),
    .B2(_05166_),
    .X(_02170_));
 sky130_fd_sc_hd__a22o_2 _26606_ (.A1(_18421_),
    .A2(_05165_),
    .B1(_18442_),
    .B2(_05166_),
    .X(_02171_));
 sky130_fd_sc_hd__a22o_2 _26607_ (.A1(_18420_),
    .A2(_05165_),
    .B1(_18440_),
    .B2(_05166_),
    .X(_02172_));
 sky130_fd_sc_hd__a22o_2 _26608_ (.A1(_18418_),
    .A2(_05165_),
    .B1(_18437_),
    .B2(_05166_),
    .X(_02173_));
 sky130_fd_sc_hd__a22o_2 _26609_ (.A1(_18416_),
    .A2(_04593_),
    .B1(_18434_),
    .B2(_04077_),
    .X(_02174_));
 sky130_fd_sc_hd__buf_1 _26610_ (.A(_04077_),
    .X(_05167_));
 sky130_fd_sc_hd__o21a_2 _26611_ (.A1(_04577_),
    .A2(_05167_),
    .B1(_18455_),
    .X(_02175_));
 sky130_fd_sc_hd__o21a_2 _26612_ (.A1(_04577_),
    .A2(_05167_),
    .B1(_18527_),
    .X(_02176_));
 sky130_fd_sc_hd__buf_1 _26613_ (.A(_18448_),
    .X(_05168_));
 sky130_fd_sc_hd__o21a_2 _26614_ (.A1(_04577_),
    .A2(_05167_),
    .B1(_05168_),
    .X(_02177_));
 sky130_fd_sc_hd__buf_1 _26615_ (.A(_04593_),
    .X(_05169_));
 sky130_fd_sc_hd__o21a_2 _26616_ (.A1(_05169_),
    .A2(_05167_),
    .B1(_19534_),
    .X(_02178_));
 sky130_fd_sc_hd__buf_1 _26617_ (.A(_04077_),
    .X(_05170_));
 sky130_fd_sc_hd__o21a_2 _26618_ (.A1(_05169_),
    .A2(_05170_),
    .B1(_19533_),
    .X(_02179_));
 sky130_fd_sc_hd__o21a_2 _26619_ (.A1(_05169_),
    .A2(_05170_),
    .B1(_18440_),
    .X(_02180_));
 sky130_fd_sc_hd__o21a_2 _26620_ (.A1(_05169_),
    .A2(_05170_),
    .B1(_18437_),
    .X(_02181_));
 sky130_fd_sc_hd__o21a_2 _26621_ (.A1(_05164_),
    .A2(_05170_),
    .B1(_18434_),
    .X(_02182_));
 sky130_fd_sc_hd__nand2_2 _26622_ (.A(_04080_),
    .B(_16987_),
    .Y(_02183_));
 sky130_fd_sc_hd__or2_2 _26623_ (.A(_17984_),
    .B(irq[3]),
    .X(_02214_));
 sky130_fd_sc_hd__o21a_2 _26624_ (.A1(_17984_),
    .A2(irq[3]),
    .B1(_17205_),
    .X(_02215_));
 sky130_vsdinv _26625_ (.A(_01700_),
    .Y(_02217_));
 sky130_fd_sc_hd__or2_2 _26626_ (.A(_17979_),
    .B(irq[4]),
    .X(_02218_));
 sky130_fd_sc_hd__o21a_2 _26627_ (.A1(_17979_),
    .A2(irq[4]),
    .B1(_17202_),
    .X(_02219_));
 sky130_fd_sc_hd__or2_2 _26628_ (.A(_17976_),
    .B(irq[5]),
    .X(_02221_));
 sky130_fd_sc_hd__o21a_2 _26629_ (.A1(_17976_),
    .A2(irq[5]),
    .B1(_17199_),
    .X(_02222_));
 sky130_fd_sc_hd__or2_2 _26630_ (.A(_17973_),
    .B(irq[6]),
    .X(_02224_));
 sky130_fd_sc_hd__o21a_2 _26631_ (.A1(_17973_),
    .A2(irq[6]),
    .B1(_17196_),
    .X(_02225_));
 sky130_fd_sc_hd__or2_2 _26632_ (.A(_17968_),
    .B(irq[7]),
    .X(_02227_));
 sky130_fd_sc_hd__o21a_2 _26633_ (.A1(_17968_),
    .A2(irq[7]),
    .B1(\irq_mask[7] ),
    .X(_02228_));
 sky130_fd_sc_hd__or2_2 _26634_ (.A(_17962_),
    .B(irq[8]),
    .X(_02230_));
 sky130_fd_sc_hd__o21a_2 _26635_ (.A1(_17962_),
    .A2(irq[8]),
    .B1(_17187_),
    .X(_02231_));
 sky130_fd_sc_hd__or2_2 _26636_ (.A(_17959_),
    .B(irq[9]),
    .X(_02233_));
 sky130_fd_sc_hd__o21a_2 _26637_ (.A1(_17959_),
    .A2(irq[9]),
    .B1(_17183_),
    .X(_02234_));
 sky130_fd_sc_hd__or2_2 _26638_ (.A(_17956_),
    .B(irq[10]),
    .X(_02236_));
 sky130_fd_sc_hd__o21a_2 _26639_ (.A1(_17956_),
    .A2(irq[10]),
    .B1(_17180_),
    .X(_02237_));
 sky130_fd_sc_hd__or2_2 _26640_ (.A(_17951_),
    .B(irq[11]),
    .X(_02239_));
 sky130_fd_sc_hd__o21a_2 _26641_ (.A1(_17951_),
    .A2(irq[11]),
    .B1(\irq_mask[11] ),
    .X(_02240_));
 sky130_fd_sc_hd__or2_2 _26642_ (.A(_17946_),
    .B(irq[12]),
    .X(_02242_));
 sky130_fd_sc_hd__o21a_2 _26643_ (.A1(_17946_),
    .A2(irq[12]),
    .B1(_17176_),
    .X(_02243_));
 sky130_fd_sc_hd__or2_2 _26644_ (.A(_17943_),
    .B(irq[13]),
    .X(_02245_));
 sky130_fd_sc_hd__o21a_2 _26645_ (.A1(_17943_),
    .A2(irq[13]),
    .B1(_17170_),
    .X(_02246_));
 sky130_fd_sc_hd__or2_2 _26646_ (.A(_17940_),
    .B(irq[14]),
    .X(_02248_));
 sky130_fd_sc_hd__o21a_2 _26647_ (.A1(_17940_),
    .A2(irq[14]),
    .B1(_17166_),
    .X(_02249_));
 sky130_fd_sc_hd__or2_2 _26648_ (.A(_17933_),
    .B(irq[15]),
    .X(_02251_));
 sky130_fd_sc_hd__o21a_2 _26649_ (.A1(_17933_),
    .A2(irq[15]),
    .B1(_17931_),
    .X(_02252_));
 sky130_fd_sc_hd__or2_2 _26650_ (.A(_17926_),
    .B(irq[16]),
    .X(_02254_));
 sky130_fd_sc_hd__o21a_2 _26651_ (.A1(_17926_),
    .A2(irq[16]),
    .B1(_17162_),
    .X(_02255_));
 sky130_fd_sc_hd__or2_2 _26652_ (.A(_17923_),
    .B(irq[17]),
    .X(_02257_));
 sky130_fd_sc_hd__o21a_2 _26653_ (.A1(_17923_),
    .A2(irq[17]),
    .B1(_17159_),
    .X(_02258_));
 sky130_fd_sc_hd__or2_2 _26654_ (.A(_17920_),
    .B(irq[18]),
    .X(_02260_));
 sky130_fd_sc_hd__o21a_2 _26655_ (.A1(_17920_),
    .A2(irq[18]),
    .B1(_17157_),
    .X(_02261_));
 sky130_fd_sc_hd__or2_2 _26656_ (.A(_17915_),
    .B(irq[19]),
    .X(_02263_));
 sky130_fd_sc_hd__o21a_2 _26657_ (.A1(_17915_),
    .A2(irq[19]),
    .B1(_17154_),
    .X(_02264_));
 sky130_fd_sc_hd__or2_2 _26658_ (.A(_17910_),
    .B(irq[20]),
    .X(_02266_));
 sky130_fd_sc_hd__o21a_2 _26659_ (.A1(_17910_),
    .A2(irq[20]),
    .B1(_17151_),
    .X(_02267_));
 sky130_fd_sc_hd__or2_2 _26660_ (.A(_17907_),
    .B(irq[21]),
    .X(_02269_));
 sky130_fd_sc_hd__o21a_2 _26661_ (.A1(_17907_),
    .A2(irq[21]),
    .B1(_17146_),
    .X(_02270_));
 sky130_fd_sc_hd__or2_2 _26662_ (.A(_17904_),
    .B(irq[22]),
    .X(_02272_));
 sky130_fd_sc_hd__o21a_2 _26663_ (.A1(_17904_),
    .A2(irq[22]),
    .B1(_17143_),
    .X(_02273_));
 sky130_fd_sc_hd__or2_2 _26664_ (.A(_17899_),
    .B(irq[23]),
    .X(_02275_));
 sky130_fd_sc_hd__o21a_2 _26665_ (.A1(_17899_),
    .A2(irq[23]),
    .B1(_17896_),
    .X(_02276_));
 sky130_fd_sc_hd__or2_2 _26666_ (.A(_17892_),
    .B(irq[24]),
    .X(_02278_));
 sky130_fd_sc_hd__o21a_2 _26667_ (.A1(_17892_),
    .A2(irq[24]),
    .B1(_17134_),
    .X(_02279_));
 sky130_fd_sc_hd__or2_2 _26668_ (.A(_17889_),
    .B(irq[25]),
    .X(_02281_));
 sky130_fd_sc_hd__o21a_2 _26669_ (.A1(_17889_),
    .A2(irq[25]),
    .B1(_17129_),
    .X(_02282_));
 sky130_fd_sc_hd__or2_2 _26670_ (.A(_17886_),
    .B(irq[26]),
    .X(_02284_));
 sky130_fd_sc_hd__o21a_2 _26671_ (.A1(_17886_),
    .A2(irq[26]),
    .B1(_17126_),
    .X(_02285_));
 sky130_fd_sc_hd__or2_2 _26672_ (.A(_17881_),
    .B(irq[27]),
    .X(_02287_));
 sky130_fd_sc_hd__o21a_2 _26673_ (.A1(_17881_),
    .A2(irq[27]),
    .B1(\irq_mask[27] ),
    .X(_02288_));
 sky130_fd_sc_hd__or2_2 _26674_ (.A(_17876_),
    .B(irq[28]),
    .X(_02290_));
 sky130_fd_sc_hd__o21a_2 _26675_ (.A1(_17876_),
    .A2(irq[28]),
    .B1(_17116_),
    .X(_02291_));
 sky130_fd_sc_hd__or2_2 _26676_ (.A(_17873_),
    .B(irq[29]),
    .X(_02293_));
 sky130_fd_sc_hd__o21a_2 _26677_ (.A1(_17873_),
    .A2(irq[29]),
    .B1(_17113_),
    .X(_02294_));
 sky130_fd_sc_hd__or2_2 _26678_ (.A(_17870_),
    .B(irq[30]),
    .X(_02296_));
 sky130_fd_sc_hd__o21a_2 _26679_ (.A1(_17870_),
    .A2(irq[30]),
    .B1(_17108_),
    .X(_02297_));
 sky130_fd_sc_hd__or2_2 _26680_ (.A(_17861_),
    .B(irq[31]),
    .X(_02299_));
 sky130_fd_sc_hd__o21a_2 _26681_ (.A1(_17861_),
    .A2(irq[31]),
    .B1(_17088_),
    .X(_02300_));
 sky130_fd_sc_hd__or4_2 _26682_ (.A(\timer[23] ),
    .B(\timer[22] ),
    .C(\timer[31] ),
    .D(\timer[30] ),
    .X(_05171_));
 sky130_fd_sc_hd__or4_2 _26683_ (.A(_04113_),
    .B(_04117_),
    .C(\timer[15] ),
    .D(\timer[14] ),
    .X(_05172_));
 sky130_fd_sc_hd__or4_2 _26684_ (.A(_04086_),
    .B(_04083_),
    .C(_05171_),
    .D(_05172_),
    .X(_05173_));
 sky130_fd_sc_hd__nand3b_2 _26685_ (.A_N(_04103_),
    .B(_04100_),
    .C(\timer[0] ),
    .Y(_05174_));
 sky130_fd_sc_hd__or4_2 _26686_ (.A(\timer[3] ),
    .B(_04104_),
    .C(_04111_),
    .D(\timer[6] ),
    .X(_05175_));
 sky130_fd_sc_hd__nand3b_2 _26687_ (.A_N(_05175_),
    .B(_04094_),
    .C(_04090_),
    .Y(_05176_));
 sky130_fd_sc_hd__or4_2 _26688_ (.A(_04087_),
    .B(_04130_),
    .C(_05174_),
    .D(_05176_),
    .X(_05177_));
 sky130_fd_sc_hd__o21bai_2 _26689_ (.A1(_05173_),
    .A2(_05177_),
    .B1_N(\irq_pending[0] ),
    .Y(_02302_));
 sky130_fd_sc_hd__or2_2 _26690_ (.A(_02303_),
    .B(irq[0]),
    .X(_02304_));
 sky130_fd_sc_hd__o21a_2 _26691_ (.A1(_02303_),
    .A2(irq[0]),
    .B1(_17214_),
    .X(_02305_));
 sky130_fd_sc_hd__nor2_2 _26692_ (.A(_17991_),
    .B(irq[2]),
    .Y(_02307_));
 sky130_fd_sc_hd__o21ai_2 _26693_ (.A1(_17991_),
    .A2(irq[2]),
    .B1(_19549_),
    .Y(_02308_));
 sky130_fd_sc_hd__nor2b_2 _26694_ (.A(_02310_),
    .B_N(_16832_),
    .Y(_02311_));
 sky130_fd_sc_hd__o22ai_2 _26695_ (.A1(_16936_),
    .A2(_17990_),
    .B1(_02310_),
    .B2(_17370_),
    .Y(_02312_));
 sky130_fd_sc_hd__o21bai_2 _26696_ (.A1(_19548_),
    .A2(_19549_),
    .B1_N(_02313_),
    .Y(_02314_));
 sky130_fd_sc_hd__o21bai_2 _26697_ (.A1(_19548_),
    .A2(_19549_),
    .B1_N(_02316_),
    .Y(_02317_));
 sky130_fd_sc_hd__and2b_2 _26698_ (.A_N(_16958_),
    .B(_16977_),
    .X(_05178_));
 sky130_fd_sc_hd__and2b_2 _26699_ (.A_N(_19076_),
    .B(_18415_),
    .X(_05179_));
 sky130_fd_sc_hd__and2b_2 _26700_ (.A_N(_19080_),
    .B(pcpi_rs2[14]),
    .X(_05180_));
 sky130_fd_sc_hd__and2b_2 _26701_ (.A_N(_19082_),
    .B(_18419_),
    .X(_05181_));
 sky130_fd_sc_hd__inv_2 _26702_ (.A(pcpi_rs2[12]),
    .Y(_02351_));
 sky130_fd_sc_hd__nor3_2 _26703_ (.A(_02351_),
    .B(_19084_),
    .C(_19724_),
    .Y(_05182_));
 sky130_fd_sc_hd__o21ba_2 _26704_ (.A1(_05181_),
    .A2(_05182_),
    .B1_N(_19725_),
    .X(_05183_));
 sky130_fd_sc_hd__o21ba_2 _26705_ (.A1(_05180_),
    .A2(_05183_),
    .B1_N(_19722_),
    .X(_05184_));
 sky130_fd_sc_hd__and2b_2 _26706_ (.A_N(_19098_),
    .B(_18432_),
    .X(_05185_));
 sky130_fd_sc_hd__inv_2 _26707_ (.A(_18438_),
    .Y(_02330_));
 sky130_vsdinv _26708_ (.A(_19736_),
    .Y(_05186_));
 sky130_fd_sc_hd__a211oi_2 _26709_ (.A1(_05186_),
    .A2(_05045_),
    .B1(_19537_),
    .C1(_19107_),
    .Y(_05187_));
 sky130_fd_sc_hd__o21bai_2 _26710_ (.A1(_02330_),
    .A2(_19105_),
    .B1_N(_05187_),
    .Y(_05188_));
 sky130_fd_sc_hd__o21a_2 _26711_ (.A1(_19541_),
    .A2(_00048_),
    .B1(_19115_),
    .X(_05189_));
 sky130_fd_sc_hd__a211o_2 _26712_ (.A1(_19541_),
    .A2(_00048_),
    .B1(_05189_),
    .C1(_19732_),
    .X(_05190_));
 sky130_fd_sc_hd__nand3_2 _26713_ (.A(_19727_),
    .B(_18447_),
    .C(_19728_),
    .Y(_05191_));
 sky130_fd_sc_hd__or2b_2 _26714_ (.A(_19109_),
    .B_N(_18444_),
    .X(_05192_));
 sky130_fd_sc_hd__a31oi_2 _26715_ (.A1(_05190_),
    .A2(_05191_),
    .A3(_05192_),
    .B1(_19737_),
    .Y(_05193_));
 sky130_fd_sc_hd__o21bai_2 _26716_ (.A1(_05188_),
    .A2(_05193_),
    .B1_N(_05050_),
    .Y(_05194_));
 sky130_fd_sc_hd__nand2_2 _26717_ (.A(_19738_),
    .B(_18436_),
    .Y(_05195_));
 sky130_fd_sc_hd__a21oi_2 _26718_ (.A1(_05194_),
    .A2(_05195_),
    .B1(_19742_),
    .Y(_05196_));
 sky130_fd_sc_hd__o21ai_2 _26719_ (.A1(_05185_),
    .A2(_05196_),
    .B1(_19754_),
    .Y(_05197_));
 sky130_fd_sc_hd__or2b_2 _26720_ (.A(_19087_),
    .B_N(_18423_),
    .X(_05198_));
 sky130_fd_sc_hd__or2b_2 _26721_ (.A(_19089_),
    .B_N(pcpi_rs2[10]),
    .X(_05199_));
 sky130_fd_sc_hd__and2b_2 _26722_ (.A_N(_19092_),
    .B(pcpi_rs2[9]),
    .X(_05200_));
 sky130_vsdinv _26723_ (.A(_19095_),
    .Y(_05201_));
 sky130_fd_sc_hd__and3_2 _26724_ (.A(_19747_),
    .B(_18429_),
    .C(_05201_),
    .X(_05202_));
 sky130_fd_sc_hd__o21bai_2 _26725_ (.A1(_05200_),
    .A2(_05202_),
    .B1_N(_19752_),
    .Y(_05203_));
 sky130_fd_sc_hd__o2bb2ai_2 _26726_ (.A1_N(_05199_),
    .A2_N(_05203_),
    .B1(_19749_),
    .B2(_19748_),
    .Y(_05204_));
 sky130_fd_sc_hd__a31oi_2 _26727_ (.A1(_05197_),
    .A2(_05198_),
    .A3(_05204_),
    .B1(_19726_),
    .Y(_05205_));
 sky130_fd_sc_hd__o31ai_2 _26728_ (.A1(_05179_),
    .A2(_05184_),
    .A3(_05205_),
    .B1(_19721_),
    .Y(_05206_));
 sky130_fd_sc_hd__o2bb2ai_2 _26729_ (.A1_N(_05161_),
    .A2_N(_05160_),
    .B1(_19709_),
    .B2(_19710_),
    .Y(_05207_));
 sky130_fd_sc_hd__inv_2 _26730_ (.A(pcpi_rs2[27]),
    .Y(_02396_));
 sky130_fd_sc_hd__and2b_2 _26731_ (.A_N(_19701_),
    .B(pcpi_rs2[26]),
    .X(_05208_));
 sky130_vsdinv _26732_ (.A(_19707_),
    .Y(_05209_));
 sky130_fd_sc_hd__inv_2 _26733_ (.A(pcpi_rs2[24]),
    .Y(_02387_));
 sky130_fd_sc_hd__a211o_2 _26734_ (.A1(_05209_),
    .A2(_05139_),
    .B1(_02387_),
    .C1(_19054_),
    .X(_05210_));
 sky130_fd_sc_hd__nand2_2 _26735_ (.A(_04257_),
    .B(_18394_),
    .Y(_05211_));
 sky130_fd_sc_hd__a21oi_2 _26736_ (.A1(_05210_),
    .A2(_05211_),
    .B1(_19702_),
    .Y(_05212_));
 sky130_fd_sc_hd__o21bai_2 _26737_ (.A1(_05208_),
    .A2(_05212_),
    .B1_N(_19700_),
    .Y(_05213_));
 sky130_fd_sc_hd__o21ai_2 _26738_ (.A1(_02396_),
    .A2(_19047_),
    .B1(_05213_),
    .Y(_05214_));
 sky130_fd_sc_hd__o211a_2 _26739_ (.A1(_19714_),
    .A2(_19713_),
    .B1(pcpi_rs2[28]),
    .C1(_19715_),
    .X(_05215_));
 sky130_fd_sc_hd__a221oi_2 _26740_ (.A1(_18386_),
    .A2(_04278_),
    .B1(_05214_),
    .B2(_19718_),
    .C1(_05215_),
    .Y(_05216_));
 sky130_fd_sc_hd__inv_2 _26741_ (.A(pcpi_rs2[30]),
    .Y(_02405_));
 sky130_fd_sc_hd__a211o_2 _26742_ (.A1(_05160_),
    .A2(_05161_),
    .B1(_02405_),
    .C1(_19041_),
    .X(_05217_));
 sky130_fd_sc_hd__and2b_2 _26743_ (.A_N(_19068_),
    .B(_18408_),
    .X(_05218_));
 sky130_fd_sc_hd__and2b_2 _26744_ (.A_N(_19071_),
    .B(_18410_),
    .X(_05219_));
 sky130_fd_sc_hd__inv_2 _26745_ (.A(pcpi_rs2[16]),
    .Y(_02363_));
 sky130_fd_sc_hd__nor3_2 _26746_ (.A(_02363_),
    .B(_19073_),
    .C(_19697_),
    .Y(_05220_));
 sky130_fd_sc_hd__o21ba_2 _26747_ (.A1(_05219_),
    .A2(_05220_),
    .B1_N(_19698_),
    .X(_05221_));
 sky130_fd_sc_hd__o21bai_2 _26748_ (.A1(_05218_),
    .A2(_05221_),
    .B1_N(_19695_),
    .Y(_05222_));
 sky130_fd_sc_hd__or2b_2 _26749_ (.A(_19065_),
    .B_N(_18406_),
    .X(_05223_));
 sky130_fd_sc_hd__a21o_2 _26750_ (.A1(_05222_),
    .A2(_05223_),
    .B1(_19694_),
    .X(_05224_));
 sky130_fd_sc_hd__or2b_2 _26751_ (.A(_19056_),
    .B_N(_18398_),
    .X(_05225_));
 sky130_fd_sc_hd__and2b_2 _26752_ (.A_N(_19059_),
    .B(pcpi_rs2[22]),
    .X(_05226_));
 sky130_fd_sc_hd__and2b_2 _26753_ (.A_N(_19061_),
    .B(_18402_),
    .X(_05227_));
 sky130_fd_sc_hd__inv_2 _26754_ (.A(pcpi_rs2[20]),
    .Y(_02375_));
 sky130_fd_sc_hd__nor3_2 _26755_ (.A(_02375_),
    .B(_19063_),
    .C(_19692_),
    .Y(_05228_));
 sky130_fd_sc_hd__o21ba_2 _26756_ (.A1(_05227_),
    .A2(_05228_),
    .B1_N(_19693_),
    .X(_05229_));
 sky130_fd_sc_hd__o21bai_2 _26757_ (.A1(_05226_),
    .A2(_05229_),
    .B1_N(_19690_),
    .Y(_05230_));
 sky130_fd_sc_hd__a31o_2 _26758_ (.A1(_05224_),
    .A2(_05225_),
    .A3(_05230_),
    .B1(_19720_),
    .X(_05231_));
 sky130_fd_sc_hd__o211a_2 _26759_ (.A1(_05207_),
    .A2(_05216_),
    .B1(_05217_),
    .C1(_05231_),
    .X(_05232_));
 sky130_fd_sc_hd__and3b_2 _26760_ (.A_N(_05178_),
    .B(_05206_),
    .C(_05232_),
    .X(_05233_));
 sky130_fd_sc_hd__nor2_2 _26761_ (.A(_00000_),
    .B(_05233_),
    .Y(_00002_));
 sky130_fd_sc_hd__a31oi_2 _26762_ (.A1(_05206_),
    .A2(_19712_),
    .A3(_05232_),
    .B1(_00000_),
    .Y(_05234_));
 sky130_fd_sc_hd__o21a_2 _26763_ (.A1(_19712_),
    .A2(_05233_),
    .B1(_05234_),
    .X(_00001_));
 sky130_fd_sc_hd__buf_1 _26764_ (.A(\pcpi_mul.rs2[0] ),
    .X(_05235_));
 sky130_fd_sc_hd__buf_1 _26765_ (.A(_05235_),
    .X(_05236_));
 sky130_fd_sc_hd__buf_1 _26766_ (.A(_05236_),
    .X(_05237_));
 sky130_fd_sc_hd__buf_1 _26767_ (.A(\pcpi_mul.rs1[0] ),
    .X(_05238_));
 sky130_fd_sc_hd__buf_1 _26768_ (.A(_05238_),
    .X(_05239_));
 sky130_fd_sc_hd__buf_1 _26769_ (.A(_05239_),
    .X(_05240_));
 sky130_fd_sc_hd__buf_1 _26770_ (.A(_05240_),
    .X(_05241_));
 sky130_fd_sc_hd__buf_1 _26771_ (.A(_05241_),
    .X(_05242_));
 sky130_fd_sc_hd__buf_1 _26772_ (.A(_05242_),
    .X(_05243_));
 sky130_fd_sc_hd__and2_2 _26773_ (.A(_05237_),
    .B(_05243_),
    .X(_02623_));
 sky130_fd_sc_hd__xnor2_2 _26774_ (.A(_18451_),
    .B(_18454_),
    .Y(_02319_));
 sky130_fd_sc_hd__and2b_2 _26775_ (.A_N(pcpi_rs1[0]),
    .B(mem_la_wdata[0]),
    .X(_05244_));
 sky130_vsdinv _26776_ (.A(_05244_),
    .Y(_05245_));
 sky130_fd_sc_hd__xor2_2 _26777_ (.A(pcpi_rs1[1]),
    .B(_02320_),
    .X(_05246_));
 sky130_fd_sc_hd__xor2_2 _26778_ (.A(_05245_),
    .B(_05246_),
    .X(_02602_));
 sky130_vsdinv _26779_ (.A(_18453_),
    .Y(_05247_));
 sky130_fd_sc_hd__nand2_2 _26780_ (.A(_19541_),
    .B(_05247_),
    .Y(_05248_));
 sky130_fd_sc_hd__xor2_2 _26781_ (.A(_19539_),
    .B(_05248_),
    .X(_02322_));
 sky130_fd_sc_hd__xor2_2 _26782_ (.A(_19113_),
    .B(_02323_),
    .X(_05249_));
 sky130_fd_sc_hd__and2_2 _26783_ (.A(_19114_),
    .B(_02320_),
    .X(_05250_));
 sky130_fd_sc_hd__a21o_2 _26784_ (.A1(_05246_),
    .A2(_05245_),
    .B1(_05250_),
    .X(_05251_));
 sky130_fd_sc_hd__xor2_2 _26785_ (.A(_05249_),
    .B(_05251_),
    .X(_02613_));
 sky130_fd_sc_hd__nor3_2 _26786_ (.A(mem_la_wdata[2]),
    .B(mem_la_wdata[1]),
    .C(_18452_),
    .Y(_05252_));
 sky130_fd_sc_hd__xor2_2 _26787_ (.A(_18446_),
    .B(_05252_),
    .X(_02325_));
 sky130_fd_sc_hd__nor2_2 _26788_ (.A(pcpi_rs1[3]),
    .B(_02326_),
    .Y(_05253_));
 sky130_fd_sc_hd__and2_2 _26789_ (.A(pcpi_rs1[3]),
    .B(_02326_),
    .X(_05254_));
 sky130_fd_sc_hd__nor2_2 _26790_ (.A(_05253_),
    .B(_05254_),
    .Y(_05255_));
 sky130_fd_sc_hd__o21ai_2 _26791_ (.A1(pcpi_rs1[2]),
    .A2(_02323_),
    .B1(_05251_),
    .Y(_05256_));
 sky130_fd_sc_hd__nand2_2 _26792_ (.A(pcpi_rs1[2]),
    .B(_02323_),
    .Y(_05257_));
 sky130_fd_sc_hd__nand2_2 _26793_ (.A(_05256_),
    .B(_05257_),
    .Y(_05258_));
 sky130_fd_sc_hd__xor2_2 _26794_ (.A(_05255_),
    .B(_05258_),
    .X(_02616_));
 sky130_fd_sc_hd__nand2_2 _26795_ (.A(_05252_),
    .B(_19542_),
    .Y(_05259_));
 sky130_fd_sc_hd__xor2_2 _26796_ (.A(_19537_),
    .B(_05259_),
    .X(_02328_));
 sky130_fd_sc_hd__xor2_2 _26797_ (.A(_19108_),
    .B(_02329_),
    .X(_05260_));
 sky130_vsdinv _26798_ (.A(_05253_),
    .Y(_05261_));
 sky130_fd_sc_hd__a21o_2 _26799_ (.A1(_05258_),
    .A2(_05261_),
    .B1(_05254_),
    .X(_05262_));
 sky130_fd_sc_hd__xor2_2 _26800_ (.A(_05260_),
    .B(_05262_),
    .X(_02617_));
 sky130_fd_sc_hd__nand3_2 _26801_ (.A(_05252_),
    .B(_19536_),
    .C(_19538_),
    .Y(_05263_));
 sky130_fd_sc_hd__xor2_2 _26802_ (.A(_02330_),
    .B(_05263_),
    .X(_02331_));
 sky130_fd_sc_hd__nor2_2 _26803_ (.A(pcpi_rs1[5]),
    .B(_02332_),
    .Y(_05264_));
 sky130_fd_sc_hd__and2_2 _26804_ (.A(pcpi_rs1[5]),
    .B(_02332_),
    .X(_05265_));
 sky130_fd_sc_hd__nor2_2 _26805_ (.A(_05264_),
    .B(_05265_),
    .Y(_05266_));
 sky130_fd_sc_hd__or2_2 _26806_ (.A(pcpi_rs1[4]),
    .B(_02329_),
    .X(_05267_));
 sky130_fd_sc_hd__nand2_2 _26807_ (.A(_05262_),
    .B(_05267_),
    .Y(_05268_));
 sky130_fd_sc_hd__nand2_2 _26808_ (.A(_19106_),
    .B(_02329_),
    .Y(_05269_));
 sky130_fd_sc_hd__nand2_2 _26809_ (.A(_05268_),
    .B(_05269_),
    .Y(_05270_));
 sky130_fd_sc_hd__xor2_2 _26810_ (.A(_05266_),
    .B(_05270_),
    .X(_02618_));
 sky130_fd_sc_hd__nor2_2 _26811_ (.A(_18439_),
    .B(_05263_),
    .Y(_05271_));
 sky130_fd_sc_hd__xor2_2 _26812_ (.A(_18436_),
    .B(_05271_),
    .X(_02334_));
 sky130_fd_sc_hd__xor2_2 _26813_ (.A(pcpi_rs1[6]),
    .B(_02335_),
    .X(_05272_));
 sky130_vsdinv _26814_ (.A(_05264_),
    .Y(_05273_));
 sky130_fd_sc_hd__a21o_2 _26815_ (.A1(_05270_),
    .A2(_05273_),
    .B1(_05265_),
    .X(_05274_));
 sky130_fd_sc_hd__xor2_2 _26816_ (.A(_05272_),
    .B(_05274_),
    .X(_02619_));
 sky130_fd_sc_hd__inv_2 _26817_ (.A(mem_la_wdata[7]),
    .Y(_02336_));
 sky130_fd_sc_hd__nor3_2 _26818_ (.A(mem_la_wdata[6]),
    .B(mem_la_wdata[5]),
    .C(_05263_),
    .Y(_05275_));
 sky130_fd_sc_hd__xor2_2 _26819_ (.A(_18433_),
    .B(_05275_),
    .X(_02337_));
 sky130_fd_sc_hd__xnor2_2 _26820_ (.A(pcpi_rs1[7]),
    .B(_02338_),
    .Y(_05276_));
 sky130_fd_sc_hd__nand2_2 _26821_ (.A(_05274_),
    .B(_05272_),
    .Y(_05277_));
 sky130_fd_sc_hd__a21boi_2 _26822_ (.A1(_19103_),
    .A2(_02335_),
    .B1_N(_05277_),
    .Y(_05278_));
 sky130_fd_sc_hd__xor2_2 _26823_ (.A(_05276_),
    .B(_05278_),
    .X(_02620_));
 sky130_fd_sc_hd__inv_2 _26824_ (.A(pcpi_rs2[8]),
    .Y(_02339_));
 sky130_fd_sc_hd__nand3_2 _26825_ (.A(_05271_),
    .B(_02336_),
    .C(_02333_),
    .Y(_05279_));
 sky130_fd_sc_hd__xor2_2 _26826_ (.A(_02339_),
    .B(_05279_),
    .X(_02340_));
 sky130_fd_sc_hd__xor2_2 _26827_ (.A(pcpi_rs1[8]),
    .B(_02341_),
    .X(_05280_));
 sky130_fd_sc_hd__and2b_2 _26828_ (.A_N(_05276_),
    .B(_05272_),
    .X(_05281_));
 sky130_fd_sc_hd__nand2_2 _26829_ (.A(_05274_),
    .B(_05281_),
    .Y(_05282_));
 sky130_fd_sc_hd__o211a_2 _26830_ (.A1(_19097_),
    .A2(_02338_),
    .B1(_19101_),
    .C1(_02335_),
    .X(_05283_));
 sky130_fd_sc_hd__a21oi_2 _26831_ (.A1(_19098_),
    .A2(_02338_),
    .B1(_05283_),
    .Y(_05284_));
 sky130_fd_sc_hd__nand2_2 _26832_ (.A(_05282_),
    .B(_05284_),
    .Y(_05285_));
 sky130_fd_sc_hd__xor2_2 _26833_ (.A(_05280_),
    .B(_05285_),
    .X(_02621_));
 sky130_fd_sc_hd__inv_2 _26834_ (.A(_18428_),
    .Y(_02342_));
 sky130_fd_sc_hd__nand3_2 _26835_ (.A(_05275_),
    .B(_02339_),
    .C(_02336_),
    .Y(_05286_));
 sky130_fd_sc_hd__xor2_2 _26836_ (.A(_02342_),
    .B(_05286_),
    .X(_02343_));
 sky130_fd_sc_hd__xnor2_2 _26837_ (.A(pcpi_rs1[9]),
    .B(_02344_),
    .Y(_05287_));
 sky130_fd_sc_hd__a21boi_2 _26838_ (.A1(_05282_),
    .A2(_05284_),
    .B1_N(_05280_),
    .Y(_05288_));
 sky130_fd_sc_hd__a21oi_2 _26839_ (.A1(_19096_),
    .A2(_02341_),
    .B1(_05288_),
    .Y(_05289_));
 sky130_fd_sc_hd__xor2_2 _26840_ (.A(_05287_),
    .B(_05289_),
    .X(_02622_));
 sky130_fd_sc_hd__inv_2 _26841_ (.A(_18425_),
    .Y(_02345_));
 sky130_fd_sc_hd__nor2_2 _26842_ (.A(_18427_),
    .B(_05286_),
    .Y(_05290_));
 sky130_fd_sc_hd__xor2_2 _26843_ (.A(_18426_),
    .B(_05290_),
    .X(_02346_));
 sky130_fd_sc_hd__nor2_2 _26844_ (.A(pcpi_rs1[10]),
    .B(_02347_),
    .Y(_05291_));
 sky130_fd_sc_hd__and2_2 _26845_ (.A(pcpi_rs1[10]),
    .B(_02347_),
    .X(_05292_));
 sky130_fd_sc_hd__nor2_2 _26846_ (.A(_05291_),
    .B(_05292_),
    .Y(_05293_));
 sky130_fd_sc_hd__and2b_2 _26847_ (.A_N(_05287_),
    .B(_05280_),
    .X(_05294_));
 sky130_fd_sc_hd__nand2_2 _26848_ (.A(_05285_),
    .B(_05294_),
    .Y(_05295_));
 sky130_fd_sc_hd__o211a_2 _26849_ (.A1(_19091_),
    .A2(_02344_),
    .B1(_19094_),
    .C1(_02341_),
    .X(_05296_));
 sky130_fd_sc_hd__a21oi_2 _26850_ (.A1(_19092_),
    .A2(_02344_),
    .B1(_05296_),
    .Y(_05297_));
 sky130_fd_sc_hd__nand2_2 _26851_ (.A(_05295_),
    .B(_05297_),
    .Y(_05298_));
 sky130_fd_sc_hd__xor2_2 _26852_ (.A(_05293_),
    .B(_05298_),
    .X(_02592_));
 sky130_fd_sc_hd__inv_2 _26853_ (.A(pcpi_rs2[11]),
    .Y(_02348_));
 sky130_fd_sc_hd__nor3_2 _26854_ (.A(pcpi_rs2[10]),
    .B(pcpi_rs2[9]),
    .C(_05286_),
    .Y(_05299_));
 sky130_fd_sc_hd__xor2_2 _26855_ (.A(_18424_),
    .B(_05299_),
    .X(_02349_));
 sky130_fd_sc_hd__xnor2_2 _26856_ (.A(pcpi_rs1[11]),
    .B(_02350_),
    .Y(_05300_));
 sky130_fd_sc_hd__a21oi_2 _26857_ (.A1(_05298_),
    .A2(_05293_),
    .B1(_05292_),
    .Y(_05301_));
 sky130_fd_sc_hd__xor2_2 _26858_ (.A(_05300_),
    .B(_05301_),
    .X(_02593_));
 sky130_fd_sc_hd__nand3_2 _26859_ (.A(_05290_),
    .B(_02348_),
    .C(_02345_),
    .Y(_05302_));
 sky130_fd_sc_hd__xor2_2 _26860_ (.A(_02351_),
    .B(_05302_),
    .X(_02352_));
 sky130_fd_sc_hd__nor2_2 _26861_ (.A(pcpi_rs1[12]),
    .B(_02353_),
    .Y(_05303_));
 sky130_fd_sc_hd__and2_2 _26862_ (.A(pcpi_rs1[12]),
    .B(_02353_),
    .X(_05304_));
 sky130_fd_sc_hd__nor2_2 _26863_ (.A(_05303_),
    .B(_05304_),
    .Y(_05305_));
 sky130_fd_sc_hd__and2_2 _26864_ (.A(_19086_),
    .B(_02350_),
    .X(_05306_));
 sky130_fd_sc_hd__o21bai_2 _26865_ (.A1(_05300_),
    .A2(_05301_),
    .B1_N(_05306_),
    .Y(_05307_));
 sky130_fd_sc_hd__xor2_2 _26866_ (.A(_05305_),
    .B(_05307_),
    .X(_02594_));
 sky130_fd_sc_hd__nand3_2 _26867_ (.A(_05299_),
    .B(_02351_),
    .C(_02348_),
    .Y(_05308_));
 sky130_fd_sc_hd__xor2_2 _26868_ (.A(_02354_),
    .B(_05308_),
    .X(_02355_));
 sky130_fd_sc_hd__xnor2_2 _26869_ (.A(pcpi_rs1[13]),
    .B(_02356_),
    .Y(_05309_));
 sky130_fd_sc_hd__a21oi_2 _26870_ (.A1(_05307_),
    .A2(_05305_),
    .B1(_05304_),
    .Y(_05310_));
 sky130_fd_sc_hd__xor2_2 _26871_ (.A(_05309_),
    .B(_05310_),
    .X(_02595_));
 sky130_fd_sc_hd__inv_2 _26872_ (.A(_18417_),
    .Y(_02357_));
 sky130_fd_sc_hd__nor2_2 _26873_ (.A(_18419_),
    .B(_05308_),
    .Y(_05311_));
 sky130_fd_sc_hd__xor2_2 _26874_ (.A(_18418_),
    .B(_05311_),
    .X(_02358_));
 sky130_fd_sc_hd__nor2_2 _26875_ (.A(pcpi_rs1[14]),
    .B(_02359_),
    .Y(_05312_));
 sky130_fd_sc_hd__and2_2 _26876_ (.A(pcpi_rs1[14]),
    .B(_02359_),
    .X(_05313_));
 sky130_fd_sc_hd__nor2_2 _26877_ (.A(_05312_),
    .B(_05313_),
    .Y(_05314_));
 sky130_fd_sc_hd__and2_2 _26878_ (.A(_19082_),
    .B(_02356_),
    .X(_05315_));
 sky130_fd_sc_hd__o21bai_2 _26879_ (.A1(_05309_),
    .A2(_05310_),
    .B1_N(_05315_),
    .Y(_05316_));
 sky130_fd_sc_hd__xor2_2 _26880_ (.A(_05314_),
    .B(_05316_),
    .X(_02596_));
 sky130_fd_sc_hd__inv_2 _26881_ (.A(pcpi_rs2[15]),
    .Y(_02360_));
 sky130_fd_sc_hd__nor3_2 _26882_ (.A(pcpi_rs2[14]),
    .B(pcpi_rs2[13]),
    .C(_05308_),
    .Y(_05317_));
 sky130_fd_sc_hd__xor2_2 _26883_ (.A(_18416_),
    .B(_05317_),
    .X(_02361_));
 sky130_fd_sc_hd__xnor2_2 _26884_ (.A(pcpi_rs1[15]),
    .B(_02362_),
    .Y(_05318_));
 sky130_fd_sc_hd__a21oi_2 _26885_ (.A1(_05316_),
    .A2(_05314_),
    .B1(_05313_),
    .Y(_05319_));
 sky130_fd_sc_hd__xor2_2 _26886_ (.A(_05318_),
    .B(_05319_),
    .X(_02597_));
 sky130_fd_sc_hd__nand3_2 _26887_ (.A(_05311_),
    .B(_02360_),
    .C(_02357_),
    .Y(_05320_));
 sky130_fd_sc_hd__xor2_2 _26888_ (.A(_02363_),
    .B(_05320_),
    .X(_02364_));
 sky130_fd_sc_hd__xor2_2 _26889_ (.A(pcpi_rs1[16]),
    .B(_02365_),
    .X(_05321_));
 sky130_fd_sc_hd__and2_2 _26890_ (.A(_19076_),
    .B(_02362_),
    .X(_05322_));
 sky130_fd_sc_hd__o21bai_2 _26891_ (.A1(_05318_),
    .A2(_05319_),
    .B1_N(_05322_),
    .Y(_05323_));
 sky130_fd_sc_hd__xor2_2 _26892_ (.A(_05321_),
    .B(_05323_),
    .X(_02598_));
 sky130_fd_sc_hd__nand3_2 _26893_ (.A(_05317_),
    .B(_02363_),
    .C(_02360_),
    .Y(_05324_));
 sky130_fd_sc_hd__xor2_2 _26894_ (.A(_02366_),
    .B(_05324_),
    .X(_02367_));
 sky130_fd_sc_hd__xnor2_2 _26895_ (.A(pcpi_rs1[17]),
    .B(_02368_),
    .Y(_05325_));
 sky130_fd_sc_hd__nand2_2 _26896_ (.A(_05323_),
    .B(_05321_),
    .Y(_05326_));
 sky130_fd_sc_hd__a21boi_2 _26897_ (.A1(_19075_),
    .A2(_02365_),
    .B1_N(_05326_),
    .Y(_05327_));
 sky130_fd_sc_hd__xor2_2 _26898_ (.A(_05325_),
    .B(_05327_),
    .X(_02599_));
 sky130_fd_sc_hd__inv_2 _26899_ (.A(_18409_),
    .Y(_02369_));
 sky130_fd_sc_hd__nor2_2 _26900_ (.A(_18411_),
    .B(_05324_),
    .Y(_05328_));
 sky130_fd_sc_hd__xor2_2 _26901_ (.A(_18409_),
    .B(_05328_),
    .X(_02370_));
 sky130_fd_sc_hd__xnor2_2 _26902_ (.A(pcpi_rs1[18]),
    .B(_02371_),
    .Y(_05329_));
 sky130_fd_sc_hd__and2b_2 _26903_ (.A_N(_05325_),
    .B(_05321_),
    .X(_05330_));
 sky130_fd_sc_hd__o211a_2 _26904_ (.A1(_19070_),
    .A2(_02368_),
    .B1(_19073_),
    .C1(_02365_),
    .X(_05331_));
 sky130_fd_sc_hd__a21o_2 _26905_ (.A1(_19071_),
    .A2(_02368_),
    .B1(_05331_),
    .X(_05332_));
 sky130_fd_sc_hd__a21oi_2 _26906_ (.A1(_05323_),
    .A2(_05330_),
    .B1(_05332_),
    .Y(_05333_));
 sky130_fd_sc_hd__xor2_2 _26907_ (.A(_05329_),
    .B(_05333_),
    .X(_02600_));
 sky130_fd_sc_hd__inv_2 _26908_ (.A(pcpi_rs2[19]),
    .Y(_02372_));
 sky130_fd_sc_hd__nor3_2 _26909_ (.A(pcpi_rs2[18]),
    .B(_18410_),
    .C(_05324_),
    .Y(_05334_));
 sky130_fd_sc_hd__xor2_2 _26910_ (.A(_18407_),
    .B(_05334_),
    .X(_02373_));
 sky130_fd_sc_hd__nor2_2 _26911_ (.A(pcpi_rs1[19]),
    .B(_02374_),
    .Y(_05335_));
 sky130_fd_sc_hd__and2_2 _26912_ (.A(pcpi_rs1[19]),
    .B(_02374_),
    .X(_05336_));
 sky130_fd_sc_hd__nor2_2 _26913_ (.A(_05335_),
    .B(_05336_),
    .Y(_05337_));
 sky130_fd_sc_hd__and2_2 _26914_ (.A(pcpi_rs1[18]),
    .B(_02371_),
    .X(_05338_));
 sky130_fd_sc_hd__o21bai_2 _26915_ (.A1(_05329_),
    .A2(_05333_),
    .B1_N(_05338_),
    .Y(_05339_));
 sky130_fd_sc_hd__xor2_2 _26916_ (.A(_05337_),
    .B(_05339_),
    .X(_02601_));
 sky130_fd_sc_hd__nand3_2 _26917_ (.A(_05328_),
    .B(_02372_),
    .C(_02369_),
    .Y(_05340_));
 sky130_fd_sc_hd__xor2_2 _26918_ (.A(_02375_),
    .B(_05340_),
    .X(_02376_));
 sky130_fd_sc_hd__xnor2_2 _26919_ (.A(pcpi_rs1[20]),
    .B(_02377_),
    .Y(_05341_));
 sky130_fd_sc_hd__a21oi_2 _26920_ (.A1(_05339_),
    .A2(_05337_),
    .B1(_05336_),
    .Y(_05342_));
 sky130_fd_sc_hd__xor2_2 _26921_ (.A(_05341_),
    .B(_05342_),
    .X(_02603_));
 sky130_fd_sc_hd__nand3_2 _26922_ (.A(_05334_),
    .B(_02375_),
    .C(_02372_),
    .Y(_05343_));
 sky130_fd_sc_hd__xor2_2 _26923_ (.A(_02378_),
    .B(_05343_),
    .X(_02379_));
 sky130_fd_sc_hd__nor2_2 _26924_ (.A(pcpi_rs1[21]),
    .B(_02380_),
    .Y(_05344_));
 sky130_fd_sc_hd__and2_2 _26925_ (.A(pcpi_rs1[21]),
    .B(_02380_),
    .X(_05345_));
 sky130_fd_sc_hd__nor2_2 _26926_ (.A(_05344_),
    .B(_05345_),
    .Y(_05346_));
 sky130_fd_sc_hd__and2_2 _26927_ (.A(pcpi_rs1[20]),
    .B(_02377_),
    .X(_05347_));
 sky130_fd_sc_hd__o21bai_2 _26928_ (.A1(_05341_),
    .A2(_05342_),
    .B1_N(_05347_),
    .Y(_05348_));
 sky130_fd_sc_hd__xor2_2 _26929_ (.A(_05346_),
    .B(_05348_),
    .X(_02604_));
 sky130_fd_sc_hd__inv_2 _26930_ (.A(_18401_),
    .Y(_02381_));
 sky130_fd_sc_hd__nor2_2 _26931_ (.A(_18403_),
    .B(_05343_),
    .Y(_05349_));
 sky130_fd_sc_hd__xor2_2 _26932_ (.A(_18401_),
    .B(_05349_),
    .X(_02382_));
 sky130_fd_sc_hd__xnor2_2 _26933_ (.A(pcpi_rs1[22]),
    .B(_02383_),
    .Y(_05350_));
 sky130_fd_sc_hd__a21oi_2 _26934_ (.A1(_05348_),
    .A2(_05346_),
    .B1(_05345_),
    .Y(_05351_));
 sky130_fd_sc_hd__xor2_2 _26935_ (.A(_05350_),
    .B(_05351_),
    .X(_02605_));
 sky130_fd_sc_hd__inv_2 _26936_ (.A(_18398_),
    .Y(_02384_));
 sky130_fd_sc_hd__nor3_2 _26937_ (.A(_18400_),
    .B(_18402_),
    .C(_05343_),
    .Y(_05352_));
 sky130_fd_sc_hd__xor2_2 _26938_ (.A(_18399_),
    .B(_05352_),
    .X(_02385_));
 sky130_fd_sc_hd__nor2_2 _26939_ (.A(pcpi_rs1[23]),
    .B(_02386_),
    .Y(_05353_));
 sky130_fd_sc_hd__and2_2 _26940_ (.A(pcpi_rs1[23]),
    .B(_02386_),
    .X(_05354_));
 sky130_fd_sc_hd__nor2_2 _26941_ (.A(_05353_),
    .B(_05354_),
    .Y(_05355_));
 sky130_fd_sc_hd__and2_2 _26942_ (.A(pcpi_rs1[22]),
    .B(_02383_),
    .X(_05356_));
 sky130_fd_sc_hd__o21bai_2 _26943_ (.A1(_05350_),
    .A2(_05351_),
    .B1_N(_05356_),
    .Y(_05357_));
 sky130_fd_sc_hd__xor2_2 _26944_ (.A(_05355_),
    .B(_05357_),
    .X(_02606_));
 sky130_fd_sc_hd__nand3_2 _26945_ (.A(_05349_),
    .B(_02384_),
    .C(_02381_),
    .Y(_05358_));
 sky130_fd_sc_hd__xor2_2 _26946_ (.A(_02387_),
    .B(_05358_),
    .X(_02388_));
 sky130_fd_sc_hd__xor2_2 _26947_ (.A(_19703_),
    .B(_02389_),
    .X(_05359_));
 sky130_fd_sc_hd__a21oi_2 _26948_ (.A1(_05357_),
    .A2(_05355_),
    .B1(_05354_),
    .Y(_05360_));
 sky130_fd_sc_hd__xnor2_2 _26949_ (.A(_05359_),
    .B(_05360_),
    .Y(_02607_));
 sky130_fd_sc_hd__inv_2 _26950_ (.A(_18395_),
    .Y(_02390_));
 sky130_fd_sc_hd__nand3_2 _26951_ (.A(_05352_),
    .B(_02387_),
    .C(_02384_),
    .Y(_05361_));
 sky130_fd_sc_hd__xor2_2 _26952_ (.A(_02390_),
    .B(_05361_),
    .X(_02391_));
 sky130_fd_sc_hd__xor2_2 _26953_ (.A(_04251_),
    .B(_02392_),
    .X(_05362_));
 sky130_fd_sc_hd__and2b_2 _26954_ (.A_N(_05360_),
    .B(_05359_),
    .X(_05363_));
 sky130_fd_sc_hd__a21oi_2 _26955_ (.A1(_19055_),
    .A2(_02389_),
    .B1(_05363_),
    .Y(_05364_));
 sky130_fd_sc_hd__xnor2_2 _26956_ (.A(_05362_),
    .B(_05364_),
    .Y(_02608_));
 sky130_fd_sc_hd__inv_2 _26957_ (.A(_18392_),
    .Y(_02393_));
 sky130_fd_sc_hd__nor2_2 _26958_ (.A(_18394_),
    .B(_05361_),
    .Y(_05365_));
 sky130_fd_sc_hd__xor2_2 _26959_ (.A(_18393_),
    .B(_05365_),
    .X(_02394_));
 sky130_fd_sc_hd__xor2_2 _26960_ (.A(pcpi_rs1[26]),
    .B(_02395_),
    .X(_05366_));
 sky130_fd_sc_hd__nand2_2 _26961_ (.A(_05359_),
    .B(_05362_),
    .Y(_05367_));
 sky130_fd_sc_hd__o211a_2 _26962_ (.A1(_19052_),
    .A2(_02392_),
    .B1(_19703_),
    .C1(_02389_),
    .X(_05368_));
 sky130_fd_sc_hd__a21o_2 _26963_ (.A1(_19053_),
    .A2(_02392_),
    .B1(_05368_),
    .X(_05369_));
 sky130_fd_sc_hd__o21bai_2 _26964_ (.A1(_05367_),
    .A2(_05360_),
    .B1_N(_05369_),
    .Y(_05370_));
 sky130_fd_sc_hd__xor2_2 _26965_ (.A(_05366_),
    .B(_05370_),
    .X(_02609_));
 sky130_fd_sc_hd__nor3_2 _26966_ (.A(_18393_),
    .B(_18395_),
    .C(_05361_),
    .Y(_05371_));
 sky130_fd_sc_hd__xor2_2 _26967_ (.A(_18391_),
    .B(_05371_),
    .X(_02397_));
 sky130_fd_sc_hd__xnor2_2 _26968_ (.A(_04261_),
    .B(_02398_),
    .Y(_05372_));
 sky130_fd_sc_hd__and2_2 _26969_ (.A(_19051_),
    .B(_02395_),
    .X(_05373_));
 sky130_fd_sc_hd__a21oi_2 _26970_ (.A1(_05370_),
    .A2(_05366_),
    .B1(_05373_),
    .Y(_05374_));
 sky130_fd_sc_hd__xor2_2 _26971_ (.A(_05372_),
    .B(_05374_),
    .X(_02610_));
 sky130_fd_sc_hd__nand3_2 _26972_ (.A(_05365_),
    .B(_02396_),
    .C(_02393_),
    .Y(_05375_));
 sky130_fd_sc_hd__xor2_2 _26973_ (.A(_02399_),
    .B(_05375_),
    .X(_02400_));
 sky130_fd_sc_hd__xnor2_2 _26974_ (.A(_19046_),
    .B(_02401_),
    .Y(_05376_));
 sky130_fd_sc_hd__and2b_2 _26975_ (.A_N(_05372_),
    .B(_05366_),
    .X(_05377_));
 sky130_fd_sc_hd__o211a_2 _26976_ (.A1(_04261_),
    .A2(_02398_),
    .B1(_19050_),
    .C1(_02395_),
    .X(_05378_));
 sky130_fd_sc_hd__a21oi_2 _26977_ (.A1(_19047_),
    .A2(_02398_),
    .B1(_05378_),
    .Y(_05379_));
 sky130_fd_sc_hd__a21boi_2 _26978_ (.A1(_05370_),
    .A2(_05377_),
    .B1_N(_05379_),
    .Y(_05380_));
 sky130_fd_sc_hd__xor2_2 _26979_ (.A(_05376_),
    .B(_05380_),
    .X(_02611_));
 sky130_fd_sc_hd__inv_2 _26980_ (.A(_18386_),
    .Y(_02402_));
 sky130_fd_sc_hd__nor2_2 _26981_ (.A(_18388_),
    .B(_05375_),
    .Y(_05381_));
 sky130_fd_sc_hd__xor2_2 _26982_ (.A(_18387_),
    .B(_05381_),
    .X(_02403_));
 sky130_fd_sc_hd__nor2_2 _26983_ (.A(_19043_),
    .B(_02404_),
    .Y(_05382_));
 sky130_fd_sc_hd__and2_2 _26984_ (.A(_19043_),
    .B(_02404_),
    .X(_05383_));
 sky130_fd_sc_hd__nor2_2 _26985_ (.A(_05382_),
    .B(_05383_),
    .Y(_05384_));
 sky130_fd_sc_hd__nor2_2 _26986_ (.A(_19045_),
    .B(_02401_),
    .Y(_05385_));
 sky130_fd_sc_hd__and2_2 _26987_ (.A(pcpi_rs1[28]),
    .B(_02401_),
    .X(_05386_));
 sky130_fd_sc_hd__o21bai_2 _26988_ (.A1(_05385_),
    .A2(_05380_),
    .B1_N(_05386_),
    .Y(_05387_));
 sky130_fd_sc_hd__xor2_2 _26989_ (.A(_05384_),
    .B(_05387_),
    .X(_02612_));
 sky130_fd_sc_hd__nor3_2 _26990_ (.A(_18387_),
    .B(_18388_),
    .C(_05375_),
    .Y(_05388_));
 sky130_fd_sc_hd__xor2_2 _26991_ (.A(_18385_),
    .B(_05388_),
    .X(_02406_));
 sky130_fd_sc_hd__xnor2_2 _26992_ (.A(_04276_),
    .B(_02407_),
    .Y(_05389_));
 sky130_vsdinv _26993_ (.A(_05382_),
    .Y(_05390_));
 sky130_fd_sc_hd__a21oi_2 _26994_ (.A1(_05387_),
    .A2(_05390_),
    .B1(_05383_),
    .Y(_05391_));
 sky130_fd_sc_hd__xor2_2 _26995_ (.A(_05389_),
    .B(_05391_),
    .X(_02614_));
 sky130_fd_sc_hd__nand3_2 _26996_ (.A(_05381_),
    .B(_02405_),
    .C(_02402_),
    .Y(_05392_));
 sky130_fd_sc_hd__xor2_2 _26997_ (.A(_16978_),
    .B(_05392_),
    .X(_02408_));
 sky130_fd_sc_hd__nor2_2 _26998_ (.A(_19042_),
    .B(_02407_),
    .Y(_05393_));
 sky130_fd_sc_hd__and2_2 _26999_ (.A(_19041_),
    .B(_02407_),
    .X(_05394_));
 sky130_fd_sc_hd__o21bai_2 _27000_ (.A1(_05393_),
    .A2(_05391_),
    .B1_N(_05394_),
    .Y(_05395_));
 sky130_fd_sc_hd__xor2_2 _27001_ (.A(_16957_),
    .B(_02409_),
    .X(_05396_));
 sky130_fd_sc_hd__nand2_2 _27002_ (.A(_05395_),
    .B(_05396_),
    .Y(_05397_));
 sky130_vsdinv _27003_ (.A(_05394_),
    .Y(_05398_));
 sky130_vsdinv _27004_ (.A(_05396_),
    .Y(_05399_));
 sky130_fd_sc_hd__o211ai_2 _27005_ (.A1(_05393_),
    .A2(_05391_),
    .B1(_05398_),
    .C1(_05399_),
    .Y(_05400_));
 sky130_fd_sc_hd__nand2_2 _27006_ (.A(_05397_),
    .B(_05400_),
    .Y(_02615_));
 sky130_fd_sc_hd__buf_1 _27007_ (.A(\pcpi_mul.rs1[1] ),
    .X(_05401_));
 sky130_fd_sc_hd__buf_1 _27008_ (.A(_05401_),
    .X(_05402_));
 sky130_fd_sc_hd__buf_1 _27009_ (.A(_05402_),
    .X(_05403_));
 sky130_fd_sc_hd__buf_1 _27010_ (.A(_05403_),
    .X(_05404_));
 sky130_fd_sc_hd__nand2_2 _27011_ (.A(_05237_),
    .B(_05404_),
    .Y(_05405_));
 sky130_fd_sc_hd__nand2_2 _27012_ (.A(_18875_),
    .B(_05243_),
    .Y(_05406_));
 sky130_fd_sc_hd__xor2_2 _27013_ (.A(_05405_),
    .B(_05406_),
    .X(_02624_));
 sky130_fd_sc_hd__nor2_2 _27014_ (.A(_05405_),
    .B(_05406_),
    .Y(_05407_));
 sky130_fd_sc_hd__buf_1 _27015_ (.A(_18874_),
    .X(_05408_));
 sky130_fd_sc_hd__a22oi_2 _27016_ (.A1(_18868_),
    .A2(_05242_),
    .B1(_05408_),
    .B2(_05404_),
    .Y(_05409_));
 sky130_fd_sc_hd__and4_2 _27017_ (.A(_18868_),
    .B(_18874_),
    .C(_05404_),
    .D(_05241_),
    .X(_05410_));
 sky130_vsdinv _27018_ (.A(_05410_),
    .Y(_05411_));
 sky130_fd_sc_hd__buf_1 _27019_ (.A(_19292_),
    .X(_05412_));
 sky130_fd_sc_hd__buf_1 _27020_ (.A(_05412_),
    .X(_05413_));
 sky130_fd_sc_hd__buf_1 _27021_ (.A(_05413_),
    .X(_05414_));
 sky130_fd_sc_hd__and2_2 _27022_ (.A(_05237_),
    .B(_05414_),
    .X(_05415_));
 sky130_fd_sc_hd__nand3b_2 _27023_ (.A_N(_05409_),
    .B(_05411_),
    .C(_05415_),
    .Y(_05416_));
 sky130_fd_sc_hd__o21bai_2 _27024_ (.A1(_05409_),
    .A2(_05410_),
    .B1_N(_05415_),
    .Y(_05417_));
 sky130_fd_sc_hd__and2_2 _27025_ (.A(_05416_),
    .B(_05417_),
    .X(_05418_));
 sky130_fd_sc_hd__xor2_2 _27026_ (.A(_05407_),
    .B(_05418_),
    .X(_02625_));
 sky130_fd_sc_hd__nand3_2 _27027_ (.A(_05416_),
    .B(_05407_),
    .C(_05417_),
    .Y(_05419_));
 sky130_fd_sc_hd__buf_1 _27028_ (.A(\pcpi_mul.rs2[2] ),
    .X(_05420_));
 sky130_fd_sc_hd__buf_1 _27029_ (.A(_05420_),
    .X(_05421_));
 sky130_fd_sc_hd__buf_1 _27030_ (.A(_05421_),
    .X(_05422_));
 sky130_fd_sc_hd__buf_1 _27031_ (.A(\pcpi_mul.rs1[1] ),
    .X(_05423_));
 sky130_fd_sc_hd__buf_1 _27032_ (.A(_05423_),
    .X(_05424_));
 sky130_fd_sc_hd__buf_1 _27033_ (.A(_05424_),
    .X(_05425_));
 sky130_fd_sc_hd__nand2_2 _27034_ (.A(_05422_),
    .B(_05425_),
    .Y(_05426_));
 sky130_fd_sc_hd__buf_1 _27035_ (.A(\pcpi_mul.rs2[1] ),
    .X(_05427_));
 sky130_fd_sc_hd__buf_1 _27036_ (.A(_05427_),
    .X(_05428_));
 sky130_fd_sc_hd__buf_1 _27037_ (.A(_05428_),
    .X(_05429_));
 sky130_fd_sc_hd__buf_1 _27038_ (.A(\pcpi_mul.rs1[2] ),
    .X(_05430_));
 sky130_fd_sc_hd__buf_1 _27039_ (.A(_05430_),
    .X(_05431_));
 sky130_fd_sc_hd__buf_1 _27040_ (.A(_05431_),
    .X(_05432_));
 sky130_fd_sc_hd__nand2_2 _27041_ (.A(_05429_),
    .B(_05432_),
    .Y(_05433_));
 sky130_fd_sc_hd__xnor2_2 _27042_ (.A(_05426_),
    .B(_05433_),
    .Y(_05434_));
 sky130_fd_sc_hd__o21ai_2 _27043_ (.A1(_18858_),
    .A2(_19302_),
    .B1(_05434_),
    .Y(_05435_));
 sky130_vsdinv _27044_ (.A(_05434_),
    .Y(_05436_));
 sky130_fd_sc_hd__buf_1 _27045_ (.A(_18854_),
    .X(_05437_));
 sky130_fd_sc_hd__buf_1 _27046_ (.A(_05437_),
    .X(_05438_));
 sky130_fd_sc_hd__buf_1 _27047_ (.A(_05438_),
    .X(_05439_));
 sky130_fd_sc_hd__and2_2 _27048_ (.A(_05439_),
    .B(_05240_),
    .X(_05440_));
 sky130_fd_sc_hd__nand2_2 _27049_ (.A(_05436_),
    .B(_05440_),
    .Y(_05441_));
 sky130_fd_sc_hd__o2bb2ai_2 _27050_ (.A1_N(_05435_),
    .A2_N(_05441_),
    .B1(_18881_),
    .B2(_19290_),
    .Y(_05442_));
 sky130_fd_sc_hd__buf_1 _27051_ (.A(\pcpi_mul.rs1[3] ),
    .X(_05443_));
 sky130_fd_sc_hd__buf_1 _27052_ (.A(_05443_),
    .X(_05444_));
 sky130_fd_sc_hd__buf_1 _27053_ (.A(_05444_),
    .X(_05445_));
 sky130_fd_sc_hd__buf_1 _27054_ (.A(_05445_),
    .X(_05446_));
 sky130_fd_sc_hd__and2_2 _27055_ (.A(_05237_),
    .B(_05446_),
    .X(_05447_));
 sky130_fd_sc_hd__nand3_2 _27056_ (.A(_05441_),
    .B(_05435_),
    .C(_05447_),
    .Y(_05448_));
 sky130_fd_sc_hd__buf_1 _27057_ (.A(_05448_),
    .X(_05449_));
 sky130_fd_sc_hd__nand2_2 _27058_ (.A(_05442_),
    .B(_05449_),
    .Y(_05450_));
 sky130_fd_sc_hd__xnor2_2 _27059_ (.A(_05416_),
    .B(_05450_),
    .Y(_05451_));
 sky130_fd_sc_hd__and3_2 _27060_ (.A(_05442_),
    .B(_05410_),
    .C(_05449_),
    .X(_05452_));
 sky130_fd_sc_hd__a21oi_2 _27061_ (.A1(_05451_),
    .A2(_05411_),
    .B1(_05452_),
    .Y(_05453_));
 sky130_fd_sc_hd__xnor2_2 _27062_ (.A(_05419_),
    .B(_05453_),
    .Y(_02626_));
 sky130_fd_sc_hd__a21o_2 _27063_ (.A1(_05411_),
    .A2(_05416_),
    .B1(_05450_),
    .X(_05454_));
 sky130_fd_sc_hd__a22oi_2 _27064_ (.A1(_18867_),
    .A2(_05414_),
    .B1(_18873_),
    .B2(_05446_),
    .Y(_05455_));
 sky130_fd_sc_hd__and4_2 _27065_ (.A(_18867_),
    .B(_18873_),
    .C(_05446_),
    .D(_05414_),
    .X(_05456_));
 sky130_fd_sc_hd__nor2_2 _27066_ (.A(_05455_),
    .B(_05456_),
    .Y(_05457_));
 sky130_fd_sc_hd__buf_1 _27067_ (.A(\pcpi_mul.rs2[3] ),
    .X(_05458_));
 sky130_fd_sc_hd__buf_1 _27068_ (.A(_05458_),
    .X(_05459_));
 sky130_fd_sc_hd__buf_1 _27069_ (.A(_05459_),
    .X(_05460_));
 sky130_fd_sc_hd__and2_2 _27070_ (.A(_05460_),
    .B(_05403_),
    .X(_05461_));
 sky130_fd_sc_hd__nand2_2 _27071_ (.A(_05457_),
    .B(_05461_),
    .Y(_05462_));
 sky130_fd_sc_hd__buf_1 _27072_ (.A(_18849_),
    .X(_05463_));
 sky130_fd_sc_hd__buf_1 _27073_ (.A(_05463_),
    .X(_05464_));
 sky130_fd_sc_hd__buf_1 _27074_ (.A(_19300_),
    .X(_05465_));
 sky130_fd_sc_hd__buf_1 _27075_ (.A(_05465_),
    .X(_05466_));
 sky130_fd_sc_hd__nand2_2 _27076_ (.A(_05464_),
    .B(_05466_),
    .Y(_05467_));
 sky130_fd_sc_hd__buf_1 _27077_ (.A(\pcpi_mul.rs1[4] ),
    .X(_05468_));
 sky130_fd_sc_hd__buf_1 _27078_ (.A(_05468_),
    .X(_05469_));
 sky130_fd_sc_hd__buf_1 _27079_ (.A(_05469_),
    .X(_05470_));
 sky130_fd_sc_hd__buf_1 _27080_ (.A(_05470_),
    .X(_05471_));
 sky130_fd_sc_hd__nand2_2 _27081_ (.A(_05236_),
    .B(_05471_),
    .Y(_05472_));
 sky130_fd_sc_hd__xor2_2 _27082_ (.A(_05467_),
    .B(_05472_),
    .X(_05473_));
 sky130_fd_sc_hd__o21bai_2 _27083_ (.A1(_05455_),
    .A2(_05456_),
    .B1_N(_05461_),
    .Y(_05474_));
 sky130_fd_sc_hd__nand3_2 _27084_ (.A(_05462_),
    .B(_05473_),
    .C(_05474_),
    .Y(_05475_));
 sky130_fd_sc_hd__a21o_2 _27085_ (.A1(_05462_),
    .A2(_05474_),
    .B1(_05473_),
    .X(_05476_));
 sky130_fd_sc_hd__nand3b_2 _27086_ (.A_N(_05448_),
    .B(_05475_),
    .C(_05476_),
    .Y(_05477_));
 sky130_fd_sc_hd__nand2_2 _27087_ (.A(_05476_),
    .B(_05475_),
    .Y(_05478_));
 sky130_fd_sc_hd__nand2_2 _27088_ (.A(_05478_),
    .B(_05449_),
    .Y(_05479_));
 sky130_fd_sc_hd__nand3b_2 _27089_ (.A_N(_05426_),
    .B(_18874_),
    .C(_05414_),
    .Y(_05480_));
 sky130_fd_sc_hd__a21boi_2 _27090_ (.A1(_05436_),
    .A2(_05440_),
    .B1_N(_05480_),
    .Y(_05481_));
 sky130_vsdinv _27091_ (.A(_05481_),
    .Y(_05482_));
 sky130_fd_sc_hd__a21o_2 _27092_ (.A1(_05477_),
    .A2(_05479_),
    .B1(_05482_),
    .X(_05483_));
 sky130_fd_sc_hd__nand3_2 _27093_ (.A(_05477_),
    .B(_05479_),
    .C(_05482_),
    .Y(_05484_));
 sky130_fd_sc_hd__and3b_2 _27094_ (.A_N(_05454_),
    .B(_05483_),
    .C(_05484_),
    .X(_05485_));
 sky130_fd_sc_hd__buf_1 _27095_ (.A(_05485_),
    .X(_05486_));
 sky130_fd_sc_hd__a21boi_2 _27096_ (.A1(_05483_),
    .A2(_05484_),
    .B1_N(_05454_),
    .Y(_05487_));
 sky130_fd_sc_hd__nand3_2 _27097_ (.A(_05453_),
    .B(_05407_),
    .C(_05418_),
    .Y(_05488_));
 sky130_fd_sc_hd__o21a_2 _27098_ (.A1(_05486_),
    .A2(_05487_),
    .B1(_05488_),
    .X(_05489_));
 sky130_fd_sc_hd__nor3_2 _27099_ (.A(_05486_),
    .B(_05487_),
    .C(_05488_),
    .Y(_05490_));
 sky130_fd_sc_hd__nor2_2 _27100_ (.A(_05489_),
    .B(_05490_),
    .Y(_02627_));
 sky130_fd_sc_hd__buf_1 _27101_ (.A(\pcpi_mul.rs2[5] ),
    .X(_05491_));
 sky130_fd_sc_hd__buf_1 _27102_ (.A(_05491_),
    .X(_05492_));
 sky130_fd_sc_hd__buf_1 _27103_ (.A(_05423_),
    .X(_05493_));
 sky130_fd_sc_hd__buf_1 _27104_ (.A(_05412_),
    .X(_05494_));
 sky130_fd_sc_hd__a22oi_2 _27105_ (.A1(_05492_),
    .A2(_05493_),
    .B1(_18850_),
    .B2(_05494_),
    .Y(_05495_));
 sky130_fd_sc_hd__buf_1 _27106_ (.A(\pcpi_mul.rs2[5] ),
    .X(_05496_));
 sky130_fd_sc_hd__nand2_2 _27107_ (.A(_05496_),
    .B(_05401_),
    .Y(_05497_));
 sky130_fd_sc_hd__nand2_2 _27108_ (.A(_18849_),
    .B(_05412_),
    .Y(_05498_));
 sky130_fd_sc_hd__nor2_2 _27109_ (.A(_05497_),
    .B(_05498_),
    .Y(_05499_));
 sky130_fd_sc_hd__buf_1 _27110_ (.A(_19271_),
    .X(_05500_));
 sky130_fd_sc_hd__and2_2 _27111_ (.A(_05235_),
    .B(_05500_),
    .X(_05501_));
 sky130_fd_sc_hd__o21bai_2 _27112_ (.A1(_05495_),
    .A2(_05499_),
    .B1_N(_05501_),
    .Y(_05502_));
 sky130_fd_sc_hd__buf_1 _27113_ (.A(_18848_),
    .X(_05503_));
 sky130_fd_sc_hd__buf_1 _27114_ (.A(_05503_),
    .X(_05504_));
 sky130_fd_sc_hd__nand3b_2 _27115_ (.A_N(_05497_),
    .B(_05504_),
    .C(_05413_),
    .Y(_05505_));
 sky130_fd_sc_hd__nand2_2 _27116_ (.A(_05497_),
    .B(_05498_),
    .Y(_05506_));
 sky130_fd_sc_hd__nand3_2 _27117_ (.A(_05505_),
    .B(_05506_),
    .C(_05501_),
    .Y(_05507_));
 sky130_fd_sc_hd__nand2_2 _27118_ (.A(_05502_),
    .B(_05507_),
    .Y(_05508_));
 sky130_fd_sc_hd__buf_1 _27119_ (.A(_18848_),
    .X(_05509_));
 sky130_fd_sc_hd__buf_1 _27120_ (.A(_05423_),
    .X(_05510_));
 sky130_fd_sc_hd__nand2_2 _27121_ (.A(_05509_),
    .B(_05510_),
    .Y(_05511_));
 sky130_fd_sc_hd__buf_1 _27122_ (.A(\pcpi_mul.rs2[5] ),
    .X(_05512_));
 sky130_fd_sc_hd__buf_1 _27123_ (.A(_05512_),
    .X(_05513_));
 sky130_fd_sc_hd__nand2_2 _27124_ (.A(_05513_),
    .B(_19301_),
    .Y(_05514_));
 sky130_fd_sc_hd__nand2_2 _27125_ (.A(_05511_),
    .B(_05514_),
    .Y(_05515_));
 sky130_fd_sc_hd__buf_1 _27126_ (.A(\pcpi_mul.rs2[0] ),
    .X(_05516_));
 sky130_fd_sc_hd__buf_1 _27127_ (.A(\pcpi_mul.rs1[5] ),
    .X(_05517_));
 sky130_fd_sc_hd__buf_1 _27128_ (.A(_05517_),
    .X(_05518_));
 sky130_fd_sc_hd__and2_2 _27129_ (.A(_05516_),
    .B(_05518_),
    .X(_05519_));
 sky130_fd_sc_hd__nor2_2 _27130_ (.A(_05511_),
    .B(_05514_),
    .Y(_05520_));
 sky130_fd_sc_hd__a21o_2 _27131_ (.A1(_05515_),
    .A2(_05519_),
    .B1(_05520_),
    .X(_05521_));
 sky130_vsdinv _27132_ (.A(_05521_),
    .Y(_05522_));
 sky130_fd_sc_hd__nand2_2 _27133_ (.A(_05508_),
    .B(_05522_),
    .Y(_05523_));
 sky130_fd_sc_hd__nand3_2 _27134_ (.A(_05502_),
    .B(_05521_),
    .C(_05507_),
    .Y(_05524_));
 sky130_fd_sc_hd__buf_1 _27135_ (.A(_05524_),
    .X(_05525_));
 sky130_fd_sc_hd__buf_1 _27136_ (.A(_18871_),
    .X(_05526_));
 sky130_fd_sc_hd__buf_1 _27137_ (.A(\pcpi_mul.rs1[5] ),
    .X(_05527_));
 sky130_fd_sc_hd__buf_1 _27138_ (.A(_05527_),
    .X(_05528_));
 sky130_fd_sc_hd__buf_1 _27139_ (.A(_05528_),
    .X(_05529_));
 sky130_fd_sc_hd__a22oi_2 _27140_ (.A1(_05421_),
    .A2(_05470_),
    .B1(_05526_),
    .B2(_05529_),
    .Y(_05530_));
 sky130_fd_sc_hd__buf_1 _27141_ (.A(_05420_),
    .X(_05531_));
 sky130_fd_sc_hd__buf_1 _27142_ (.A(\pcpi_mul.rs1[4] ),
    .X(_05532_));
 sky130_fd_sc_hd__buf_1 _27143_ (.A(_05532_),
    .X(_05533_));
 sky130_fd_sc_hd__nand2_2 _27144_ (.A(_05531_),
    .B(_05533_),
    .Y(_05534_));
 sky130_fd_sc_hd__buf_1 _27145_ (.A(\pcpi_mul.rs2[1] ),
    .X(_05535_));
 sky130_fd_sc_hd__buf_1 _27146_ (.A(_05517_),
    .X(_05536_));
 sky130_fd_sc_hd__nand2_2 _27147_ (.A(_05535_),
    .B(_05536_),
    .Y(_05537_));
 sky130_fd_sc_hd__nor2_2 _27148_ (.A(_05534_),
    .B(_05537_),
    .Y(_05538_));
 sky130_vsdinv _27149_ (.A(_05538_),
    .Y(_05539_));
 sky130_fd_sc_hd__buf_1 _27150_ (.A(_19287_),
    .X(_05540_));
 sky130_fd_sc_hd__and2_2 _27151_ (.A(_05458_),
    .B(_05540_),
    .X(_05541_));
 sky130_fd_sc_hd__nand3b_2 _27152_ (.A_N(_05530_),
    .B(_05539_),
    .C(_05541_),
    .Y(_05542_));
 sky130_fd_sc_hd__o21bai_2 _27153_ (.A1(_05530_),
    .A2(_05538_),
    .B1_N(_05541_),
    .Y(_05543_));
 sky130_fd_sc_hd__nand2_2 _27154_ (.A(_05542_),
    .B(_05543_),
    .Y(_05544_));
 sky130_fd_sc_hd__buf_1 _27155_ (.A(_05544_),
    .X(_05545_));
 sky130_fd_sc_hd__a21boi_2 _27156_ (.A1(_05523_),
    .A2(_05525_),
    .B1_N(_05545_),
    .Y(_05546_));
 sky130_fd_sc_hd__a21oi_2 _27157_ (.A1(_05502_),
    .A2(_05507_),
    .B1(_05521_),
    .Y(_05547_));
 sky130_fd_sc_hd__nor3b_2 _27158_ (.A(_05545_),
    .B(_05547_),
    .C_N(_05525_),
    .Y(_05548_));
 sky130_fd_sc_hd__buf_1 _27159_ (.A(_05420_),
    .X(_05549_));
 sky130_fd_sc_hd__buf_1 _27160_ (.A(_05549_),
    .X(_05550_));
 sky130_fd_sc_hd__buf_1 _27161_ (.A(_19287_),
    .X(_05551_));
 sky130_fd_sc_hd__buf_1 _27162_ (.A(_05551_),
    .X(_05552_));
 sky130_fd_sc_hd__nand2_2 _27163_ (.A(_05550_),
    .B(_05552_),
    .Y(_05553_));
 sky130_fd_sc_hd__buf_1 _27164_ (.A(_05428_),
    .X(_05554_));
 sky130_fd_sc_hd__buf_1 _27165_ (.A(_05532_),
    .X(_05555_));
 sky130_fd_sc_hd__buf_1 _27166_ (.A(_05555_),
    .X(_05556_));
 sky130_fd_sc_hd__nand2_2 _27167_ (.A(_05554_),
    .B(_05556_),
    .Y(_05557_));
 sky130_fd_sc_hd__nor2_2 _27168_ (.A(_05553_),
    .B(_05557_),
    .Y(_05558_));
 sky130_fd_sc_hd__nand2_2 _27169_ (.A(_05553_),
    .B(_05557_),
    .Y(_05559_));
 sky130_vsdinv _27170_ (.A(_05559_),
    .Y(_05560_));
 sky130_fd_sc_hd__and2_2 _27171_ (.A(_05438_),
    .B(_05432_),
    .X(_05561_));
 sky130_fd_sc_hd__o21bai_2 _27172_ (.A1(_05558_),
    .A2(_05560_),
    .B1_N(_05561_),
    .Y(_05562_));
 sky130_fd_sc_hd__nand3b_2 _27173_ (.A_N(_05558_),
    .B(_05561_),
    .C(_05559_),
    .Y(_05563_));
 sky130_fd_sc_hd__nand2_2 _27174_ (.A(_05562_),
    .B(_05563_),
    .Y(_05564_));
 sky130_fd_sc_hd__nand3b_2 _27175_ (.A_N(_05520_),
    .B(_05519_),
    .C(_05515_),
    .Y(_05565_));
 sky130_fd_sc_hd__buf_1 _27176_ (.A(_18844_),
    .X(_05566_));
 sky130_fd_sc_hd__buf_1 _27177_ (.A(_05465_),
    .X(_05567_));
 sky130_fd_sc_hd__buf_1 _27178_ (.A(_05493_),
    .X(_05568_));
 sky130_fd_sc_hd__a22oi_2 _27179_ (.A1(_05566_),
    .A2(_05567_),
    .B1(_05464_),
    .B2(_05568_),
    .Y(_05569_));
 sky130_fd_sc_hd__o21bai_2 _27180_ (.A1(_05569_),
    .A2(_05520_),
    .B1_N(_05519_),
    .Y(_05570_));
 sky130_fd_sc_hd__nor2_2 _27181_ (.A(_05467_),
    .B(_05472_),
    .Y(_05571_));
 sky130_fd_sc_hd__a21oi_2 _27182_ (.A1(_05565_),
    .A2(_05570_),
    .B1(_05571_),
    .Y(_05572_));
 sky130_fd_sc_hd__nand3_2 _27183_ (.A(_05565_),
    .B(_05570_),
    .C(_05571_),
    .Y(_05573_));
 sky130_fd_sc_hd__o21ai_2 _27184_ (.A1(_05564_),
    .A2(_05572_),
    .B1(_05573_),
    .Y(_05574_));
 sky130_fd_sc_hd__o21bai_2 _27185_ (.A1(_05546_),
    .A2(_05548_),
    .B1_N(_05574_),
    .Y(_05575_));
 sky130_fd_sc_hd__nand2_2 _27186_ (.A(_05523_),
    .B(_05524_),
    .Y(_05576_));
 sky130_fd_sc_hd__nand2_2 _27187_ (.A(_05576_),
    .B(_05545_),
    .Y(_05577_));
 sky130_fd_sc_hd__nand3b_2 _27188_ (.A_N(_05544_),
    .B(_05523_),
    .C(_05525_),
    .Y(_05578_));
 sky130_fd_sc_hd__nand3_2 _27189_ (.A(_05577_),
    .B(_05574_),
    .C(_05578_),
    .Y(_05579_));
 sky130_fd_sc_hd__a21oi_2 _27190_ (.A1(_05559_),
    .A2(_05561_),
    .B1(_05558_),
    .Y(_05580_));
 sky130_vsdinv _27191_ (.A(_05580_),
    .Y(_05581_));
 sky130_fd_sc_hd__a21oi_2 _27192_ (.A1(_05575_),
    .A2(_05579_),
    .B1(_05581_),
    .Y(_05582_));
 sky130_fd_sc_hd__nand3_2 _27193_ (.A(_05575_),
    .B(_05581_),
    .C(_05579_),
    .Y(_05583_));
 sky130_vsdinv _27194_ (.A(_05583_),
    .Y(_05584_));
 sky130_fd_sc_hd__buf_1 _27195_ (.A(\pcpi_mul.rs2[6] ),
    .X(_05585_));
 sky130_fd_sc_hd__buf_1 _27196_ (.A(_05585_),
    .X(_05586_));
 sky130_fd_sc_hd__buf_1 _27197_ (.A(_05586_),
    .X(_05587_));
 sky130_fd_sc_hd__buf_1 _27198_ (.A(_05587_),
    .X(_05588_));
 sky130_fd_sc_hd__buf_1 _27199_ (.A(_05242_),
    .X(_05589_));
 sky130_fd_sc_hd__and2_2 _27200_ (.A(_05588_),
    .B(_05589_),
    .X(_05590_));
 sky130_fd_sc_hd__o21bai_2 _27201_ (.A1(_05582_),
    .A2(_05584_),
    .B1_N(_05590_),
    .Y(_05591_));
 sky130_fd_sc_hd__a21oi_2 _27202_ (.A1(_05577_),
    .A2(_05578_),
    .B1(_05574_),
    .Y(_05592_));
 sky130_vsdinv _27203_ (.A(_05579_),
    .Y(_05593_));
 sky130_fd_sc_hd__o21bai_2 _27204_ (.A1(_05592_),
    .A2(_05593_),
    .B1_N(_05581_),
    .Y(_05594_));
 sky130_fd_sc_hd__nand3_2 _27205_ (.A(_05594_),
    .B(_05590_),
    .C(_05583_),
    .Y(_05595_));
 sky130_fd_sc_hd__buf_1 _27206_ (.A(_05595_),
    .X(_05596_));
 sky130_fd_sc_hd__o2bb2ai_2 _27207_ (.A1_N(_05565_),
    .A2_N(_05570_),
    .B1(_05467_),
    .B2(_05472_),
    .Y(_05597_));
 sky130_vsdinv _27208_ (.A(_05564_),
    .Y(_05598_));
 sky130_fd_sc_hd__a21oi_2 _27209_ (.A1(_05597_),
    .A2(_05573_),
    .B1(_05598_),
    .Y(_05599_));
 sky130_fd_sc_hd__nand3_2 _27210_ (.A(_05598_),
    .B(_05597_),
    .C(_05573_),
    .Y(_05600_));
 sky130_vsdinv _27211_ (.A(_05600_),
    .Y(_05601_));
 sky130_vsdinv _27212_ (.A(_05475_),
    .Y(_05602_));
 sky130_fd_sc_hd__o21bai_2 _27213_ (.A1(_05599_),
    .A2(_05601_),
    .B1_N(_05602_),
    .Y(_05603_));
 sky130_fd_sc_hd__a21oi_2 _27214_ (.A1(_05457_),
    .A2(_05461_),
    .B1(_05456_),
    .Y(_05604_));
 sky130_vsdinv _27215_ (.A(_05604_),
    .Y(_05605_));
 sky130_fd_sc_hd__a21o_2 _27216_ (.A1(_05597_),
    .A2(_05573_),
    .B1(_05598_),
    .X(_05606_));
 sky130_fd_sc_hd__nand3_2 _27217_ (.A(_05606_),
    .B(_05602_),
    .C(_05600_),
    .Y(_05607_));
 sky130_fd_sc_hd__a21boi_2 _27218_ (.A1(_05603_),
    .A2(_05605_),
    .B1_N(_05607_),
    .Y(_05608_));
 sky130_vsdinv _27219_ (.A(_05608_),
    .Y(_05609_));
 sky130_fd_sc_hd__a21oi_2 _27220_ (.A1(_05591_),
    .A2(_05596_),
    .B1(_05609_),
    .Y(_05610_));
 sky130_fd_sc_hd__nand3_2 _27221_ (.A(_05591_),
    .B(_05595_),
    .C(_05609_),
    .Y(_05611_));
 sky130_vsdinv _27222_ (.A(_05611_),
    .Y(_05612_));
 sky130_fd_sc_hd__a21oi_2 _27223_ (.A1(_05603_),
    .A2(_05607_),
    .B1(_05605_),
    .Y(_05613_));
 sky130_vsdinv _27224_ (.A(_05462_),
    .Y(_05614_));
 sky130_fd_sc_hd__o211a_2 _27225_ (.A1(_05456_),
    .A2(_05614_),
    .B1(_05607_),
    .C1(_05603_),
    .X(_05615_));
 sky130_fd_sc_hd__nor2_2 _27226_ (.A(_05449_),
    .B(_05478_),
    .Y(_05616_));
 sky130_fd_sc_hd__a21oi_2 _27227_ (.A1(_05479_),
    .A2(_05482_),
    .B1(_05616_),
    .Y(_05617_));
 sky130_fd_sc_hd__o21ai_2 _27228_ (.A1(_05613_),
    .A2(_05615_),
    .B1(_05617_),
    .Y(_05618_));
 sky130_fd_sc_hd__nor3_2 _27229_ (.A(_05617_),
    .B(_05613_),
    .C(_05615_),
    .Y(_05619_));
 sky130_fd_sc_hd__a21oi_2 _27230_ (.A1(_05618_),
    .A2(_05485_),
    .B1(_05619_),
    .Y(_05620_));
 sky130_fd_sc_hd__o21bai_2 _27231_ (.A1(_05610_),
    .A2(_05612_),
    .B1_N(_05620_),
    .Y(_05621_));
 sky130_fd_sc_hd__a21oi_2 _27232_ (.A1(_05594_),
    .A2(_05583_),
    .B1(_05590_),
    .Y(_05622_));
 sky130_vsdinv _27233_ (.A(_05595_),
    .Y(_05623_));
 sky130_fd_sc_hd__o21bai_2 _27234_ (.A1(_05622_),
    .A2(_05623_),
    .B1_N(_05609_),
    .Y(_05624_));
 sky130_fd_sc_hd__buf_1 _27235_ (.A(_05611_),
    .X(_05625_));
 sky130_fd_sc_hd__nand3_2 _27236_ (.A(_05620_),
    .B(_05624_),
    .C(_05625_),
    .Y(_05626_));
 sky130_vsdinv _27237_ (.A(_05619_),
    .Y(_05627_));
 sky130_fd_sc_hd__nand3_2 _27238_ (.A(_05490_),
    .B(_05627_),
    .C(_05618_),
    .Y(_05628_));
 sky130_fd_sc_hd__a21oi_2 _27239_ (.A1(_05621_),
    .A2(_05626_),
    .B1(_05628_),
    .Y(_05629_));
 sky130_fd_sc_hd__and3_2 _27240_ (.A(_05621_),
    .B(_05628_),
    .C(_05626_),
    .X(_05630_));
 sky130_fd_sc_hd__nor2_2 _27241_ (.A(_05629_),
    .B(_05630_),
    .Y(_02683_));
 sky130_fd_sc_hd__nand3b_2 _27242_ (.A_N(_05619_),
    .B(_05486_),
    .C(_05618_),
    .Y(_05631_));
 sky130_fd_sc_hd__nor3_2 _27243_ (.A(_05610_),
    .B(_05612_),
    .C(_05631_),
    .Y(_05632_));
 sky130_fd_sc_hd__nor2_2 _27244_ (.A(_05632_),
    .B(_05629_),
    .Y(_05633_));
 sky130_fd_sc_hd__buf_1 _27245_ (.A(_18843_),
    .X(_05634_));
 sky130_fd_sc_hd__buf_1 _27246_ (.A(_19292_),
    .X(_05635_));
 sky130_fd_sc_hd__buf_1 _27247_ (.A(_05635_),
    .X(_05636_));
 sky130_fd_sc_hd__buf_1 _27248_ (.A(_18848_),
    .X(_05637_));
 sky130_fd_sc_hd__buf_1 _27249_ (.A(_05637_),
    .X(_05638_));
 sky130_fd_sc_hd__buf_1 _27250_ (.A(_05444_),
    .X(_05639_));
 sky130_fd_sc_hd__a22oi_2 _27251_ (.A1(_05634_),
    .A2(_05636_),
    .B1(_05638_),
    .B2(_05639_),
    .Y(_05640_));
 sky130_fd_sc_hd__nand2_2 _27252_ (.A(_05496_),
    .B(_19293_),
    .Y(_05641_));
 sky130_fd_sc_hd__buf_1 _27253_ (.A(\pcpi_mul.rs2[4] ),
    .X(_05642_));
 sky130_fd_sc_hd__buf_1 _27254_ (.A(_05642_),
    .X(_05643_));
 sky130_fd_sc_hd__buf_1 _27255_ (.A(_19287_),
    .X(_05644_));
 sky130_fd_sc_hd__nand2_2 _27256_ (.A(_05643_),
    .B(_05644_),
    .Y(_05645_));
 sky130_fd_sc_hd__nor2_2 _27257_ (.A(_05641_),
    .B(_05645_),
    .Y(_05646_));
 sky130_fd_sc_hd__buf_1 _27258_ (.A(\pcpi_mul.rs2[0] ),
    .X(_05647_));
 sky130_fd_sc_hd__buf_1 _27259_ (.A(\pcpi_mul.rs1[7] ),
    .X(_05648_));
 sky130_fd_sc_hd__buf_1 _27260_ (.A(_05648_),
    .X(_05649_));
 sky130_fd_sc_hd__and2_2 _27261_ (.A(_05647_),
    .B(_05649_),
    .X(_05650_));
 sky130_fd_sc_hd__o21bai_2 _27262_ (.A1(_05640_),
    .A2(_05646_),
    .B1_N(_05650_),
    .Y(_05651_));
 sky130_fd_sc_hd__buf_1 _27263_ (.A(_05503_),
    .X(_05652_));
 sky130_fd_sc_hd__nand3b_2 _27264_ (.A_N(_05641_),
    .B(_05652_),
    .C(_05445_),
    .Y(_05653_));
 sky130_fd_sc_hd__nand2_2 _27265_ (.A(_05641_),
    .B(_05645_),
    .Y(_05654_));
 sky130_fd_sc_hd__nand3_2 _27266_ (.A(_05653_),
    .B(_05654_),
    .C(_05650_),
    .Y(_05655_));
 sky130_fd_sc_hd__nand2_2 _27267_ (.A(_05651_),
    .B(_05655_),
    .Y(_05656_));
 sky130_fd_sc_hd__a21o_2 _27268_ (.A1(_05506_),
    .A2(_05501_),
    .B1(_05499_),
    .X(_05657_));
 sky130_vsdinv _27269_ (.A(_05657_),
    .Y(_05658_));
 sky130_fd_sc_hd__nand2_2 _27270_ (.A(_05656_),
    .B(_05658_),
    .Y(_05659_));
 sky130_fd_sc_hd__nand3_2 _27271_ (.A(_05651_),
    .B(_05657_),
    .C(_05655_),
    .Y(_05660_));
 sky130_fd_sc_hd__buf_1 _27272_ (.A(_05420_),
    .X(_05661_));
 sky130_fd_sc_hd__buf_1 _27273_ (.A(_05661_),
    .X(_05662_));
 sky130_fd_sc_hd__buf_1 _27274_ (.A(_05427_),
    .X(_05663_));
 sky130_fd_sc_hd__buf_1 _27275_ (.A(\pcpi_mul.rs1[6] ),
    .X(_05664_));
 sky130_fd_sc_hd__buf_1 _27276_ (.A(_05664_),
    .X(_05665_));
 sky130_fd_sc_hd__buf_1 _27277_ (.A(_05665_),
    .X(_05666_));
 sky130_fd_sc_hd__a22oi_2 _27278_ (.A1(_05662_),
    .A2(_05529_),
    .B1(_05663_),
    .B2(_05666_),
    .Y(_05667_));
 sky130_fd_sc_hd__buf_1 _27279_ (.A(\pcpi_mul.rs1[5] ),
    .X(_05668_));
 sky130_fd_sc_hd__buf_1 _27280_ (.A(_05668_),
    .X(_05669_));
 sky130_fd_sc_hd__nand2_2 _27281_ (.A(_05549_),
    .B(_05669_),
    .Y(_05670_));
 sky130_fd_sc_hd__buf_1 _27282_ (.A(_05665_),
    .X(_05671_));
 sky130_fd_sc_hd__nand2_2 _27283_ (.A(_05428_),
    .B(_05671_),
    .Y(_05672_));
 sky130_fd_sc_hd__nor2_2 _27284_ (.A(_05670_),
    .B(_05672_),
    .Y(_05673_));
 sky130_fd_sc_hd__buf_1 _27285_ (.A(_05468_),
    .X(_05674_));
 sky130_fd_sc_hd__and2_2 _27286_ (.A(_18854_),
    .B(_05674_),
    .X(_05675_));
 sky130_vsdinv _27287_ (.A(_05675_),
    .Y(_05676_));
 sky130_fd_sc_hd__nor3_2 _27288_ (.A(_05667_),
    .B(_05673_),
    .C(_05676_),
    .Y(_05677_));
 sky130_fd_sc_hd__o21a_2 _27289_ (.A1(_05667_),
    .A2(_05673_),
    .B1(_05676_),
    .X(_05678_));
 sky130_fd_sc_hd__nor2_2 _27290_ (.A(_05677_),
    .B(_05678_),
    .Y(_05679_));
 sky130_fd_sc_hd__a21oi_2 _27291_ (.A1(_05659_),
    .A2(_05660_),
    .B1(_05679_),
    .Y(_05680_));
 sky130_fd_sc_hd__nand3_2 _27292_ (.A(_05659_),
    .B(_05679_),
    .C(_05660_),
    .Y(_05681_));
 sky130_vsdinv _27293_ (.A(_05681_),
    .Y(_05682_));
 sky130_fd_sc_hd__o21ai_2 _27294_ (.A1(_05545_),
    .A2(_05547_),
    .B1(_05525_),
    .Y(_05683_));
 sky130_fd_sc_hd__o21bai_2 _27295_ (.A1(_05680_),
    .A2(_05682_),
    .B1_N(_05683_),
    .Y(_05684_));
 sky130_fd_sc_hd__buf_1 _27296_ (.A(_05684_),
    .X(_05685_));
 sky130_fd_sc_hd__o2bb2ai_2 _27297_ (.A1_N(_05660_),
    .A2_N(_05659_),
    .B1(_05678_),
    .B2(_05677_),
    .Y(_05686_));
 sky130_fd_sc_hd__nand3_2 _27298_ (.A(_05686_),
    .B(_05683_),
    .C(_05681_),
    .Y(_05687_));
 sky130_fd_sc_hd__buf_1 _27299_ (.A(_05687_),
    .X(_05688_));
 sky130_fd_sc_hd__nand2_2 _27300_ (.A(_05685_),
    .B(_05688_),
    .Y(_05689_));
 sky130_fd_sc_hd__buf_1 _27301_ (.A(_18858_),
    .X(_05690_));
 sky130_fd_sc_hd__o31a_2 _27302_ (.A1(_05690_),
    .A2(_19290_),
    .A3(_05530_),
    .B1(_05539_),
    .X(_05691_));
 sky130_fd_sc_hd__nand2_2 _27303_ (.A(_05689_),
    .B(_05691_),
    .Y(_05692_));
 sky130_vsdinv _27304_ (.A(_05691_),
    .Y(_05693_));
 sky130_fd_sc_hd__nand3_2 _27305_ (.A(_05685_),
    .B(_05693_),
    .C(_05688_),
    .Y(_05694_));
 sky130_fd_sc_hd__nand2_2 _27306_ (.A(_18835_),
    .B(_05240_),
    .Y(_05695_));
 sky130_fd_sc_hd__nand2_2 _27307_ (.A(_05588_),
    .B(_05404_),
    .Y(_05696_));
 sky130_fd_sc_hd__xor2_2 _27308_ (.A(_05695_),
    .B(_05696_),
    .X(_05697_));
 sky130_fd_sc_hd__a21oi_2 _27309_ (.A1(_05692_),
    .A2(_05694_),
    .B1(_05697_),
    .Y(_05698_));
 sky130_vsdinv _27310_ (.A(_05697_),
    .Y(_05699_));
 sky130_fd_sc_hd__a21oi_2 _27311_ (.A1(_05685_),
    .A2(_05688_),
    .B1(_05693_),
    .Y(_05700_));
 sky130_vsdinv _27312_ (.A(_05542_),
    .Y(_05701_));
 sky130_fd_sc_hd__o211a_2 _27313_ (.A1(_05538_),
    .A2(_05701_),
    .B1(_05687_),
    .C1(_05684_),
    .X(_05702_));
 sky130_fd_sc_hd__nor3_2 _27314_ (.A(_05699_),
    .B(_05700_),
    .C(_05702_),
    .Y(_05703_));
 sky130_fd_sc_hd__o21ai_2 _27315_ (.A1(_05698_),
    .A2(_05703_),
    .B1(_05596_),
    .Y(_05704_));
 sky130_fd_sc_hd__o21bai_2 _27316_ (.A1(_05700_),
    .A2(_05702_),
    .B1_N(_05697_),
    .Y(_05705_));
 sky130_fd_sc_hd__nand3_2 _27317_ (.A(_05692_),
    .B(_05697_),
    .C(_05694_),
    .Y(_05706_));
 sky130_fd_sc_hd__nand3b_2 _27318_ (.A_N(_05595_),
    .B(_05705_),
    .C(_05706_),
    .Y(_05707_));
 sky130_fd_sc_hd__buf_1 _27319_ (.A(_05707_),
    .X(_05708_));
 sky130_fd_sc_hd__a21boi_2 _27320_ (.A1(_05575_),
    .A2(_05581_),
    .B1_N(_05579_),
    .Y(_05709_));
 sky130_vsdinv _27321_ (.A(_05709_),
    .Y(_05710_));
 sky130_fd_sc_hd__a21oi_2 _27322_ (.A1(_05704_),
    .A2(_05708_),
    .B1(_05710_),
    .Y(_05711_));
 sky130_fd_sc_hd__a21boi_2 _27323_ (.A1(_05705_),
    .A2(_05706_),
    .B1_N(_05596_),
    .Y(_05712_));
 sky130_fd_sc_hd__buf_1 _27324_ (.A(_05703_),
    .X(_05713_));
 sky130_fd_sc_hd__nor3_2 _27325_ (.A(_05596_),
    .B(_05698_),
    .C(_05713_),
    .Y(_05714_));
 sky130_fd_sc_hd__nor3_2 _27326_ (.A(_05709_),
    .B(_05712_),
    .C(_05714_),
    .Y(_05715_));
 sky130_fd_sc_hd__a21oi_2 _27327_ (.A1(_05624_),
    .A2(_05619_),
    .B1(_05612_),
    .Y(_05716_));
 sky130_fd_sc_hd__o21bai_2 _27328_ (.A1(_05711_),
    .A2(_05715_),
    .B1_N(_05716_),
    .Y(_05717_));
 sky130_fd_sc_hd__o21bai_2 _27329_ (.A1(_05712_),
    .A2(_05714_),
    .B1_N(_05710_),
    .Y(_05718_));
 sky130_fd_sc_hd__nand3_2 _27330_ (.A(_05704_),
    .B(_05708_),
    .C(_05710_),
    .Y(_05719_));
 sky130_fd_sc_hd__nand3_2 _27331_ (.A(_05718_),
    .B(_05716_),
    .C(_05719_),
    .Y(_05720_));
 sky130_fd_sc_hd__and2_2 _27332_ (.A(_05717_),
    .B(_05720_),
    .X(_05721_));
 sky130_fd_sc_hd__xor2_2 _27333_ (.A(_05633_),
    .B(_05721_),
    .X(_02684_));
 sky130_fd_sc_hd__buf_1 _27334_ (.A(_05468_),
    .X(_05722_));
 sky130_fd_sc_hd__nand2_2 _27335_ (.A(_05503_),
    .B(_05722_),
    .Y(_05723_));
 sky130_fd_sc_hd__buf_1 _27336_ (.A(_05512_),
    .X(_05724_));
 sky130_fd_sc_hd__nand2_2 _27337_ (.A(_05724_),
    .B(_05551_),
    .Y(_05725_));
 sky130_fd_sc_hd__nor2_2 _27338_ (.A(_05723_),
    .B(_05725_),
    .Y(_05726_));
 sky130_fd_sc_hd__buf_1 _27339_ (.A(\pcpi_mul.rs1[8] ),
    .X(_05727_));
 sky130_fd_sc_hd__buf_1 _27340_ (.A(_05727_),
    .X(_05728_));
 sky130_fd_sc_hd__and2_2 _27341_ (.A(_05235_),
    .B(_05728_),
    .X(_05729_));
 sky130_fd_sc_hd__nand2_2 _27342_ (.A(_05723_),
    .B(_05725_),
    .Y(_05730_));
 sky130_fd_sc_hd__nand3b_2 _27343_ (.A_N(_05726_),
    .B(_05729_),
    .C(_05730_),
    .Y(_05731_));
 sky130_fd_sc_hd__buf_1 _27344_ (.A(_05503_),
    .X(_05732_));
 sky130_fd_sc_hd__buf_1 _27345_ (.A(_05722_),
    .X(_05733_));
 sky130_fd_sc_hd__a22oi_2 _27346_ (.A1(_05492_),
    .A2(_05445_),
    .B1(_05732_),
    .B2(_05733_),
    .Y(_05734_));
 sky130_fd_sc_hd__o21bai_2 _27347_ (.A1(_05734_),
    .A2(_05726_),
    .B1_N(_05729_),
    .Y(_05735_));
 sky130_fd_sc_hd__a21oi_2 _27348_ (.A1(_05654_),
    .A2(_05650_),
    .B1(_05646_),
    .Y(_05736_));
 sky130_fd_sc_hd__a21bo_2 _27349_ (.A1(_05731_),
    .A2(_05735_),
    .B1_N(_05736_),
    .X(_05737_));
 sky130_fd_sc_hd__nand3b_2 _27350_ (.A_N(_05736_),
    .B(_05731_),
    .C(_05735_),
    .Y(_05738_));
 sky130_fd_sc_hd__buf_1 _27351_ (.A(_05664_),
    .X(_05739_));
 sky130_fd_sc_hd__nand2_2 _27352_ (.A(_18865_),
    .B(_05739_),
    .Y(_05740_));
 sky130_fd_sc_hd__buf_1 _27353_ (.A(_05648_),
    .X(_05741_));
 sky130_fd_sc_hd__nand2_2 _27354_ (.A(_18871_),
    .B(_05741_),
    .Y(_05742_));
 sky130_fd_sc_hd__xor2_2 _27355_ (.A(_05740_),
    .B(_05742_),
    .X(_05743_));
 sky130_fd_sc_hd__buf_1 _27356_ (.A(_05458_),
    .X(_05744_));
 sky130_fd_sc_hd__buf_1 _27357_ (.A(_05527_),
    .X(_05745_));
 sky130_fd_sc_hd__buf_1 _27358_ (.A(_05745_),
    .X(_05746_));
 sky130_fd_sc_hd__and2_2 _27359_ (.A(_05744_),
    .B(_05746_),
    .X(_05747_));
 sky130_fd_sc_hd__nand2_2 _27360_ (.A(_05743_),
    .B(_05747_),
    .Y(_05748_));
 sky130_fd_sc_hd__xnor2_2 _27361_ (.A(_05740_),
    .B(_05742_),
    .Y(_05749_));
 sky130_fd_sc_hd__o21ai_2 _27362_ (.A1(_18856_),
    .A2(_19279_),
    .B1(_05749_),
    .Y(_05750_));
 sky130_fd_sc_hd__nand2_2 _27363_ (.A(_05748_),
    .B(_05750_),
    .Y(_05751_));
 sky130_fd_sc_hd__a21boi_2 _27364_ (.A1(_05737_),
    .A2(_05738_),
    .B1_N(_05751_),
    .Y(_05752_));
 sky130_fd_sc_hd__a21boi_2 _27365_ (.A1(_05731_),
    .A2(_05735_),
    .B1_N(_05736_),
    .Y(_05753_));
 sky130_fd_sc_hd__nor3b_2 _27366_ (.A(_05753_),
    .B(_05751_),
    .C_N(_05738_),
    .Y(_05754_));
 sky130_fd_sc_hd__a21boi_2 _27367_ (.A1(_05659_),
    .A2(_05679_),
    .B1_N(_05660_),
    .Y(_05755_));
 sky130_fd_sc_hd__o21ai_2 _27368_ (.A1(_05752_),
    .A2(_05754_),
    .B1(_05755_),
    .Y(_05756_));
 sky130_vsdinv _27369_ (.A(_05755_),
    .Y(_05757_));
 sky130_fd_sc_hd__nand3b_2 _27370_ (.A_N(_05751_),
    .B(_05738_),
    .C(_05737_),
    .Y(_05758_));
 sky130_fd_sc_hd__nand3b_2 _27371_ (.A_N(_05752_),
    .B(_05757_),
    .C(_05758_),
    .Y(_05759_));
 sky130_fd_sc_hd__buf_1 _27372_ (.A(_05759_),
    .X(_05760_));
 sky130_fd_sc_hd__o21ba_2 _27373_ (.A1(_05667_),
    .A2(_05676_),
    .B1_N(_05673_),
    .X(_05761_));
 sky130_fd_sc_hd__a21boi_2 _27374_ (.A1(_05756_),
    .A2(_05760_),
    .B1_N(_05761_),
    .Y(_05762_));
 sky130_fd_sc_hd__nand3b_2 _27375_ (.A_N(_05761_),
    .B(_05756_),
    .C(_05759_),
    .Y(_05763_));
 sky130_vsdinv _27376_ (.A(_05763_),
    .Y(_05764_));
 sky130_fd_sc_hd__nor2_2 _27377_ (.A(_05695_),
    .B(_05696_),
    .Y(_05765_));
 sky130_fd_sc_hd__buf_1 _27378_ (.A(\pcpi_mul.rs2[7] ),
    .X(_05766_));
 sky130_fd_sc_hd__buf_1 _27379_ (.A(_05766_),
    .X(_05767_));
 sky130_fd_sc_hd__buf_1 _27380_ (.A(_05767_),
    .X(_05768_));
 sky130_fd_sc_hd__buf_1 _27381_ (.A(_05768_),
    .X(_05769_));
 sky130_fd_sc_hd__nand2_2 _27382_ (.A(_05769_),
    .B(_05568_),
    .Y(_05770_));
 sky130_fd_sc_hd__buf_1 _27383_ (.A(\pcpi_mul.rs2[8] ),
    .X(_05771_));
 sky130_fd_sc_hd__buf_1 _27384_ (.A(_05771_),
    .X(_05772_));
 sky130_fd_sc_hd__buf_1 _27385_ (.A(_05772_),
    .X(_05773_));
 sky130_fd_sc_hd__nand2_2 _27386_ (.A(_05773_),
    .B(_05567_),
    .Y(_05774_));
 sky130_fd_sc_hd__nand2_2 _27387_ (.A(_05770_),
    .B(_05774_),
    .Y(_05775_));
 sky130_fd_sc_hd__nand3b_2 _27388_ (.A_N(_05770_),
    .B(_18830_),
    .C(_05241_),
    .Y(_05776_));
 sky130_fd_sc_hd__o2bb2ai_2 _27389_ (.A1_N(_05775_),
    .A2_N(_05776_),
    .B1(_18841_),
    .B2(_19295_),
    .Y(_05777_));
 sky130_fd_sc_hd__buf_1 _27390_ (.A(_05585_),
    .X(_05778_));
 sky130_fd_sc_hd__buf_1 _27391_ (.A(_05778_),
    .X(_05779_));
 sky130_fd_sc_hd__and2_2 _27392_ (.A(_05779_),
    .B(_05432_),
    .X(_05780_));
 sky130_fd_sc_hd__nand3_2 _27393_ (.A(_05776_),
    .B(_05775_),
    .C(_05780_),
    .Y(_05781_));
 sky130_fd_sc_hd__nand2_2 _27394_ (.A(_05777_),
    .B(_05781_),
    .Y(_05782_));
 sky130_fd_sc_hd__xnor2_2 _27395_ (.A(_05765_),
    .B(_05782_),
    .Y(_05783_));
 sky130_fd_sc_hd__o21bai_2 _27396_ (.A1(_05762_),
    .A2(_05764_),
    .B1_N(_05783_),
    .Y(_05784_));
 sky130_fd_sc_hd__buf_1 _27397_ (.A(_05784_),
    .X(_05785_));
 sky130_fd_sc_hd__a21bo_2 _27398_ (.A1(_05756_),
    .A2(_05760_),
    .B1_N(_05761_),
    .X(_05786_));
 sky130_fd_sc_hd__nand3_2 _27399_ (.A(_05786_),
    .B(_05783_),
    .C(_05763_),
    .Y(_05787_));
 sky130_fd_sc_hd__buf_1 _27400_ (.A(_05787_),
    .X(_05788_));
 sky130_fd_sc_hd__a21oi_2 _27401_ (.A1(_05785_),
    .A2(_05788_),
    .B1(_05713_),
    .Y(_05789_));
 sky130_fd_sc_hd__nand3_2 _27402_ (.A(_05784_),
    .B(_05703_),
    .C(_05787_),
    .Y(_05790_));
 sky130_vsdinv _27403_ (.A(_05790_),
    .Y(_05791_));
 sky130_fd_sc_hd__a21boi_2 _27404_ (.A1(_05685_),
    .A2(_05693_),
    .B1_N(_05688_),
    .Y(_05792_));
 sky130_fd_sc_hd__xnor2_2 _27405_ (.A(_05792_),
    .B(_05708_),
    .Y(_05793_));
 sky130_fd_sc_hd__o21ai_2 _27406_ (.A1(_05789_),
    .A2(_05791_),
    .B1(_05793_),
    .Y(_05794_));
 sky130_fd_sc_hd__nor2_2 _27407_ (.A(_05789_),
    .B(_05791_),
    .Y(_05795_));
 sky130_fd_sc_hd__nor2_2 _27408_ (.A(_05792_),
    .B(_05707_),
    .Y(_05796_));
 sky130_vsdinv _27409_ (.A(_05796_),
    .Y(_05797_));
 sky130_fd_sc_hd__nand2_2 _27410_ (.A(_05708_),
    .B(_05792_),
    .Y(_05798_));
 sky130_fd_sc_hd__nand3_2 _27411_ (.A(_05795_),
    .B(_05797_),
    .C(_05798_),
    .Y(_05799_));
 sky130_fd_sc_hd__nand2_2 _27412_ (.A(_05794_),
    .B(_05799_),
    .Y(_05800_));
 sky130_fd_sc_hd__o21ai_2 _27413_ (.A1(_05625_),
    .A2(_05711_),
    .B1(_05719_),
    .Y(_05801_));
 sky130_fd_sc_hd__nand2_2 _27414_ (.A(_05800_),
    .B(_05801_),
    .Y(_05802_));
 sky130_fd_sc_hd__o2111ai_2 _27415_ (.A1(_05625_),
    .A2(_05711_),
    .B1(_05719_),
    .C1(_05799_),
    .D1(_05794_),
    .Y(_05803_));
 sky130_fd_sc_hd__nand2_2 _27416_ (.A(_05802_),
    .B(_05803_),
    .Y(_05804_));
 sky130_fd_sc_hd__o2bb2ai_2 _27417_ (.A1_N(_05720_),
    .A2_N(_05717_),
    .B1(_05632_),
    .B2(_05629_),
    .Y(_05805_));
 sky130_fd_sc_hd__nor3_2 _27418_ (.A(_05627_),
    .B(_05610_),
    .C(_05612_),
    .Y(_05806_));
 sky130_fd_sc_hd__and3_2 _27419_ (.A(_05806_),
    .B(_05718_),
    .C(_05719_),
    .X(_05807_));
 sky130_vsdinv _27420_ (.A(_05807_),
    .Y(_05808_));
 sky130_fd_sc_hd__nand2_2 _27421_ (.A(_05805_),
    .B(_05808_),
    .Y(_05809_));
 sky130_fd_sc_hd__xor2_2 _27422_ (.A(_05804_),
    .B(_05809_),
    .X(_02685_));
 sky130_fd_sc_hd__nor3_2 _27423_ (.A(_05625_),
    .B(_05711_),
    .C(_05715_),
    .Y(_05810_));
 sky130_fd_sc_hd__and3_2 _27424_ (.A(_05810_),
    .B(_05799_),
    .C(_05794_),
    .X(_05811_));
 sky130_fd_sc_hd__a21oi_2 _27425_ (.A1(_05809_),
    .A2(_05804_),
    .B1(_05811_),
    .Y(_05812_));
 sky130_fd_sc_hd__buf_1 _27426_ (.A(_05512_),
    .X(_05813_));
 sky130_fd_sc_hd__buf_1 _27427_ (.A(_05532_),
    .X(_05814_));
 sky130_fd_sc_hd__nand2_2 _27428_ (.A(_05813_),
    .B(_05814_),
    .Y(_05815_));
 sky130_fd_sc_hd__buf_1 _27429_ (.A(_05642_),
    .X(_05816_));
 sky130_fd_sc_hd__nand2_2 _27430_ (.A(_05816_),
    .B(_05669_),
    .Y(_05817_));
 sky130_fd_sc_hd__nor2_2 _27431_ (.A(_05815_),
    .B(_05817_),
    .Y(_05818_));
 sky130_fd_sc_hd__nand2_2 _27432_ (.A(_05815_),
    .B(_05817_),
    .Y(_05819_));
 sky130_fd_sc_hd__buf_1 _27433_ (.A(_18877_),
    .X(_05820_));
 sky130_fd_sc_hd__buf_1 _27434_ (.A(_19256_),
    .X(_05821_));
 sky130_fd_sc_hd__buf_1 _27435_ (.A(_05821_),
    .X(_05822_));
 sky130_fd_sc_hd__and2_2 _27436_ (.A(_05820_),
    .B(_05822_),
    .X(_05823_));
 sky130_fd_sc_hd__nand3b_2 _27437_ (.A_N(_05818_),
    .B(_05819_),
    .C(_05823_),
    .Y(_05824_));
 sky130_fd_sc_hd__buf_1 _27438_ (.A(_05513_),
    .X(_05825_));
 sky130_fd_sc_hd__buf_1 _27439_ (.A(_05509_),
    .X(_05826_));
 sky130_fd_sc_hd__buf_1 _27440_ (.A(_05669_),
    .X(_05827_));
 sky130_fd_sc_hd__a22oi_2 _27441_ (.A1(_05825_),
    .A2(_05556_),
    .B1(_05826_),
    .B2(_05827_),
    .Y(_05828_));
 sky130_fd_sc_hd__o21bai_2 _27442_ (.A1(_05828_),
    .A2(_05818_),
    .B1_N(_05823_),
    .Y(_05829_));
 sky130_fd_sc_hd__nand2_2 _27443_ (.A(_05824_),
    .B(_05829_),
    .Y(_05830_));
 sky130_fd_sc_hd__a21oi_2 _27444_ (.A1(_05730_),
    .A2(_05729_),
    .B1(_05726_),
    .Y(_05831_));
 sky130_fd_sc_hd__nand2_2 _27445_ (.A(_05830_),
    .B(_05831_),
    .Y(_05832_));
 sky130_fd_sc_hd__nand3b_2 _27446_ (.A_N(_05831_),
    .B(_05829_),
    .C(_05824_),
    .Y(_05833_));
 sky130_fd_sc_hd__nand2_2 _27447_ (.A(_05832_),
    .B(_05833_),
    .Y(_05834_));
 sky130_fd_sc_hd__buf_1 _27448_ (.A(_05661_),
    .X(_05835_));
 sky130_fd_sc_hd__buf_1 _27449_ (.A(\pcpi_mul.rs1[7] ),
    .X(_05836_));
 sky130_fd_sc_hd__buf_1 _27450_ (.A(_05836_),
    .X(_05837_));
 sky130_fd_sc_hd__buf_1 _27451_ (.A(_05837_),
    .X(_05838_));
 sky130_fd_sc_hd__nand2_2 _27452_ (.A(_05835_),
    .B(_05838_),
    .Y(_05839_));
 sky130_fd_sc_hd__buf_1 _27453_ (.A(\pcpi_mul.rs1[8] ),
    .X(_05840_));
 sky130_fd_sc_hd__buf_1 _27454_ (.A(_05840_),
    .X(_05841_));
 sky130_fd_sc_hd__buf_1 _27455_ (.A(_05841_),
    .X(_05842_));
 sky130_fd_sc_hd__nand2_2 _27456_ (.A(_05554_),
    .B(_05842_),
    .Y(_05843_));
 sky130_fd_sc_hd__nand2_2 _27457_ (.A(_05839_),
    .B(_05843_),
    .Y(_05844_));
 sky130_fd_sc_hd__buf_1 _27458_ (.A(\pcpi_mul.rs1[8] ),
    .X(_05845_));
 sky130_fd_sc_hd__buf_1 _27459_ (.A(_05845_),
    .X(_05846_));
 sky130_fd_sc_hd__buf_1 _27460_ (.A(_05846_),
    .X(_05847_));
 sky130_fd_sc_hd__buf_1 _27461_ (.A(_05847_),
    .X(_05848_));
 sky130_fd_sc_hd__nand3b_2 _27462_ (.A_N(_05839_),
    .B(_18873_),
    .C(_05848_),
    .Y(_05849_));
 sky130_fd_sc_hd__o2bb2ai_2 _27463_ (.A1_N(_05844_),
    .A2_N(_05849_),
    .B1(_18857_),
    .B2(_19275_),
    .Y(_05850_));
 sky130_fd_sc_hd__buf_1 _27464_ (.A(_19271_),
    .X(_05851_));
 sky130_fd_sc_hd__buf_1 _27465_ (.A(_05851_),
    .X(_05852_));
 sky130_fd_sc_hd__and2_2 _27466_ (.A(_05438_),
    .B(_05852_),
    .X(_05853_));
 sky130_fd_sc_hd__nand3_2 _27467_ (.A(_05849_),
    .B(_05844_),
    .C(_05853_),
    .Y(_05854_));
 sky130_fd_sc_hd__nand2_2 _27468_ (.A(_05850_),
    .B(_05854_),
    .Y(_05855_));
 sky130_fd_sc_hd__nand2_2 _27469_ (.A(_05834_),
    .B(_05855_),
    .Y(_05856_));
 sky130_fd_sc_hd__nand3b_2 _27470_ (.A_N(_05855_),
    .B(_05832_),
    .C(_05833_),
    .Y(_05857_));
 sky130_fd_sc_hd__o21ai_2 _27471_ (.A1(_05753_),
    .A2(_05751_),
    .B1(_05738_),
    .Y(_05858_));
 sky130_fd_sc_hd__a21oi_2 _27472_ (.A1(_05856_),
    .A2(_05857_),
    .B1(_05858_),
    .Y(_05859_));
 sky130_fd_sc_hd__nand3_2 _27473_ (.A(_05858_),
    .B(_05856_),
    .C(_05857_),
    .Y(_05860_));
 sky130_vsdinv _27474_ (.A(_05860_),
    .Y(_05861_));
 sky130_fd_sc_hd__nor2_2 _27475_ (.A(_05740_),
    .B(_05742_),
    .Y(_05862_));
 sky130_fd_sc_hd__a21oi_2 _27476_ (.A1(_05743_),
    .A2(_05747_),
    .B1(_05862_),
    .Y(_05863_));
 sky130_vsdinv _27477_ (.A(_05863_),
    .Y(_05864_));
 sky130_fd_sc_hd__o21bai_2 _27478_ (.A1(_05859_),
    .A2(_05861_),
    .B1_N(_05864_),
    .Y(_05865_));
 sky130_fd_sc_hd__a21o_2 _27479_ (.A1(_05856_),
    .A2(_05857_),
    .B1(_05858_),
    .X(_05866_));
 sky130_fd_sc_hd__nand3_2 _27480_ (.A(_05866_),
    .B(_05864_),
    .C(_05860_),
    .Y(_05867_));
 sky130_fd_sc_hd__nand3_2 _27481_ (.A(_05777_),
    .B(_05765_),
    .C(_05781_),
    .Y(_05868_));
 sky130_fd_sc_hd__buf_1 _27482_ (.A(_18827_),
    .X(_05869_));
 sky130_fd_sc_hd__buf_1 _27483_ (.A(_05869_),
    .X(_05870_));
 sky130_fd_sc_hd__nand2_2 _27484_ (.A(_05870_),
    .B(_05493_),
    .Y(_05871_));
 sky130_fd_sc_hd__buf_1 _27485_ (.A(_05766_),
    .X(_05872_));
 sky130_fd_sc_hd__buf_1 _27486_ (.A(_05872_),
    .X(_05873_));
 sky130_fd_sc_hd__buf_1 _27487_ (.A(_19293_),
    .X(_05874_));
 sky130_fd_sc_hd__nand2_2 _27488_ (.A(_05873_),
    .B(_05874_),
    .Y(_05875_));
 sky130_fd_sc_hd__nand2_2 _27489_ (.A(_05871_),
    .B(_05875_),
    .Y(_05876_));
 sky130_fd_sc_hd__nor2_2 _27490_ (.A(_05871_),
    .B(_05875_),
    .Y(_05877_));
 sky130_vsdinv _27491_ (.A(_05877_),
    .Y(_05878_));
 sky130_fd_sc_hd__o2bb2ai_2 _27492_ (.A1_N(_05876_),
    .A2_N(_05878_),
    .B1(_18841_),
    .B2(_19289_),
    .Y(_05879_));
 sky130_fd_sc_hd__buf_1 _27493_ (.A(_05551_),
    .X(_05880_));
 sky130_fd_sc_hd__and2_2 _27494_ (.A(_05587_),
    .B(_05880_),
    .X(_05881_));
 sky130_fd_sc_hd__nand3b_2 _27495_ (.A_N(_05877_),
    .B(_05876_),
    .C(_05881_),
    .Y(_05882_));
 sky130_fd_sc_hd__nor2_2 _27496_ (.A(_05770_),
    .B(_05774_),
    .Y(_05883_));
 sky130_fd_sc_hd__a21oi_2 _27497_ (.A1(_05775_),
    .A2(_05780_),
    .B1(_05883_),
    .Y(_05884_));
 sky130_vsdinv _27498_ (.A(_05884_),
    .Y(_05885_));
 sky130_fd_sc_hd__a21oi_2 _27499_ (.A1(_05879_),
    .A2(_05882_),
    .B1(_05885_),
    .Y(_05886_));
 sky130_fd_sc_hd__nand3_2 _27500_ (.A(_05879_),
    .B(_05882_),
    .C(_05885_),
    .Y(_05887_));
 sky130_fd_sc_hd__or2b_2 _27501_ (.A(_05886_),
    .B_N(_05887_),
    .X(_05888_));
 sky130_fd_sc_hd__xor2_2 _27502_ (.A(_05868_),
    .B(_05888_),
    .X(_05889_));
 sky130_fd_sc_hd__a21oi_2 _27503_ (.A1(_05865_),
    .A2(_05867_),
    .B1(_05889_),
    .Y(_05890_));
 sky130_fd_sc_hd__nand3_2 _27504_ (.A(_05865_),
    .B(_05889_),
    .C(_05867_),
    .Y(_05891_));
 sky130_vsdinv _27505_ (.A(_05891_),
    .Y(_05892_));
 sky130_fd_sc_hd__o21ai_2 _27506_ (.A1(_05890_),
    .A2(_05892_),
    .B1(_05787_),
    .Y(_05893_));
 sky130_fd_sc_hd__buf_1 _27507_ (.A(\pcpi_mul.rs2[9] ),
    .X(_05894_));
 sky130_fd_sc_hd__buf_1 _27508_ (.A(_05894_),
    .X(_05895_));
 sky130_fd_sc_hd__buf_1 _27509_ (.A(_05895_),
    .X(_05896_));
 sky130_fd_sc_hd__and2_2 _27510_ (.A(_05896_),
    .B(_05243_),
    .X(_05897_));
 sky130_fd_sc_hd__a21o_2 _27511_ (.A1(_05865_),
    .A2(_05867_),
    .B1(_05889_),
    .X(_05898_));
 sky130_fd_sc_hd__nand3b_2 _27512_ (.A_N(_05787_),
    .B(_05898_),
    .C(_05891_),
    .Y(_05899_));
 sky130_fd_sc_hd__nand3_2 _27513_ (.A(_05893_),
    .B(_05897_),
    .C(_05899_),
    .Y(_05900_));
 sky130_fd_sc_hd__buf_1 _27514_ (.A(_05900_),
    .X(_05901_));
 sky130_fd_sc_hd__buf_1 _27515_ (.A(_05899_),
    .X(_05902_));
 sky130_fd_sc_hd__nand2_2 _27516_ (.A(_05893_),
    .B(_05902_),
    .Y(_05903_));
 sky130_vsdinv _27517_ (.A(_05897_),
    .Y(_05904_));
 sky130_fd_sc_hd__nand2_2 _27518_ (.A(_05903_),
    .B(_05904_),
    .Y(_05905_));
 sky130_vsdinv _27519_ (.A(_05760_),
    .Y(_05906_));
 sky130_fd_sc_hd__o2111ai_2 _27520_ (.A1(_05906_),
    .A2(_05764_),
    .B1(_05703_),
    .C1(_05788_),
    .D1(_05785_),
    .Y(_05907_));
 sky130_vsdinv _27521_ (.A(_05907_),
    .Y(_05908_));
 sky130_fd_sc_hd__a311oi_2 _27522_ (.A1(_05785_),
    .A2(_05713_),
    .A3(_05788_),
    .B1(_05906_),
    .C1(_05764_),
    .Y(_05909_));
 sky130_fd_sc_hd__o2bb2ai_2 _27523_ (.A1_N(_05901_),
    .A2_N(_05905_),
    .B1(_05908_),
    .B2(_05909_),
    .Y(_05910_));
 sky130_fd_sc_hd__nand3_2 _27524_ (.A(_05790_),
    .B(_05760_),
    .C(_05763_),
    .Y(_05911_));
 sky130_fd_sc_hd__and2_2 _27525_ (.A(_05911_),
    .B(_05907_),
    .X(_05912_));
 sky130_fd_sc_hd__nand3_2 _27526_ (.A(_05912_),
    .B(_05901_),
    .C(_05905_),
    .Y(_05913_));
 sky130_fd_sc_hd__nand2_2 _27527_ (.A(_05910_),
    .B(_05913_),
    .Y(_05914_));
 sky130_fd_sc_hd__a21o_2 _27528_ (.A1(_05785_),
    .A2(_05788_),
    .B1(_05713_),
    .X(_05915_));
 sky130_fd_sc_hd__a31oi_2 _27529_ (.A1(_05915_),
    .A2(_05798_),
    .A3(_05790_),
    .B1(_05796_),
    .Y(_05916_));
 sky130_fd_sc_hd__nand2_2 _27530_ (.A(_05914_),
    .B(_05916_),
    .Y(_05917_));
 sky130_vsdinv _27531_ (.A(_05916_),
    .Y(_05918_));
 sky130_fd_sc_hd__nand3_2 _27532_ (.A(_05910_),
    .B(_05913_),
    .C(_05918_),
    .Y(_05919_));
 sky130_fd_sc_hd__nand3_2 _27533_ (.A(_05794_),
    .B(_05799_),
    .C(_05715_),
    .Y(_05920_));
 sky130_fd_sc_hd__a21boi_2 _27534_ (.A1(_05917_),
    .A2(_05919_),
    .B1_N(_05920_),
    .Y(_05921_));
 sky130_fd_sc_hd__a21oi_2 _27535_ (.A1(_05910_),
    .A2(_05913_),
    .B1(_05918_),
    .Y(_05922_));
 sky130_fd_sc_hd__nor3b_2 _27536_ (.A(_05920_),
    .B(_05922_),
    .C_N(_05919_),
    .Y(_05923_));
 sky130_fd_sc_hd__nor2_2 _27537_ (.A(_05921_),
    .B(_05923_),
    .Y(_05924_));
 sky130_fd_sc_hd__xnor2_2 _27538_ (.A(_05812_),
    .B(_05924_),
    .Y(_02686_));
 sky130_fd_sc_hd__o21bai_2 _27539_ (.A1(_05921_),
    .A2(_05812_),
    .B1_N(_05923_),
    .Y(_05925_));
 sky130_fd_sc_hd__buf_1 _27540_ (.A(_18843_),
    .X(_05926_));
 sky130_fd_sc_hd__buf_1 _27541_ (.A(_05668_),
    .X(_05927_));
 sky130_fd_sc_hd__nand2_2 _27542_ (.A(_05926_),
    .B(_05927_),
    .Y(_05928_));
 sky130_fd_sc_hd__buf_1 _27543_ (.A(_05642_),
    .X(_05929_));
 sky130_fd_sc_hd__buf_1 _27544_ (.A(_05664_),
    .X(_05930_));
 sky130_fd_sc_hd__buf_1 _27545_ (.A(_05930_),
    .X(_05931_));
 sky130_fd_sc_hd__nand2_2 _27546_ (.A(_05929_),
    .B(_05931_),
    .Y(_05932_));
 sky130_fd_sc_hd__nor2_2 _27547_ (.A(_05928_),
    .B(_05932_),
    .Y(_05933_));
 sky130_fd_sc_hd__buf_1 _27548_ (.A(\pcpi_mul.rs1[10] ),
    .X(_05934_));
 sky130_fd_sc_hd__buf_1 _27549_ (.A(_05934_),
    .X(_05935_));
 sky130_fd_sc_hd__and2_2 _27550_ (.A(_05820_),
    .B(_05935_),
    .X(_05936_));
 sky130_fd_sc_hd__nand2_2 _27551_ (.A(_05928_),
    .B(_05932_),
    .Y(_05937_));
 sky130_fd_sc_hd__nand3b_2 _27552_ (.A_N(_05933_),
    .B(_05936_),
    .C(_05937_),
    .Y(_05938_));
 sky130_fd_sc_hd__buf_1 _27553_ (.A(_05637_),
    .X(_05939_));
 sky130_fd_sc_hd__buf_1 _27554_ (.A(_05939_),
    .X(_05940_));
 sky130_fd_sc_hd__buf_1 _27555_ (.A(_05666_),
    .X(_05941_));
 sky130_fd_sc_hd__a22oi_2 _27556_ (.A1(_05566_),
    .A2(_05827_),
    .B1(_05940_),
    .B2(_05941_),
    .Y(_05942_));
 sky130_fd_sc_hd__o21bai_2 _27557_ (.A1(_05942_),
    .A2(_05933_),
    .B1_N(_05936_),
    .Y(_05943_));
 sky130_fd_sc_hd__nand2_2 _27558_ (.A(_05938_),
    .B(_05943_),
    .Y(_05944_));
 sky130_fd_sc_hd__a21oi_2 _27559_ (.A1(_05819_),
    .A2(_05823_),
    .B1(_05818_),
    .Y(_05945_));
 sky130_fd_sc_hd__nand2_2 _27560_ (.A(_05944_),
    .B(_05945_),
    .Y(_05946_));
 sky130_fd_sc_hd__nand3b_2 _27561_ (.A_N(_05945_),
    .B(_05938_),
    .C(_05943_),
    .Y(_05947_));
 sky130_fd_sc_hd__nand2_2 _27562_ (.A(_05946_),
    .B(_05947_),
    .Y(_05948_));
 sky130_fd_sc_hd__buf_1 _27563_ (.A(_19256_),
    .X(_05949_));
 sky130_fd_sc_hd__buf_1 _27564_ (.A(_05949_),
    .X(_05950_));
 sky130_fd_sc_hd__buf_1 _27565_ (.A(_05950_),
    .X(_05951_));
 sky130_fd_sc_hd__a22oi_2 _27566_ (.A1(_05550_),
    .A2(_05842_),
    .B1(_05429_),
    .B2(_05951_),
    .Y(_05952_));
 sky130_fd_sc_hd__buf_1 _27567_ (.A(_05531_),
    .X(_05953_));
 sky130_fd_sc_hd__buf_1 _27568_ (.A(_05728_),
    .X(_05954_));
 sky130_fd_sc_hd__nand2_2 _27569_ (.A(_05953_),
    .B(_05954_),
    .Y(_05955_));
 sky130_fd_sc_hd__buf_1 _27570_ (.A(_05535_),
    .X(_05956_));
 sky130_fd_sc_hd__buf_1 _27571_ (.A(\pcpi_mul.rs1[9] ),
    .X(_05957_));
 sky130_fd_sc_hd__buf_1 _27572_ (.A(_05957_),
    .X(_05958_));
 sky130_fd_sc_hd__buf_1 _27573_ (.A(_05958_),
    .X(_05959_));
 sky130_fd_sc_hd__nand2_2 _27574_ (.A(_05956_),
    .B(_05959_),
    .Y(_05960_));
 sky130_fd_sc_hd__nor2_2 _27575_ (.A(_05955_),
    .B(_05960_),
    .Y(_05961_));
 sky130_vsdinv _27576_ (.A(_05961_),
    .Y(_05962_));
 sky130_fd_sc_hd__buf_1 _27577_ (.A(_05648_),
    .X(_05963_));
 sky130_fd_sc_hd__buf_1 _27578_ (.A(_05963_),
    .X(_05964_));
 sky130_fd_sc_hd__and2_2 _27579_ (.A(_05744_),
    .B(_05964_),
    .X(_05965_));
 sky130_fd_sc_hd__nand3b_2 _27580_ (.A_N(_05952_),
    .B(_05962_),
    .C(_05965_),
    .Y(_05966_));
 sky130_fd_sc_hd__o21bai_2 _27581_ (.A1(_05952_),
    .A2(_05961_),
    .B1_N(_05965_),
    .Y(_05967_));
 sky130_fd_sc_hd__nand2_2 _27582_ (.A(_05966_),
    .B(_05967_),
    .Y(_05968_));
 sky130_fd_sc_hd__nand2_2 _27583_ (.A(_05948_),
    .B(_05968_),
    .Y(_05969_));
 sky130_fd_sc_hd__nand3b_2 _27584_ (.A_N(_05968_),
    .B(_05946_),
    .C(_05947_),
    .Y(_05970_));
 sky130_fd_sc_hd__a21boi_2 _27585_ (.A1(_05824_),
    .A2(_05829_),
    .B1_N(_05831_),
    .Y(_05971_));
 sky130_fd_sc_hd__o21ai_2 _27586_ (.A1(_05855_),
    .A2(_05971_),
    .B1(_05833_),
    .Y(_05972_));
 sky130_fd_sc_hd__a21oi_2 _27587_ (.A1(_05969_),
    .A2(_05970_),
    .B1(_05972_),
    .Y(_05973_));
 sky130_fd_sc_hd__nand3_2 _27588_ (.A(_05969_),
    .B(_05972_),
    .C(_05970_),
    .Y(_05974_));
 sky130_vsdinv _27589_ (.A(_05974_),
    .Y(_05975_));
 sky130_fd_sc_hd__nor2_2 _27590_ (.A(_05839_),
    .B(_05843_),
    .Y(_05976_));
 sky130_fd_sc_hd__a21oi_2 _27591_ (.A1(_05844_),
    .A2(_05853_),
    .B1(_05976_),
    .Y(_05977_));
 sky130_vsdinv _27592_ (.A(_05977_),
    .Y(_05978_));
 sky130_fd_sc_hd__o21bai_2 _27593_ (.A1(_05973_),
    .A2(_05975_),
    .B1_N(_05978_),
    .Y(_05979_));
 sky130_fd_sc_hd__a21o_2 _27594_ (.A1(_05969_),
    .A2(_05970_),
    .B1(_05972_),
    .X(_05980_));
 sky130_fd_sc_hd__nand3_2 _27595_ (.A(_05980_),
    .B(_05978_),
    .C(_05974_),
    .Y(_05981_));
 sky130_fd_sc_hd__buf_1 _27596_ (.A(_05771_),
    .X(_05982_));
 sky130_fd_sc_hd__buf_1 _27597_ (.A(_05982_),
    .X(_05983_));
 sky130_fd_sc_hd__buf_1 _27598_ (.A(_05430_),
    .X(_05984_));
 sky130_fd_sc_hd__buf_1 _27599_ (.A(_05984_),
    .X(_05985_));
 sky130_fd_sc_hd__buf_1 _27600_ (.A(_05443_),
    .X(_05986_));
 sky130_fd_sc_hd__buf_1 _27601_ (.A(_05986_),
    .X(_05987_));
 sky130_fd_sc_hd__buf_1 _27602_ (.A(_05987_),
    .X(_05988_));
 sky130_fd_sc_hd__a22oi_2 _27603_ (.A1(_05983_),
    .A2(_05985_),
    .B1(_18834_),
    .B2(_05988_),
    .Y(_05989_));
 sky130_fd_sc_hd__buf_1 _27604_ (.A(_05869_),
    .X(_05990_));
 sky130_fd_sc_hd__nand2_2 _27605_ (.A(_05990_),
    .B(_05494_),
    .Y(_05991_));
 sky130_fd_sc_hd__buf_1 _27606_ (.A(_05766_),
    .X(_05992_));
 sky130_fd_sc_hd__buf_1 _27607_ (.A(_05992_),
    .X(_05993_));
 sky130_fd_sc_hd__nand2_2 _27608_ (.A(_05993_),
    .B(_05880_),
    .Y(_05994_));
 sky130_fd_sc_hd__nor2_2 _27609_ (.A(_05991_),
    .B(_05994_),
    .Y(_05995_));
 sky130_vsdinv _27610_ (.A(_05995_),
    .Y(_05996_));
 sky130_fd_sc_hd__buf_1 _27611_ (.A(_05722_),
    .X(_05997_));
 sky130_fd_sc_hd__and2_2 _27612_ (.A(_05587_),
    .B(_05997_),
    .X(_05998_));
 sky130_fd_sc_hd__nand3b_2 _27613_ (.A_N(_05989_),
    .B(_05996_),
    .C(_05998_),
    .Y(_05999_));
 sky130_fd_sc_hd__o21bai_2 _27614_ (.A1(_05989_),
    .A2(_05995_),
    .B1_N(_05998_),
    .Y(_06000_));
 sky130_fd_sc_hd__a21oi_2 _27615_ (.A1(_05876_),
    .A2(_05881_),
    .B1(_05877_),
    .Y(_06001_));
 sky130_vsdinv _27616_ (.A(_06001_),
    .Y(_06002_));
 sky130_fd_sc_hd__a21oi_2 _27617_ (.A1(_05999_),
    .A2(_06000_),
    .B1(_06002_),
    .Y(_06003_));
 sky130_fd_sc_hd__nand3_2 _27618_ (.A(_06002_),
    .B(_05999_),
    .C(_06000_),
    .Y(_06004_));
 sky130_fd_sc_hd__or2b_2 _27619_ (.A(_06003_),
    .B_N(_06004_),
    .X(_06005_));
 sky130_fd_sc_hd__o21ai_2 _27620_ (.A1(_05868_),
    .A2(_05886_),
    .B1(_05887_),
    .Y(_06006_));
 sky130_fd_sc_hd__xnor2_2 _27621_ (.A(_06005_),
    .B(_06006_),
    .Y(_06007_));
 sky130_fd_sc_hd__a21o_2 _27622_ (.A1(_05979_),
    .A2(_05981_),
    .B1(_06007_),
    .X(_06008_));
 sky130_fd_sc_hd__nand3_2 _27623_ (.A(_05979_),
    .B(_05981_),
    .C(_06007_),
    .Y(_06009_));
 sky130_fd_sc_hd__nand2_2 _27624_ (.A(_06008_),
    .B(_06009_),
    .Y(_06010_));
 sky130_fd_sc_hd__nand2_2 _27625_ (.A(_06010_),
    .B(_05891_),
    .Y(_06011_));
 sky130_fd_sc_hd__nand3_2 _27626_ (.A(_05892_),
    .B(_06008_),
    .C(_06009_),
    .Y(_06012_));
 sky130_fd_sc_hd__buf_1 _27627_ (.A(_06012_),
    .X(_06013_));
 sky130_fd_sc_hd__nand2_2 _27628_ (.A(_06011_),
    .B(_06013_),
    .Y(_06014_));
 sky130_fd_sc_hd__nand2_2 _27629_ (.A(_18820_),
    .B(_05567_),
    .Y(_06015_));
 sky130_fd_sc_hd__nand2_2 _27630_ (.A(_05896_),
    .B(_05568_),
    .Y(_06016_));
 sky130_fd_sc_hd__xor2_2 _27631_ (.A(_06015_),
    .B(_06016_),
    .X(_06017_));
 sky130_vsdinv _27632_ (.A(_06017_),
    .Y(_06018_));
 sky130_fd_sc_hd__nand2_2 _27633_ (.A(_06014_),
    .B(_06018_),
    .Y(_06019_));
 sky130_fd_sc_hd__nand3_2 _27634_ (.A(_06011_),
    .B(_06017_),
    .C(_06012_),
    .Y(_06020_));
 sky130_fd_sc_hd__buf_1 _27635_ (.A(_06020_),
    .X(_06021_));
 sky130_fd_sc_hd__a21boi_2 _27636_ (.A1(_06019_),
    .A2(_06021_),
    .B1_N(_05900_),
    .Y(_06022_));
 sky130_fd_sc_hd__a21oi_2 _27637_ (.A1(_06011_),
    .A2(_06013_),
    .B1(_06017_),
    .Y(_06023_));
 sky130_vsdinv _27638_ (.A(_06021_),
    .Y(_06024_));
 sky130_fd_sc_hd__nor3_2 _27639_ (.A(_05901_),
    .B(_06023_),
    .C(_06024_),
    .Y(_06025_));
 sky130_fd_sc_hd__a21oi_2 _27640_ (.A1(_05866_),
    .A2(_05864_),
    .B1(_05861_),
    .Y(_06026_));
 sky130_fd_sc_hd__xnor2_2 _27641_ (.A(_06026_),
    .B(_05902_),
    .Y(_06027_));
 sky130_vsdinv _27642_ (.A(_06027_),
    .Y(_06028_));
 sky130_fd_sc_hd__o21bai_2 _27643_ (.A1(_06022_),
    .A2(_06025_),
    .B1_N(_06028_),
    .Y(_06029_));
 sky130_fd_sc_hd__o22ai_2 _27644_ (.A1(_05904_),
    .A2(_05903_),
    .B1(_06023_),
    .B2(_06024_),
    .Y(_06030_));
 sky130_fd_sc_hd__nand3b_2 _27645_ (.A_N(_05900_),
    .B(_06019_),
    .C(_06021_),
    .Y(_06031_));
 sky130_fd_sc_hd__nand3_2 _27646_ (.A(_06030_),
    .B(_06028_),
    .C(_06031_),
    .Y(_06032_));
 sky130_fd_sc_hd__a31o_2 _27647_ (.A1(_05905_),
    .A2(_05901_),
    .A3(_05911_),
    .B1(_05908_),
    .X(_06033_));
 sky130_fd_sc_hd__a21oi_2 _27648_ (.A1(_06029_),
    .A2(_06032_),
    .B1(_06033_),
    .Y(_06034_));
 sky130_fd_sc_hd__and3_2 _27649_ (.A(_06029_),
    .B(_06033_),
    .C(_06032_),
    .X(_06035_));
 sky130_fd_sc_hd__nor3_2 _27650_ (.A(_05919_),
    .B(_06034_),
    .C(_06035_),
    .Y(_06036_));
 sky130_fd_sc_hd__o22ai_2 _27651_ (.A1(_05914_),
    .A2(_05916_),
    .B1(_06034_),
    .B2(_06035_),
    .Y(_06037_));
 sky130_fd_sc_hd__and2b_2 _27652_ (.A_N(_06036_),
    .B(_06037_),
    .X(_06038_));
 sky130_fd_sc_hd__xor2_2 _27653_ (.A(_05925_),
    .B(_06038_),
    .X(_02629_));
 sky130_fd_sc_hd__a21oi_2 _27654_ (.A1(_05925_),
    .A2(_06037_),
    .B1(_06036_),
    .Y(_06039_));
 sky130_fd_sc_hd__buf_1 _27655_ (.A(_05512_),
    .X(_06040_));
 sky130_fd_sc_hd__buf_1 _27656_ (.A(_05930_),
    .X(_06041_));
 sky130_fd_sc_hd__nand2_2 _27657_ (.A(_06040_),
    .B(_06041_),
    .Y(_06042_));
 sky130_fd_sc_hd__buf_1 _27658_ (.A(_19267_),
    .X(_06043_));
 sky130_fd_sc_hd__nand2_2 _27659_ (.A(_05643_),
    .B(_06043_),
    .Y(_06044_));
 sky130_fd_sc_hd__nor2_2 _27660_ (.A(_06042_),
    .B(_06044_),
    .Y(_06045_));
 sky130_fd_sc_hd__buf_1 _27661_ (.A(\pcpi_mul.rs1[11] ),
    .X(_06046_));
 sky130_fd_sc_hd__buf_1 _27662_ (.A(_06046_),
    .X(_06047_));
 sky130_fd_sc_hd__and2_2 _27663_ (.A(_18878_),
    .B(_06047_),
    .X(_06048_));
 sky130_fd_sc_hd__nand2_2 _27664_ (.A(_06042_),
    .B(_06044_),
    .Y(_06049_));
 sky130_fd_sc_hd__nand3b_2 _27665_ (.A_N(_06045_),
    .B(_06048_),
    .C(_06049_),
    .Y(_06050_));
 sky130_fd_sc_hd__buf_1 _27666_ (.A(_05724_),
    .X(_06051_));
 sky130_fd_sc_hd__buf_1 _27667_ (.A(_05500_),
    .X(_06052_));
 sky130_fd_sc_hd__a22oi_2 _27668_ (.A1(_06051_),
    .A2(_06052_),
    .B1(_05463_),
    .B2(_05964_),
    .Y(_06053_));
 sky130_fd_sc_hd__o21bai_2 _27669_ (.A1(_06053_),
    .A2(_06045_),
    .B1_N(_06048_),
    .Y(_06054_));
 sky130_fd_sc_hd__nand2_2 _27670_ (.A(_06050_),
    .B(_06054_),
    .Y(_06055_));
 sky130_fd_sc_hd__a21oi_2 _27671_ (.A1(_05937_),
    .A2(_05936_),
    .B1(_05933_),
    .Y(_06056_));
 sky130_fd_sc_hd__nand2_2 _27672_ (.A(_06055_),
    .B(_06056_),
    .Y(_06057_));
 sky130_fd_sc_hd__nand3b_2 _27673_ (.A_N(_06056_),
    .B(_06050_),
    .C(_06054_),
    .Y(_06058_));
 sky130_fd_sc_hd__nand2_2 _27674_ (.A(_06057_),
    .B(_06058_),
    .Y(_06059_));
 sky130_fd_sc_hd__buf_1 _27675_ (.A(_05957_),
    .X(_06060_));
 sky130_fd_sc_hd__buf_1 _27676_ (.A(_06060_),
    .X(_06061_));
 sky130_fd_sc_hd__buf_1 _27677_ (.A(\pcpi_mul.rs1[10] ),
    .X(_06062_));
 sky130_fd_sc_hd__buf_1 _27678_ (.A(_06062_),
    .X(_06063_));
 sky130_fd_sc_hd__buf_1 _27679_ (.A(_06063_),
    .X(_06064_));
 sky130_fd_sc_hd__a22oi_2 _27680_ (.A1(_05835_),
    .A2(_06061_),
    .B1(_05956_),
    .B2(_06064_),
    .Y(_06065_));
 sky130_fd_sc_hd__nand2_2 _27681_ (.A(_18866_),
    .B(_05822_),
    .Y(_06066_));
 sky130_fd_sc_hd__buf_1 _27682_ (.A(\pcpi_mul.rs1[10] ),
    .X(_06067_));
 sky130_fd_sc_hd__buf_1 _27683_ (.A(_06067_),
    .X(_06068_));
 sky130_fd_sc_hd__buf_1 _27684_ (.A(_06068_),
    .X(_06069_));
 sky130_fd_sc_hd__nand2_2 _27685_ (.A(_05526_),
    .B(_06069_),
    .Y(_06070_));
 sky130_fd_sc_hd__nor2_2 _27686_ (.A(_06066_),
    .B(_06070_),
    .Y(_06071_));
 sky130_vsdinv _27687_ (.A(_06071_),
    .Y(_06072_));
 sky130_fd_sc_hd__buf_1 _27688_ (.A(_18854_),
    .X(_06073_));
 sky130_fd_sc_hd__buf_1 _27689_ (.A(_05845_),
    .X(_06074_));
 sky130_fd_sc_hd__buf_1 _27690_ (.A(_06074_),
    .X(_06075_));
 sky130_fd_sc_hd__and2_2 _27691_ (.A(_06073_),
    .B(_06075_),
    .X(_06076_));
 sky130_fd_sc_hd__nand3b_2 _27692_ (.A_N(_06065_),
    .B(_06072_),
    .C(_06076_),
    .Y(_06077_));
 sky130_fd_sc_hd__o21bai_2 _27693_ (.A1(_06065_),
    .A2(_06071_),
    .B1_N(_06076_),
    .Y(_06078_));
 sky130_fd_sc_hd__nand2_2 _27694_ (.A(_06077_),
    .B(_06078_),
    .Y(_06079_));
 sky130_fd_sc_hd__nand2_2 _27695_ (.A(_06059_),
    .B(_06079_),
    .Y(_06080_));
 sky130_fd_sc_hd__nand3b_2 _27696_ (.A_N(_06079_),
    .B(_06057_),
    .C(_06058_),
    .Y(_06081_));
 sky130_fd_sc_hd__nand2_2 _27697_ (.A(_06080_),
    .B(_06081_),
    .Y(_06082_));
 sky130_fd_sc_hd__a21boi_2 _27698_ (.A1(_05938_),
    .A2(_05943_),
    .B1_N(_05945_),
    .Y(_06083_));
 sky130_fd_sc_hd__o21ai_2 _27699_ (.A1(_05968_),
    .A2(_06083_),
    .B1(_05947_),
    .Y(_06084_));
 sky130_vsdinv _27700_ (.A(_06084_),
    .Y(_06085_));
 sky130_fd_sc_hd__nand2_2 _27701_ (.A(_06082_),
    .B(_06085_),
    .Y(_06086_));
 sky130_fd_sc_hd__nand3_2 _27702_ (.A(_06080_),
    .B(_06084_),
    .C(_06081_),
    .Y(_06087_));
 sky130_fd_sc_hd__o31a_2 _27703_ (.A1(_05690_),
    .A2(_19269_),
    .A3(_05952_),
    .B1(_05962_),
    .X(_06088_));
 sky130_vsdinv _27704_ (.A(_06088_),
    .Y(_06089_));
 sky130_fd_sc_hd__a21oi_2 _27705_ (.A1(_06086_),
    .A2(_06087_),
    .B1(_06089_),
    .Y(_06090_));
 sky130_fd_sc_hd__nand3_2 _27706_ (.A(_06086_),
    .B(_06089_),
    .C(_06087_),
    .Y(_06091_));
 sky130_vsdinv _27707_ (.A(_06091_),
    .Y(_06092_));
 sky130_vsdinv _27708_ (.A(_06004_),
    .Y(_06093_));
 sky130_fd_sc_hd__nor3_2 _27709_ (.A(_05887_),
    .B(_06003_),
    .C(_06093_),
    .Y(_06094_));
 sky130_fd_sc_hd__buf_1 _27710_ (.A(\pcpi_mul.rs2[7] ),
    .X(_06095_));
 sky130_fd_sc_hd__buf_1 _27711_ (.A(_06095_),
    .X(_06096_));
 sky130_fd_sc_hd__buf_1 _27712_ (.A(_06096_),
    .X(_06097_));
 sky130_fd_sc_hd__a22oi_2 _27713_ (.A1(_05990_),
    .A2(_05880_),
    .B1(_06097_),
    .B2(_05997_),
    .Y(_06098_));
 sky130_fd_sc_hd__and4_2 _27714_ (.A(_05990_),
    .B(_05993_),
    .C(_05997_),
    .D(_05552_),
    .X(_06099_));
 sky130_fd_sc_hd__buf_1 _27715_ (.A(\pcpi_mul.rs2[6] ),
    .X(_06100_));
 sky130_fd_sc_hd__buf_1 _27716_ (.A(_06100_),
    .X(_06101_));
 sky130_fd_sc_hd__buf_1 _27717_ (.A(_05528_),
    .X(_06102_));
 sky130_fd_sc_hd__and2_2 _27718_ (.A(_06101_),
    .B(_06102_),
    .X(_06103_));
 sky130_fd_sc_hd__o21bai_2 _27719_ (.A1(_06098_),
    .A2(_06099_),
    .B1_N(_06103_),
    .Y(_06104_));
 sky130_fd_sc_hd__buf_1 _27720_ (.A(_18828_),
    .X(_06105_));
 sky130_fd_sc_hd__nand2_2 _27721_ (.A(_06105_),
    .B(_05639_),
    .Y(_06106_));
 sky130_fd_sc_hd__nand3b_2 _27722_ (.A_N(_06106_),
    .B(_05769_),
    .C(_05471_),
    .Y(_06107_));
 sky130_fd_sc_hd__nand3b_2 _27723_ (.A_N(_06098_),
    .B(_06107_),
    .C(_06103_),
    .Y(_06108_));
 sky130_fd_sc_hd__nor2_2 _27724_ (.A(_06015_),
    .B(_06016_),
    .Y(_06109_));
 sky130_fd_sc_hd__a21oi_2 _27725_ (.A1(_06104_),
    .A2(_06108_),
    .B1(_06109_),
    .Y(_06110_));
 sky130_fd_sc_hd__nand3_2 _27726_ (.A(_06104_),
    .B(_06108_),
    .C(_06109_),
    .Y(_06111_));
 sky130_vsdinv _27727_ (.A(_06111_),
    .Y(_06112_));
 sky130_fd_sc_hd__buf_1 _27728_ (.A(_18839_),
    .X(_06113_));
 sky130_fd_sc_hd__buf_1 _27729_ (.A(_06113_),
    .X(_06114_));
 sky130_fd_sc_hd__o31a_2 _27730_ (.A1(_06114_),
    .A2(_19282_),
    .A3(_05989_),
    .B1(_05996_),
    .X(_06115_));
 sky130_vsdinv _27731_ (.A(_06115_),
    .Y(_06116_));
 sky130_fd_sc_hd__o21bai_2 _27732_ (.A1(_06110_),
    .A2(_06112_),
    .B1_N(_06116_),
    .Y(_06117_));
 sky130_fd_sc_hd__nand3b_2 _27733_ (.A_N(_06110_),
    .B(_06116_),
    .C(_06111_),
    .Y(_06118_));
 sky130_fd_sc_hd__nand2_2 _27734_ (.A(_06117_),
    .B(_06118_),
    .Y(_06119_));
 sky130_fd_sc_hd__o21ai_2 _27735_ (.A1(_06093_),
    .A2(_06094_),
    .B1(_06119_),
    .Y(_06120_));
 sky130_fd_sc_hd__o2111ai_2 _27736_ (.A1(_05887_),
    .A2(_06003_),
    .B1(_06004_),
    .C1(_06118_),
    .D1(_06117_),
    .Y(_06121_));
 sky130_fd_sc_hd__nand2_2 _27737_ (.A(_06120_),
    .B(_06121_),
    .Y(_06122_));
 sky130_fd_sc_hd__o21bai_2 _27738_ (.A1(_06090_),
    .A2(_06092_),
    .B1_N(_06122_),
    .Y(_06123_));
 sky130_fd_sc_hd__nand2_2 _27739_ (.A(_06086_),
    .B(_06087_),
    .Y(_06124_));
 sky130_fd_sc_hd__nand2_2 _27740_ (.A(_06124_),
    .B(_06088_),
    .Y(_06125_));
 sky130_fd_sc_hd__nand3_2 _27741_ (.A(_06125_),
    .B(_06091_),
    .C(_06122_),
    .Y(_06126_));
 sky130_fd_sc_hd__nand2_2 _27742_ (.A(_06123_),
    .B(_06126_),
    .Y(_06127_));
 sky130_fd_sc_hd__nor3_2 _27743_ (.A(_05868_),
    .B(_06005_),
    .C(_05888_),
    .Y(_06128_));
 sky130_fd_sc_hd__a31oi_2 _27744_ (.A1(_05979_),
    .A2(_06007_),
    .A3(_05981_),
    .B1(_06128_),
    .Y(_06129_));
 sky130_fd_sc_hd__nand2_2 _27745_ (.A(_06127_),
    .B(_06129_),
    .Y(_06130_));
 sky130_vsdinv _27746_ (.A(_06128_),
    .Y(_06131_));
 sky130_fd_sc_hd__nand2_2 _27747_ (.A(_06009_),
    .B(_06131_),
    .Y(_06132_));
 sky130_fd_sc_hd__nand3_2 _27748_ (.A(_06132_),
    .B(_06123_),
    .C(_06126_),
    .Y(_06133_));
 sky130_fd_sc_hd__buf_1 _27749_ (.A(_06133_),
    .X(_06134_));
 sky130_fd_sc_hd__nand2_2 _27750_ (.A(_06130_),
    .B(_06134_),
    .Y(_06135_));
 sky130_fd_sc_hd__buf_1 _27751_ (.A(\pcpi_mul.rs2[9] ),
    .X(_06136_));
 sky130_fd_sc_hd__buf_1 _27752_ (.A(_06136_),
    .X(_06137_));
 sky130_fd_sc_hd__buf_1 _27753_ (.A(_06137_),
    .X(_06138_));
 sky130_fd_sc_hd__and2_2 _27754_ (.A(_06138_),
    .B(_05985_),
    .X(_06139_));
 sky130_fd_sc_hd__buf_1 _27755_ (.A(\pcpi_mul.rs2[10] ),
    .X(_06140_));
 sky130_fd_sc_hd__buf_1 _27756_ (.A(_06140_),
    .X(_06141_));
 sky130_fd_sc_hd__buf_1 _27757_ (.A(_06141_),
    .X(_06142_));
 sky130_fd_sc_hd__buf_1 _27758_ (.A(\pcpi_mul.rs1[1] ),
    .X(_06143_));
 sky130_fd_sc_hd__buf_1 _27759_ (.A(_06143_),
    .X(_06144_));
 sky130_fd_sc_hd__nand2_2 _27760_ (.A(_06142_),
    .B(_06144_),
    .Y(_06145_));
 sky130_fd_sc_hd__buf_1 _27761_ (.A(\pcpi_mul.rs2[11] ),
    .X(_06146_));
 sky130_fd_sc_hd__buf_1 _27762_ (.A(_06146_),
    .X(_06147_));
 sky130_fd_sc_hd__buf_1 _27763_ (.A(_06147_),
    .X(_06148_));
 sky130_fd_sc_hd__nand2_2 _27764_ (.A(_06148_),
    .B(_05239_),
    .Y(_06149_));
 sky130_fd_sc_hd__xnor2_2 _27765_ (.A(_06145_),
    .B(_06149_),
    .Y(_06150_));
 sky130_fd_sc_hd__xnor2_2 _27766_ (.A(_06139_),
    .B(_06150_),
    .Y(_06151_));
 sky130_vsdinv _27767_ (.A(_06151_),
    .Y(_06152_));
 sky130_fd_sc_hd__nand2_2 _27768_ (.A(_06135_),
    .B(_06152_),
    .Y(_06153_));
 sky130_fd_sc_hd__nand3_2 _27769_ (.A(_06130_),
    .B(_06151_),
    .C(_06133_),
    .Y(_06154_));
 sky130_fd_sc_hd__a21boi_2 _27770_ (.A1(_06153_),
    .A2(_06154_),
    .B1_N(_06020_),
    .Y(_06155_));
 sky130_fd_sc_hd__a21oi_2 _27771_ (.A1(_06130_),
    .A2(_06134_),
    .B1(_06151_),
    .Y(_06156_));
 sky130_vsdinv _27772_ (.A(_06154_),
    .Y(_06157_));
 sky130_fd_sc_hd__buf_1 _27773_ (.A(_06157_),
    .X(_06158_));
 sky130_fd_sc_hd__nor3_2 _27774_ (.A(_06021_),
    .B(_06156_),
    .C(_06158_),
    .Y(_06159_));
 sky130_fd_sc_hd__a21oi_2 _27775_ (.A1(_05980_),
    .A2(_05978_),
    .B1(_05975_),
    .Y(_06160_));
 sky130_fd_sc_hd__xor2_2 _27776_ (.A(_06160_),
    .B(_06012_),
    .X(_06161_));
 sky130_fd_sc_hd__o21bai_2 _27777_ (.A1(_06155_),
    .A2(_06159_),
    .B1_N(_06161_),
    .Y(_06162_));
 sky130_fd_sc_hd__o21ai_2 _27778_ (.A1(_06027_),
    .A2(_06022_),
    .B1(_06031_),
    .Y(_06163_));
 sky130_fd_sc_hd__o22ai_2 _27779_ (.A1(_06018_),
    .A2(_06014_),
    .B1(_06156_),
    .B2(_06158_),
    .Y(_06164_));
 sky130_fd_sc_hd__nand3b_2 _27780_ (.A_N(_06020_),
    .B(_06153_),
    .C(_06154_),
    .Y(_06165_));
 sky130_fd_sc_hd__nand3_2 _27781_ (.A(_06164_),
    .B(_06161_),
    .C(_06165_),
    .Y(_06166_));
 sky130_fd_sc_hd__nand3_2 _27782_ (.A(_06162_),
    .B(_06163_),
    .C(_06166_),
    .Y(_06167_));
 sky130_fd_sc_hd__a21oi_2 _27783_ (.A1(_06164_),
    .A2(_06165_),
    .B1(_06161_),
    .Y(_06168_));
 sky130_vsdinv _27784_ (.A(_06161_),
    .Y(_06169_));
 sky130_fd_sc_hd__nor3_2 _27785_ (.A(_06169_),
    .B(_06155_),
    .C(_06159_),
    .Y(_06170_));
 sky130_fd_sc_hd__o21bai_2 _27786_ (.A1(_06168_),
    .A2(_06170_),
    .B1_N(_06163_),
    .Y(_06171_));
 sky130_fd_sc_hd__o2bb2ai_2 _27787_ (.A1_N(_06167_),
    .A2_N(_06171_),
    .B1(_05902_),
    .B2(_06026_),
    .Y(_06172_));
 sky130_fd_sc_hd__nor2_2 _27788_ (.A(_06026_),
    .B(_05902_),
    .Y(_06173_));
 sky130_fd_sc_hd__nand3_2 _27789_ (.A(_06171_),
    .B(_06173_),
    .C(_06167_),
    .Y(_06174_));
 sky130_fd_sc_hd__a21oi_2 _27790_ (.A1(_06172_),
    .A2(_06174_),
    .B1(_06035_),
    .Y(_06175_));
 sky130_vsdinv _27791_ (.A(_06035_),
    .Y(_06176_));
 sky130_fd_sc_hd__a21oi_2 _27792_ (.A1(_06171_),
    .A2(_06167_),
    .B1(_06173_),
    .Y(_06177_));
 sky130_fd_sc_hd__nor3b_2 _27793_ (.A(_06176_),
    .B(_06177_),
    .C_N(_06174_),
    .Y(_06178_));
 sky130_fd_sc_hd__nor2_2 _27794_ (.A(_06175_),
    .B(_06178_),
    .Y(_06179_));
 sky130_fd_sc_hd__xnor2_2 _27795_ (.A(_06039_),
    .B(_06179_),
    .Y(_02630_));
 sky130_fd_sc_hd__buf_1 _27796_ (.A(_19267_),
    .X(_06180_));
 sky130_fd_sc_hd__buf_1 _27797_ (.A(_06074_),
    .X(_06181_));
 sky130_fd_sc_hd__a22oi_2 _27798_ (.A1(_05513_),
    .A2(_06180_),
    .B1(_05509_),
    .B2(_06181_),
    .Y(_06182_));
 sky130_fd_sc_hd__nand2_2 _27799_ (.A(_05491_),
    .B(_05963_),
    .Y(_06183_));
 sky130_fd_sc_hd__nand2_2 _27800_ (.A(_05652_),
    .B(_05847_),
    .Y(_06184_));
 sky130_fd_sc_hd__nor2_2 _27801_ (.A(_06183_),
    .B(_06184_),
    .Y(_06185_));
 sky130_fd_sc_hd__buf_1 _27802_ (.A(_19241_),
    .X(_06186_));
 sky130_fd_sc_hd__buf_1 _27803_ (.A(_06186_),
    .X(_06187_));
 sky130_fd_sc_hd__and2_2 _27804_ (.A(_05516_),
    .B(_06187_),
    .X(_06188_));
 sky130_fd_sc_hd__o21bai_2 _27805_ (.A1(_06182_),
    .A2(_06185_),
    .B1_N(_06188_),
    .Y(_06189_));
 sky130_fd_sc_hd__nand3b_2 _27806_ (.A_N(_06183_),
    .B(_18850_),
    .C(_05954_),
    .Y(_06190_));
 sky130_fd_sc_hd__nand3b_2 _27807_ (.A_N(_06182_),
    .B(_06190_),
    .C(_06188_),
    .Y(_06191_));
 sky130_fd_sc_hd__nand2_2 _27808_ (.A(_06189_),
    .B(_06191_),
    .Y(_06192_));
 sky130_fd_sc_hd__a21oi_2 _27809_ (.A1(_06049_),
    .A2(_06048_),
    .B1(_06045_),
    .Y(_06193_));
 sky130_fd_sc_hd__nand2_2 _27810_ (.A(_06192_),
    .B(_06193_),
    .Y(_06194_));
 sky130_fd_sc_hd__nand3b_2 _27811_ (.A_N(_06193_),
    .B(_06191_),
    .C(_06189_),
    .Y(_06195_));
 sky130_fd_sc_hd__nand2_2 _27812_ (.A(_06194_),
    .B(_06195_),
    .Y(_06196_));
 sky130_fd_sc_hd__buf_1 _27813_ (.A(_06047_),
    .X(_06197_));
 sky130_fd_sc_hd__a22oi_2 _27814_ (.A1(_05953_),
    .A2(_06064_),
    .B1(_05554_),
    .B2(_06197_),
    .Y(_06198_));
 sky130_fd_sc_hd__buf_1 _27815_ (.A(_06068_),
    .X(_06199_));
 sky130_fd_sc_hd__nand2_2 _27816_ (.A(_05662_),
    .B(_06199_),
    .Y(_06200_));
 sky130_fd_sc_hd__buf_1 _27817_ (.A(\pcpi_mul.rs1[11] ),
    .X(_06201_));
 sky130_fd_sc_hd__buf_1 _27818_ (.A(_06201_),
    .X(_06202_));
 sky130_fd_sc_hd__buf_1 _27819_ (.A(_06202_),
    .X(_06203_));
 sky130_fd_sc_hd__nand2_2 _27820_ (.A(_05663_),
    .B(_06203_),
    .Y(_06204_));
 sky130_fd_sc_hd__nor2_2 _27821_ (.A(_06200_),
    .B(_06204_),
    .Y(_06205_));
 sky130_fd_sc_hd__and2_2 _27822_ (.A(_06073_),
    .B(_05822_),
    .X(_06206_));
 sky130_fd_sc_hd__nor3b_2 _27823_ (.A(_06198_),
    .B(_06205_),
    .C_N(_06206_),
    .Y(_06207_));
 sky130_fd_sc_hd__o21ba_2 _27824_ (.A1(_06198_),
    .A2(_06205_),
    .B1_N(_06206_),
    .X(_06208_));
 sky130_fd_sc_hd__nor2_2 _27825_ (.A(_06207_),
    .B(_06208_),
    .Y(_06209_));
 sky130_vsdinv _27826_ (.A(_06209_),
    .Y(_06210_));
 sky130_fd_sc_hd__nand2_2 _27827_ (.A(_06196_),
    .B(_06210_),
    .Y(_06211_));
 sky130_fd_sc_hd__nand3_2 _27828_ (.A(_06194_),
    .B(_06209_),
    .C(_06195_),
    .Y(_06212_));
 sky130_fd_sc_hd__a21boi_2 _27829_ (.A1(_06050_),
    .A2(_06054_),
    .B1_N(_06056_),
    .Y(_06213_));
 sky130_fd_sc_hd__o21ai_2 _27830_ (.A1(_06079_),
    .A2(_06213_),
    .B1(_06058_),
    .Y(_06214_));
 sky130_fd_sc_hd__a21oi_2 _27831_ (.A1(_06211_),
    .A2(_06212_),
    .B1(_06214_),
    .Y(_06215_));
 sky130_fd_sc_hd__nand3_2 _27832_ (.A(_06211_),
    .B(_06214_),
    .C(_06212_),
    .Y(_06216_));
 sky130_vsdinv _27833_ (.A(_06216_),
    .Y(_06217_));
 sky130_fd_sc_hd__o31a_2 _27834_ (.A1(_05690_),
    .A2(_19263_),
    .A3(_06065_),
    .B1(_06072_),
    .X(_06218_));
 sky130_fd_sc_hd__o21ai_2 _27835_ (.A1(_06215_),
    .A2(_06217_),
    .B1(_06218_),
    .Y(_06219_));
 sky130_fd_sc_hd__a21o_2 _27836_ (.A1(_06211_),
    .A2(_06212_),
    .B1(_06214_),
    .X(_06220_));
 sky130_fd_sc_hd__nand3b_2 _27837_ (.A_N(_06218_),
    .B(_06220_),
    .C(_06216_),
    .Y(_06221_));
 sky130_fd_sc_hd__nand2_2 _27838_ (.A(_06219_),
    .B(_06221_),
    .Y(_06222_));
 sky130_fd_sc_hd__nand3_2 _27839_ (.A(_06117_),
    .B(_06118_),
    .C(_06093_),
    .Y(_06223_));
 sky130_fd_sc_hd__buf_1 _27840_ (.A(_05771_),
    .X(_06224_));
 sky130_fd_sc_hd__buf_1 _27841_ (.A(_06224_),
    .X(_06225_));
 sky130_fd_sc_hd__buf_1 _27842_ (.A(_18832_),
    .X(_06226_));
 sky130_fd_sc_hd__buf_1 _27843_ (.A(_06226_),
    .X(_06227_));
 sky130_fd_sc_hd__a22oi_2 _27844_ (.A1(_06225_),
    .A2(_05556_),
    .B1(_06227_),
    .B2(_05827_),
    .Y(_06228_));
 sky130_fd_sc_hd__nand2_2 _27845_ (.A(_18829_),
    .B(_05733_),
    .Y(_06229_));
 sky130_fd_sc_hd__buf_1 _27846_ (.A(_05872_),
    .X(_06230_));
 sky130_fd_sc_hd__buf_1 _27847_ (.A(_06230_),
    .X(_06231_));
 sky130_fd_sc_hd__buf_1 _27848_ (.A(_05529_),
    .X(_06232_));
 sky130_fd_sc_hd__nand2_2 _27849_ (.A(_06231_),
    .B(_06232_),
    .Y(_06233_));
 sky130_fd_sc_hd__nor2_2 _27850_ (.A(_06229_),
    .B(_06233_),
    .Y(_06234_));
 sky130_fd_sc_hd__and2_2 _27851_ (.A(_05587_),
    .B(_05852_),
    .X(_06235_));
 sky130_fd_sc_hd__o21bai_2 _27852_ (.A1(_06228_),
    .A2(_06234_),
    .B1_N(_06235_),
    .Y(_06236_));
 sky130_fd_sc_hd__buf_1 _27853_ (.A(_05992_),
    .X(_06237_));
 sky130_fd_sc_hd__buf_1 _27854_ (.A(_06237_),
    .X(_06238_));
 sky130_fd_sc_hd__nand3b_2 _27855_ (.A_N(_06229_),
    .B(_06238_),
    .C(_06232_),
    .Y(_06239_));
 sky130_fd_sc_hd__nand3b_2 _27856_ (.A_N(_06228_),
    .B(_06239_),
    .C(_06235_),
    .Y(_06240_));
 sky130_fd_sc_hd__nand2_2 _27857_ (.A(_06236_),
    .B(_06240_),
    .Y(_06241_));
 sky130_fd_sc_hd__nand2_2 _27858_ (.A(_06145_),
    .B(_06149_),
    .Y(_06242_));
 sky130_fd_sc_hd__nor2_2 _27859_ (.A(_06145_),
    .B(_06149_),
    .Y(_06243_));
 sky130_fd_sc_hd__a21oi_2 _27860_ (.A1(_06242_),
    .A2(_06139_),
    .B1(_06243_),
    .Y(_06244_));
 sky130_fd_sc_hd__nand2_2 _27861_ (.A(_06241_),
    .B(_06244_),
    .Y(_06245_));
 sky130_fd_sc_hd__nand3b_2 _27862_ (.A_N(_06244_),
    .B(_06240_),
    .C(_06236_),
    .Y(_06246_));
 sky130_fd_sc_hd__nand2_2 _27863_ (.A(_06245_),
    .B(_06246_),
    .Y(_06247_));
 sky130_fd_sc_hd__buf_1 _27864_ (.A(_18840_),
    .X(_06248_));
 sky130_fd_sc_hd__o31a_2 _27865_ (.A1(_06248_),
    .A2(_19279_),
    .A3(_06098_),
    .B1(_06107_),
    .X(_06249_));
 sky130_fd_sc_hd__nand2_2 _27866_ (.A(_06247_),
    .B(_06249_),
    .Y(_06250_));
 sky130_fd_sc_hd__nand3b_2 _27867_ (.A_N(_06249_),
    .B(_06245_),
    .C(_06246_),
    .Y(_06251_));
 sky130_fd_sc_hd__o21ai_2 _27868_ (.A1(_06115_),
    .A2(_06110_),
    .B1(_06111_),
    .Y(_06252_));
 sky130_fd_sc_hd__a21o_2 _27869_ (.A1(_06250_),
    .A2(_06251_),
    .B1(_06252_),
    .X(_06253_));
 sky130_fd_sc_hd__nand3_2 _27870_ (.A(_06250_),
    .B(_06252_),
    .C(_06251_),
    .Y(_06254_));
 sky130_fd_sc_hd__nand3b_2 _27871_ (.A_N(_06223_),
    .B(_06253_),
    .C(_06254_),
    .Y(_06255_));
 sky130_fd_sc_hd__o2bb2ai_2 _27872_ (.A1_N(_06254_),
    .A2_N(_06253_),
    .B1(_06004_),
    .B2(_06119_),
    .Y(_06256_));
 sky130_fd_sc_hd__nand3b_2 _27873_ (.A_N(_06222_),
    .B(_06255_),
    .C(_06256_),
    .Y(_06257_));
 sky130_fd_sc_hd__nand2_2 _27874_ (.A(_06256_),
    .B(_06255_),
    .Y(_06258_));
 sky130_fd_sc_hd__nand2_2 _27875_ (.A(_06258_),
    .B(_06222_),
    .Y(_06259_));
 sky130_fd_sc_hd__nand3_2 _27876_ (.A(_06094_),
    .B(_06118_),
    .C(_06117_),
    .Y(_06260_));
 sky130_fd_sc_hd__nand2_2 _27877_ (.A(_06126_),
    .B(_06260_),
    .Y(_06261_));
 sky130_fd_sc_hd__nand3_2 _27878_ (.A(_06257_),
    .B(_06259_),
    .C(_06261_),
    .Y(_06262_));
 sky130_fd_sc_hd__buf_1 _27879_ (.A(_06262_),
    .X(_06263_));
 sky130_fd_sc_hd__a22oi_2 _27880_ (.A1(_06219_),
    .A2(_06221_),
    .B1(_06256_),
    .B2(_06255_),
    .Y(_06264_));
 sky130_fd_sc_hd__nor2_2 _27881_ (.A(_06222_),
    .B(_06258_),
    .Y(_06265_));
 sky130_fd_sc_hd__o21bai_2 _27882_ (.A1(_06264_),
    .A2(_06265_),
    .B1_N(_06261_),
    .Y(_06266_));
 sky130_fd_sc_hd__nand2_2 _27883_ (.A(_18815_),
    .B(_05425_),
    .Y(_06267_));
 sky130_fd_sc_hd__buf_1 _27884_ (.A(_18819_),
    .X(_06268_));
 sky130_fd_sc_hd__nand2_2 _27885_ (.A(_06268_),
    .B(_05985_),
    .Y(_06269_));
 sky130_fd_sc_hd__nand2_2 _27886_ (.A(_06267_),
    .B(_06269_),
    .Y(_06270_));
 sky130_fd_sc_hd__nor2_2 _27887_ (.A(_06267_),
    .B(_06269_),
    .Y(_06271_));
 sky130_vsdinv _27888_ (.A(_06271_),
    .Y(_06272_));
 sky130_fd_sc_hd__o2bb2ai_2 _27889_ (.A1_N(_06270_),
    .A2_N(_06272_),
    .B1(_18825_),
    .B2(_19290_),
    .Y(_06273_));
 sky130_fd_sc_hd__buf_1 _27890_ (.A(_18807_),
    .X(_06274_));
 sky130_fd_sc_hd__buf_1 _27891_ (.A(_06274_),
    .X(_06275_));
 sky130_fd_sc_hd__buf_1 _27892_ (.A(_06275_),
    .X(_06276_));
 sky130_fd_sc_hd__and2_2 _27893_ (.A(_06276_),
    .B(_05241_),
    .X(_06277_));
 sky130_fd_sc_hd__and2_2 _27894_ (.A(_05896_),
    .B(_05988_),
    .X(_06278_));
 sky130_fd_sc_hd__nand3b_2 _27895_ (.A_N(_06271_),
    .B(_06278_),
    .C(_06270_),
    .Y(_06279_));
 sky130_fd_sc_hd__nand3_2 _27896_ (.A(_06273_),
    .B(_06277_),
    .C(_06279_),
    .Y(_06280_));
 sky130_vsdinv _27897_ (.A(_06280_),
    .Y(_06281_));
 sky130_fd_sc_hd__a21oi_2 _27898_ (.A1(_06273_),
    .A2(_06279_),
    .B1(_06277_),
    .Y(_06282_));
 sky130_fd_sc_hd__o2bb2ai_2 _27899_ (.A1_N(_06263_),
    .A2_N(_06266_),
    .B1(_06281_),
    .B2(_06282_),
    .Y(_06283_));
 sky130_fd_sc_hd__nor2_2 _27900_ (.A(_06282_),
    .B(_06281_),
    .Y(_06284_));
 sky130_fd_sc_hd__nand3_2 _27901_ (.A(_06266_),
    .B(_06262_),
    .C(_06284_),
    .Y(_06285_));
 sky130_fd_sc_hd__a21oi_2 _27902_ (.A1(_06283_),
    .A2(_06285_),
    .B1(_06158_),
    .Y(_06286_));
 sky130_fd_sc_hd__a21oi_2 _27903_ (.A1(_06266_),
    .A2(_06263_),
    .B1(_06284_),
    .Y(_06287_));
 sky130_vsdinv _27904_ (.A(_06285_),
    .Y(_06288_));
 sky130_fd_sc_hd__buf_1 _27905_ (.A(_06288_),
    .X(_06289_));
 sky130_fd_sc_hd__nor3_2 _27906_ (.A(_06154_),
    .B(_06287_),
    .C(_06289_),
    .Y(_06290_));
 sky130_fd_sc_hd__a21boi_2 _27907_ (.A1(_06086_),
    .A2(_06089_),
    .B1_N(_06087_),
    .Y(_06291_));
 sky130_fd_sc_hd__xor2_2 _27908_ (.A(_06291_),
    .B(_06134_),
    .X(_06292_));
 sky130_fd_sc_hd__o21bai_2 _27909_ (.A1(_06286_),
    .A2(_06290_),
    .B1_N(_06292_),
    .Y(_06293_));
 sky130_fd_sc_hd__o21ai_2 _27910_ (.A1(_06169_),
    .A2(_06155_),
    .B1(_06165_),
    .Y(_06294_));
 sky130_fd_sc_hd__o21bai_2 _27911_ (.A1(_06287_),
    .A2(_06288_),
    .B1_N(_06157_),
    .Y(_06295_));
 sky130_fd_sc_hd__nand3_2 _27912_ (.A(_06283_),
    .B(_06158_),
    .C(_06285_),
    .Y(_06296_));
 sky130_fd_sc_hd__nand3_2 _27913_ (.A(_06295_),
    .B(_06296_),
    .C(_06292_),
    .Y(_06297_));
 sky130_fd_sc_hd__nand3_2 _27914_ (.A(_06293_),
    .B(_06294_),
    .C(_06297_),
    .Y(_06298_));
 sky130_fd_sc_hd__nand2_2 _27915_ (.A(_06293_),
    .B(_06297_),
    .Y(_06299_));
 sky130_vsdinv _27916_ (.A(_06294_),
    .Y(_06300_));
 sky130_fd_sc_hd__nand2_2 _27917_ (.A(_06299_),
    .B(_06300_),
    .Y(_06301_));
 sky130_fd_sc_hd__o2bb2ai_2 _27918_ (.A1_N(_06298_),
    .A2_N(_06301_),
    .B1(_06013_),
    .B2(_06160_),
    .Y(_06302_));
 sky130_fd_sc_hd__nor2_2 _27919_ (.A(_06160_),
    .B(_06013_),
    .Y(_06303_));
 sky130_fd_sc_hd__nand3_2 _27920_ (.A(_06301_),
    .B(_06303_),
    .C(_06298_),
    .Y(_06304_));
 sky130_fd_sc_hd__a21boi_2 _27921_ (.A1(_06171_),
    .A2(_06173_),
    .B1_N(_06167_),
    .Y(_06305_));
 sky130_fd_sc_hd__a21boi_2 _27922_ (.A1(_06302_),
    .A2(_06304_),
    .B1_N(_06305_),
    .Y(_06306_));
 sky130_fd_sc_hd__a21oi_2 _27923_ (.A1(_06301_),
    .A2(_06298_),
    .B1(_06303_),
    .Y(_06307_));
 sky130_fd_sc_hd__nor3b_2 _27924_ (.A(_06305_),
    .B(_06307_),
    .C_N(_06304_),
    .Y(_06308_));
 sky130_fd_sc_hd__nor2_2 _27925_ (.A(_06306_),
    .B(_06308_),
    .Y(_06309_));
 sky130_fd_sc_hd__o21bai_2 _27926_ (.A1(_06175_),
    .A2(_06039_),
    .B1_N(_06178_),
    .Y(_06310_));
 sky130_fd_sc_hd__xor2_2 _27927_ (.A(_06309_),
    .B(_06310_),
    .X(_02631_));
 sky130_fd_sc_hd__buf_1 _27928_ (.A(_06224_),
    .X(_06311_));
 sky130_fd_sc_hd__nand2_2 _27929_ (.A(_06311_),
    .B(_05827_),
    .Y(_06312_));
 sky130_fd_sc_hd__nand2_2 _27930_ (.A(_06238_),
    .B(_05941_),
    .Y(_06313_));
 sky130_fd_sc_hd__nand2_2 _27931_ (.A(_06312_),
    .B(_06313_),
    .Y(_06314_));
 sky130_fd_sc_hd__nand3b_2 _27932_ (.A_N(_06312_),
    .B(_18835_),
    .C(_05941_),
    .Y(_06315_));
 sky130_fd_sc_hd__o2bb2ai_2 _27933_ (.A1_N(_06314_),
    .A2_N(_06315_),
    .B1(_18841_),
    .B2(_19269_),
    .Y(_06316_));
 sky130_fd_sc_hd__buf_1 _27934_ (.A(_05838_),
    .X(_06317_));
 sky130_fd_sc_hd__and2_2 _27935_ (.A(_05588_),
    .B(_06317_),
    .X(_06318_));
 sky130_fd_sc_hd__nand3_2 _27936_ (.A(_06315_),
    .B(_06318_),
    .C(_06314_),
    .Y(_06319_));
 sky130_fd_sc_hd__a21oi_2 _27937_ (.A1(_06270_),
    .A2(_06278_),
    .B1(_06271_),
    .Y(_06320_));
 sky130_vsdinv _27938_ (.A(_06320_),
    .Y(_06321_));
 sky130_fd_sc_hd__a21o_2 _27939_ (.A1(_06316_),
    .A2(_06319_),
    .B1(_06321_),
    .X(_06322_));
 sky130_fd_sc_hd__nand3_2 _27940_ (.A(_06316_),
    .B(_06321_),
    .C(_06319_),
    .Y(_06323_));
 sky130_fd_sc_hd__o31a_2 _27941_ (.A1(_06248_),
    .A2(_19275_),
    .A3(_06228_),
    .B1(_06239_),
    .X(_06324_));
 sky130_vsdinv _27942_ (.A(_06324_),
    .Y(_06325_));
 sky130_fd_sc_hd__a21o_2 _27943_ (.A1(_06322_),
    .A2(_06323_),
    .B1(_06325_),
    .X(_06326_));
 sky130_fd_sc_hd__nand3_2 _27944_ (.A(_06322_),
    .B(_06325_),
    .C(_06323_),
    .Y(_06327_));
 sky130_fd_sc_hd__nand2_2 _27945_ (.A(_06326_),
    .B(_06327_),
    .Y(_06328_));
 sky130_fd_sc_hd__nand2_2 _27946_ (.A(_06328_),
    .B(_06280_),
    .Y(_06329_));
 sky130_fd_sc_hd__nand3_2 _27947_ (.A(_06326_),
    .B(_06281_),
    .C(_06327_),
    .Y(_06330_));
 sky130_fd_sc_hd__nand2_2 _27948_ (.A(_06329_),
    .B(_06330_),
    .Y(_06331_));
 sky130_fd_sc_hd__o21a_2 _27949_ (.A1(_06244_),
    .A2(_06241_),
    .B1(_06251_),
    .X(_06332_));
 sky130_fd_sc_hd__nand2_2 _27950_ (.A(_06331_),
    .B(_06332_),
    .Y(_06333_));
 sky130_fd_sc_hd__nand3b_2 _27951_ (.A_N(_06332_),
    .B(_06329_),
    .C(_06330_),
    .Y(_06334_));
 sky130_fd_sc_hd__nand2_2 _27952_ (.A(_06333_),
    .B(_06334_),
    .Y(_06335_));
 sky130_fd_sc_hd__nand2_2 _27953_ (.A(_06335_),
    .B(_06254_),
    .Y(_06336_));
 sky130_vsdinv _27954_ (.A(_06254_),
    .Y(_06337_));
 sky130_fd_sc_hd__nand3_2 _27955_ (.A(_06333_),
    .B(_06337_),
    .C(_06334_),
    .Y(_06338_));
 sky130_fd_sc_hd__nand2_2 _27956_ (.A(_06051_),
    .B(_05954_),
    .Y(_06339_));
 sky130_fd_sc_hd__nand2_2 _27957_ (.A(_05652_),
    .B(_06061_),
    .Y(_06340_));
 sky130_fd_sc_hd__nand2_2 _27958_ (.A(_06339_),
    .B(_06340_),
    .Y(_06341_));
 sky130_fd_sc_hd__buf_1 _27959_ (.A(_05957_),
    .X(_06342_));
 sky130_fd_sc_hd__buf_1 _27960_ (.A(_06342_),
    .X(_06343_));
 sky130_fd_sc_hd__buf_1 _27961_ (.A(_06343_),
    .X(_06344_));
 sky130_fd_sc_hd__nand3b_2 _27962_ (.A_N(_06339_),
    .B(_18851_),
    .C(_06344_),
    .Y(_06345_));
 sky130_fd_sc_hd__buf_1 _27963_ (.A(_18879_),
    .X(_06346_));
 sky130_fd_sc_hd__buf_1 _27964_ (.A(_06346_),
    .X(_06347_));
 sky130_fd_sc_hd__o2bb2ai_2 _27965_ (.A1_N(_06341_),
    .A2_N(_06345_),
    .B1(_06347_),
    .B2(_19239_),
    .Y(_06348_));
 sky130_fd_sc_hd__buf_1 _27966_ (.A(_05235_),
    .X(_06349_));
 sky130_fd_sc_hd__buf_1 _27967_ (.A(_19236_),
    .X(_06350_));
 sky130_fd_sc_hd__buf_1 _27968_ (.A(_06350_),
    .X(_06351_));
 sky130_fd_sc_hd__and2_2 _27969_ (.A(_06349_),
    .B(_06351_),
    .X(_06352_));
 sky130_fd_sc_hd__nand3_2 _27970_ (.A(_06345_),
    .B(_06352_),
    .C(_06341_),
    .Y(_06353_));
 sky130_fd_sc_hd__o31ai_2 _27971_ (.A1(_06347_),
    .A2(_19244_),
    .A3(_06182_),
    .B1(_06190_),
    .Y(_06354_));
 sky130_fd_sc_hd__a21o_2 _27972_ (.A1(_06348_),
    .A2(_06353_),
    .B1(_06354_),
    .X(_06355_));
 sky130_fd_sc_hd__nand3_2 _27973_ (.A(_06354_),
    .B(_06348_),
    .C(_06353_),
    .Y(_06356_));
 sky130_fd_sc_hd__buf_1 _27974_ (.A(_06062_),
    .X(_06357_));
 sky130_fd_sc_hd__buf_1 _27975_ (.A(_06357_),
    .X(_06358_));
 sky130_fd_sc_hd__and2_2 _27976_ (.A(_05460_),
    .B(_06358_),
    .X(_06359_));
 sky130_fd_sc_hd__buf_1 _27977_ (.A(_06202_),
    .X(_06360_));
 sky130_fd_sc_hd__buf_1 _27978_ (.A(_06360_),
    .X(_06361_));
 sky130_fd_sc_hd__nand2_2 _27979_ (.A(_05422_),
    .B(_06361_),
    .Y(_06362_));
 sky130_fd_sc_hd__buf_1 _27980_ (.A(_05663_),
    .X(_06363_));
 sky130_fd_sc_hd__buf_1 _27981_ (.A(_19241_),
    .X(_06364_));
 sky130_fd_sc_hd__buf_1 _27982_ (.A(_06364_),
    .X(_06365_));
 sky130_fd_sc_hd__buf_1 _27983_ (.A(_06365_),
    .X(_06366_));
 sky130_fd_sc_hd__nand2_2 _27984_ (.A(_06363_),
    .B(_06366_),
    .Y(_06367_));
 sky130_fd_sc_hd__xnor2_2 _27985_ (.A(_06362_),
    .B(_06367_),
    .Y(_06368_));
 sky130_fd_sc_hd__xnor2_2 _27986_ (.A(_06359_),
    .B(_06368_),
    .Y(_06369_));
 sky130_fd_sc_hd__a21oi_2 _27987_ (.A1(_06355_),
    .A2(_06356_),
    .B1(_06369_),
    .Y(_06370_));
 sky130_fd_sc_hd__nand3_2 _27988_ (.A(_06369_),
    .B(_06355_),
    .C(_06356_),
    .Y(_06371_));
 sky130_vsdinv _27989_ (.A(_06371_),
    .Y(_06372_));
 sky130_fd_sc_hd__a21boi_2 _27990_ (.A1(_06194_),
    .A2(_06209_),
    .B1_N(_06195_),
    .Y(_06373_));
 sky130_vsdinv _27991_ (.A(_06373_),
    .Y(_06374_));
 sky130_fd_sc_hd__o21bai_2 _27992_ (.A1(_06370_),
    .A2(_06372_),
    .B1_N(_06374_),
    .Y(_06375_));
 sky130_fd_sc_hd__nand3b_2 _27993_ (.A_N(_06370_),
    .B(_06371_),
    .C(_06374_),
    .Y(_06376_));
 sky130_fd_sc_hd__nor2_2 _27994_ (.A(_06205_),
    .B(_06207_),
    .Y(_06377_));
 sky130_vsdinv _27995_ (.A(_06377_),
    .Y(_06378_));
 sky130_fd_sc_hd__a21oi_2 _27996_ (.A1(_06375_),
    .A2(_06376_),
    .B1(_06378_),
    .Y(_06379_));
 sky130_fd_sc_hd__nand3_2 _27997_ (.A(_06375_),
    .B(_06378_),
    .C(_06376_),
    .Y(_06380_));
 sky130_vsdinv _27998_ (.A(_06380_),
    .Y(_06381_));
 sky130_fd_sc_hd__nor2_2 _27999_ (.A(_06379_),
    .B(_06381_),
    .Y(_06382_));
 sky130_fd_sc_hd__a21oi_2 _28000_ (.A1(_06336_),
    .A2(_06338_),
    .B1(_06382_),
    .Y(_06383_));
 sky130_fd_sc_hd__nand3_2 _28001_ (.A(_06336_),
    .B(_06382_),
    .C(_06338_),
    .Y(_06384_));
 sky130_vsdinv _28002_ (.A(_06384_),
    .Y(_06385_));
 sky130_vsdinv _28003_ (.A(_06255_),
    .Y(_06386_));
 sky130_fd_sc_hd__a31oi_2 _28004_ (.A1(_06256_),
    .A2(_06219_),
    .A3(_06221_),
    .B1(_06386_),
    .Y(_06387_));
 sky130_vsdinv _28005_ (.A(_06387_),
    .Y(_06388_));
 sky130_fd_sc_hd__o21bai_2 _28006_ (.A1(_06383_),
    .A2(_06385_),
    .B1_N(_06388_),
    .Y(_06389_));
 sky130_fd_sc_hd__o2bb2ai_2 _28007_ (.A1_N(_06338_),
    .A2_N(_06336_),
    .B1(_06381_),
    .B2(_06379_),
    .Y(_06390_));
 sky130_fd_sc_hd__nand3_2 _28008_ (.A(_06390_),
    .B(_06388_),
    .C(_06384_),
    .Y(_06391_));
 sky130_fd_sc_hd__buf_1 _28009_ (.A(_18801_),
    .X(_06392_));
 sky130_fd_sc_hd__buf_1 _28010_ (.A(_06392_),
    .X(_06393_));
 sky130_fd_sc_hd__buf_1 _28011_ (.A(_06393_),
    .X(_06394_));
 sky130_fd_sc_hd__nand2_2 _28012_ (.A(_06394_),
    .B(_05466_),
    .Y(_06395_));
 sky130_fd_sc_hd__nand2_2 _28013_ (.A(_06276_),
    .B(_05568_),
    .Y(_06396_));
 sky130_fd_sc_hd__xor2_2 _28014_ (.A(_06395_),
    .B(_06396_),
    .X(_06397_));
 sky130_fd_sc_hd__nand2_2 _28015_ (.A(_06148_),
    .B(_05985_),
    .Y(_06398_));
 sky130_fd_sc_hd__nand2_2 _28016_ (.A(_06268_),
    .B(_05552_),
    .Y(_06399_));
 sky130_fd_sc_hd__nand2_2 _28017_ (.A(_06398_),
    .B(_06399_),
    .Y(_06400_));
 sky130_fd_sc_hd__nor2_2 _28018_ (.A(_06398_),
    .B(_06399_),
    .Y(_06401_));
 sky130_vsdinv _28019_ (.A(_06401_),
    .Y(_06402_));
 sky130_fd_sc_hd__o2bb2ai_2 _28020_ (.A1_N(_06400_),
    .A2_N(_06402_),
    .B1(_18825_),
    .B2(_19283_),
    .Y(_06403_));
 sky130_fd_sc_hd__and2_2 _28021_ (.A(_06138_),
    .B(_05471_),
    .X(_06404_));
 sky130_fd_sc_hd__nand3b_2 _28022_ (.A_N(_06401_),
    .B(_06404_),
    .C(_06400_),
    .Y(_06405_));
 sky130_fd_sc_hd__nand2_2 _28023_ (.A(_06403_),
    .B(_06405_),
    .Y(_06406_));
 sky130_fd_sc_hd__xnor2_2 _28024_ (.A(_06397_),
    .B(_06406_),
    .Y(_06407_));
 sky130_fd_sc_hd__a21oi_2 _28025_ (.A1(_06389_),
    .A2(_06391_),
    .B1(_06407_),
    .Y(_06408_));
 sky130_vsdinv _28026_ (.A(_06407_),
    .Y(_06409_));
 sky130_fd_sc_hd__a21oi_2 _28027_ (.A1(_06390_),
    .A2(_06384_),
    .B1(_06388_),
    .Y(_06410_));
 sky130_fd_sc_hd__nor3_2 _28028_ (.A(_06387_),
    .B(_06383_),
    .C(_06385_),
    .Y(_06411_));
 sky130_fd_sc_hd__nor3_2 _28029_ (.A(_06409_),
    .B(_06410_),
    .C(_06411_),
    .Y(_06412_));
 sky130_fd_sc_hd__o21bai_2 _28030_ (.A1(_06408_),
    .A2(_06412_),
    .B1_N(_06289_),
    .Y(_06413_));
 sky130_fd_sc_hd__o21bai_2 _28031_ (.A1(_06410_),
    .A2(_06411_),
    .B1_N(_06407_),
    .Y(_06414_));
 sky130_fd_sc_hd__nand3_2 _28032_ (.A(_06389_),
    .B(_06407_),
    .C(_06391_),
    .Y(_06415_));
 sky130_fd_sc_hd__nand3_2 _28033_ (.A(_06414_),
    .B(_06289_),
    .C(_06415_),
    .Y(_06416_));
 sky130_fd_sc_hd__o21a_2 _28034_ (.A1(_06218_),
    .A2(_06215_),
    .B1(_06216_),
    .X(_06417_));
 sky130_fd_sc_hd__xor2_2 _28035_ (.A(_06417_),
    .B(_06263_),
    .X(_06418_));
 sky130_fd_sc_hd__a21oi_2 _28036_ (.A1(_06413_),
    .A2(_06416_),
    .B1(_06418_),
    .Y(_06419_));
 sky130_vsdinv _28037_ (.A(_06418_),
    .Y(_06420_));
 sky130_fd_sc_hd__a21oi_2 _28038_ (.A1(_06414_),
    .A2(_06415_),
    .B1(_06289_),
    .Y(_06421_));
 sky130_fd_sc_hd__nor3_2 _28039_ (.A(_06285_),
    .B(_06408_),
    .C(_06412_),
    .Y(_06422_));
 sky130_fd_sc_hd__nor3_2 _28040_ (.A(_06420_),
    .B(_06421_),
    .C(_06422_),
    .Y(_06423_));
 sky130_fd_sc_hd__a21o_2 _28041_ (.A1(_06295_),
    .A2(_06292_),
    .B1(_06290_),
    .X(_06424_));
 sky130_fd_sc_hd__o21bai_2 _28042_ (.A1(_06419_),
    .A2(_06423_),
    .B1_N(_06424_),
    .Y(_06425_));
 sky130_fd_sc_hd__o21bai_2 _28043_ (.A1(_06421_),
    .A2(_06422_),
    .B1_N(_06418_),
    .Y(_06426_));
 sky130_fd_sc_hd__nand3_2 _28044_ (.A(_06413_),
    .B(_06416_),
    .C(_06418_),
    .Y(_06427_));
 sky130_fd_sc_hd__nand3_2 _28045_ (.A(_06426_),
    .B(_06427_),
    .C(_06424_),
    .Y(_06428_));
 sky130_fd_sc_hd__nor2_2 _28046_ (.A(_06291_),
    .B(_06134_),
    .Y(_06429_));
 sky130_fd_sc_hd__buf_1 _28047_ (.A(_06429_),
    .X(_06430_));
 sky130_fd_sc_hd__a21oi_2 _28048_ (.A1(_06425_),
    .A2(_06428_),
    .B1(_06430_),
    .Y(_06431_));
 sky130_vsdinv _28049_ (.A(_06429_),
    .Y(_06432_));
 sky130_fd_sc_hd__a21oi_2 _28050_ (.A1(_06426_),
    .A2(_06427_),
    .B1(_06424_),
    .Y(_06433_));
 sky130_vsdinv _28051_ (.A(_06428_),
    .Y(_06434_));
 sky130_fd_sc_hd__nor3_2 _28052_ (.A(_06432_),
    .B(_06433_),
    .C(_06434_),
    .Y(_06435_));
 sky130_fd_sc_hd__nand2_2 _28053_ (.A(_06304_),
    .B(_06298_),
    .Y(_06436_));
 sky130_fd_sc_hd__o21bai_2 _28054_ (.A1(_06431_),
    .A2(_06435_),
    .B1_N(_06436_),
    .Y(_06437_));
 sky130_fd_sc_hd__o21bai_2 _28055_ (.A1(_06433_),
    .A2(_06434_),
    .B1_N(_06430_),
    .Y(_06438_));
 sky130_fd_sc_hd__nand3_2 _28056_ (.A(_06425_),
    .B(_06430_),
    .C(_06428_),
    .Y(_06439_));
 sky130_fd_sc_hd__nand3_2 _28057_ (.A(_06438_),
    .B(_06439_),
    .C(_06436_),
    .Y(_06440_));
 sky130_fd_sc_hd__nand2_2 _28058_ (.A(_06437_),
    .B(_06440_),
    .Y(_06441_));
 sky130_fd_sc_hd__a21oi_2 _28059_ (.A1(_06310_),
    .A2(_06309_),
    .B1(_06308_),
    .Y(_06442_));
 sky130_fd_sc_hd__xor2_2 _28060_ (.A(_06441_),
    .B(_06442_),
    .X(_02632_));
 sky130_fd_sc_hd__nand2_2 _28061_ (.A(_06051_),
    .B(_05959_),
    .Y(_06443_));
 sky130_fd_sc_hd__buf_1 _28062_ (.A(_06357_),
    .X(_06444_));
 sky130_fd_sc_hd__nand2_2 _28063_ (.A(_05826_),
    .B(_06444_),
    .Y(_06445_));
 sky130_fd_sc_hd__nand2_2 _28064_ (.A(_06443_),
    .B(_06445_),
    .Y(_06446_));
 sky130_fd_sc_hd__nand3b_2 _28065_ (.A_N(_06443_),
    .B(_18851_),
    .C(_06358_),
    .Y(_06447_));
 sky130_fd_sc_hd__o2bb2ai_2 _28066_ (.A1_N(_06446_),
    .A2_N(_06447_),
    .B1(_06347_),
    .B2(_19234_),
    .Y(_06448_));
 sky130_fd_sc_hd__nor2_2 _28067_ (.A(_06339_),
    .B(_06340_),
    .Y(_06449_));
 sky130_fd_sc_hd__a21oi_2 _28068_ (.A1(_06341_),
    .A2(_06352_),
    .B1(_06449_),
    .Y(_06450_));
 sky130_vsdinv _28069_ (.A(_06450_),
    .Y(_06451_));
 sky130_fd_sc_hd__buf_1 _28070_ (.A(\pcpi_mul.rs1[14] ),
    .X(_06452_));
 sky130_fd_sc_hd__buf_1 _28071_ (.A(_06452_),
    .X(_06453_));
 sky130_fd_sc_hd__buf_1 _28072_ (.A(_06453_),
    .X(_06454_));
 sky130_fd_sc_hd__and2_2 _28073_ (.A(_05236_),
    .B(_06454_),
    .X(_06455_));
 sky130_fd_sc_hd__nand3_2 _28074_ (.A(_06447_),
    .B(_06455_),
    .C(_06446_),
    .Y(_06456_));
 sky130_fd_sc_hd__nand3_2 _28075_ (.A(_06448_),
    .B(_06451_),
    .C(_06456_),
    .Y(_06457_));
 sky130_vsdinv _28076_ (.A(_06457_),
    .Y(_06458_));
 sky130_fd_sc_hd__a21oi_2 _28077_ (.A1(_06448_),
    .A2(_06456_),
    .B1(_06451_),
    .Y(_06459_));
 sky130_fd_sc_hd__buf_1 _28078_ (.A(_05744_),
    .X(_06460_));
 sky130_fd_sc_hd__and2_2 _28079_ (.A(_06460_),
    .B(_06361_),
    .X(_06461_));
 sky130_fd_sc_hd__buf_1 _28080_ (.A(\pcpi_mul.rs1[12] ),
    .X(_06462_));
 sky130_fd_sc_hd__buf_1 _28081_ (.A(_06462_),
    .X(_06463_));
 sky130_fd_sc_hd__buf_1 _28082_ (.A(_06463_),
    .X(_06464_));
 sky130_fd_sc_hd__nand2_2 _28083_ (.A(_05550_),
    .B(_06464_),
    .Y(_06465_));
 sky130_fd_sc_hd__buf_1 _28084_ (.A(_19236_),
    .X(_06466_));
 sky130_fd_sc_hd__buf_1 _28085_ (.A(_06466_),
    .X(_06467_));
 sky130_fd_sc_hd__nand2_2 _28086_ (.A(_05429_),
    .B(_06467_),
    .Y(_06468_));
 sky130_fd_sc_hd__xnor2_2 _28087_ (.A(_06465_),
    .B(_06468_),
    .Y(_06469_));
 sky130_fd_sc_hd__xnor2_2 _28088_ (.A(_06461_),
    .B(_06469_),
    .Y(_06470_));
 sky130_fd_sc_hd__o21ba_2 _28089_ (.A1(_06458_),
    .A2(_06459_),
    .B1_N(_06470_),
    .X(_06471_));
 sky130_fd_sc_hd__nand3b_2 _28090_ (.A_N(_06459_),
    .B(_06470_),
    .C(_06457_),
    .Y(_06472_));
 sky130_fd_sc_hd__nand2_2 _28091_ (.A(_06371_),
    .B(_06356_),
    .Y(_06473_));
 sky130_fd_sc_hd__nand3b_2 _28092_ (.A_N(_06471_),
    .B(_06472_),
    .C(_06473_),
    .Y(_06474_));
 sky130_vsdinv _28093_ (.A(_06472_),
    .Y(_06475_));
 sky130_fd_sc_hd__o21bai_2 _28094_ (.A1(_06475_),
    .A2(_06471_),
    .B1_N(_06473_),
    .Y(_06476_));
 sky130_fd_sc_hd__buf_1 _28095_ (.A(_19241_),
    .X(_06477_));
 sky130_fd_sc_hd__buf_1 _28096_ (.A(_06477_),
    .X(_06478_));
 sky130_fd_sc_hd__buf_1 _28097_ (.A(_06478_),
    .X(_06479_));
 sky130_fd_sc_hd__nor3_2 _28098_ (.A(_18859_),
    .B(_19254_),
    .C(_06368_),
    .Y(_06480_));
 sky130_fd_sc_hd__a41oi_2 _28099_ (.A1(_18869_),
    .A2(_18875_),
    .A3(_06479_),
    .A4(_06361_),
    .B1(_06480_),
    .Y(_06481_));
 sky130_vsdinv _28100_ (.A(_06481_),
    .Y(_06482_));
 sky130_fd_sc_hd__nand3_2 _28101_ (.A(_06474_),
    .B(_06476_),
    .C(_06482_),
    .Y(_06483_));
 sky130_fd_sc_hd__a21o_2 _28102_ (.A1(_06474_),
    .A2(_06476_),
    .B1(_06482_),
    .X(_06484_));
 sky130_fd_sc_hd__nand2_2 _28103_ (.A(_05983_),
    .B(_05852_),
    .Y(_06485_));
 sky130_fd_sc_hd__buf_1 _28104_ (.A(_06180_),
    .X(_06486_));
 sky130_fd_sc_hd__nand2_2 _28105_ (.A(_06238_),
    .B(_06486_),
    .Y(_06487_));
 sky130_fd_sc_hd__nand2_2 _28106_ (.A(_06485_),
    .B(_06487_),
    .Y(_06488_));
 sky130_fd_sc_hd__nand3b_2 _28107_ (.A_N(_06485_),
    .B(_18835_),
    .C(_06317_),
    .Y(_06489_));
 sky130_fd_sc_hd__o2bb2ai_2 _28108_ (.A1_N(_06488_),
    .A2_N(_06489_),
    .B1(_06248_),
    .B2(_19263_),
    .Y(_06490_));
 sky130_fd_sc_hd__and2_2 _28109_ (.A(_05588_),
    .B(_05848_),
    .X(_06491_));
 sky130_fd_sc_hd__nand3_2 _28110_ (.A(_06489_),
    .B(_06491_),
    .C(_06488_),
    .Y(_06492_));
 sky130_fd_sc_hd__a21oi_2 _28111_ (.A1(_06400_),
    .A2(_06404_),
    .B1(_06401_),
    .Y(_06493_));
 sky130_vsdinv _28112_ (.A(_06493_),
    .Y(_06494_));
 sky130_fd_sc_hd__a21o_2 _28113_ (.A1(_06490_),
    .A2(_06492_),
    .B1(_06494_),
    .X(_06495_));
 sky130_fd_sc_hd__a21boi_2 _28114_ (.A1(_06318_),
    .A2(_06314_),
    .B1_N(_06315_),
    .Y(_06496_));
 sky130_vsdinv _28115_ (.A(_06496_),
    .Y(_06497_));
 sky130_fd_sc_hd__nand3_2 _28116_ (.A(_06490_),
    .B(_06494_),
    .C(_06492_),
    .Y(_06498_));
 sky130_fd_sc_hd__nand3_2 _28117_ (.A(_06495_),
    .B(_06497_),
    .C(_06498_),
    .Y(_06499_));
 sky130_fd_sc_hd__a21o_2 _28118_ (.A1(_06495_),
    .A2(_06498_),
    .B1(_06497_),
    .X(_06500_));
 sky130_fd_sc_hd__xnor2_2 _28119_ (.A(_06395_),
    .B(_06396_),
    .Y(_06501_));
 sky130_fd_sc_hd__o2bb2ai_2 _28120_ (.A1_N(_06499_),
    .A2_N(_06500_),
    .B1(_06501_),
    .B2(_06406_),
    .Y(_06502_));
 sky130_fd_sc_hd__nand3_2 _28121_ (.A(_06403_),
    .B(_06397_),
    .C(_06405_),
    .Y(_06503_));
 sky130_vsdinv _28122_ (.A(_06503_),
    .Y(_06504_));
 sky130_fd_sc_hd__nand3_2 _28123_ (.A(_06500_),
    .B(_06504_),
    .C(_06499_),
    .Y(_06505_));
 sky130_vsdinv _28124_ (.A(_06323_),
    .Y(_06506_));
 sky130_fd_sc_hd__a21oi_2 _28125_ (.A1(_06322_),
    .A2(_06325_),
    .B1(_06506_),
    .Y(_06507_));
 sky130_vsdinv _28126_ (.A(_06507_),
    .Y(_06508_));
 sky130_fd_sc_hd__a21oi_2 _28127_ (.A1(_06502_),
    .A2(_06505_),
    .B1(_06508_),
    .Y(_06509_));
 sky130_fd_sc_hd__nand3_2 _28128_ (.A(_06502_),
    .B(_06508_),
    .C(_06505_),
    .Y(_06510_));
 sky130_vsdinv _28129_ (.A(_06510_),
    .Y(_06511_));
 sky130_fd_sc_hd__a21oi_2 _28130_ (.A1(_06326_),
    .A2(_06327_),
    .B1(_06281_),
    .Y(_06512_));
 sky130_fd_sc_hd__o21ai_2 _28131_ (.A1(_06332_),
    .A2(_06512_),
    .B1(_06330_),
    .Y(_06513_));
 sky130_fd_sc_hd__o21bai_2 _28132_ (.A1(_06509_),
    .A2(_06511_),
    .B1_N(_06513_),
    .Y(_06514_));
 sky130_fd_sc_hd__a21o_2 _28133_ (.A1(_06502_),
    .A2(_06505_),
    .B1(_06508_),
    .X(_06515_));
 sky130_fd_sc_hd__nand3_2 _28134_ (.A(_06515_),
    .B(_06510_),
    .C(_06513_),
    .Y(_06516_));
 sky130_fd_sc_hd__a22oi_2 _28135_ (.A1(_06483_),
    .A2(_06484_),
    .B1(_06514_),
    .B2(_06516_),
    .Y(_06517_));
 sky130_fd_sc_hd__nand2_2 _28136_ (.A(_06484_),
    .B(_06483_),
    .Y(_06518_));
 sky130_fd_sc_hd__nand2_2 _28137_ (.A(_06514_),
    .B(_06516_),
    .Y(_06519_));
 sky130_fd_sc_hd__nor2_2 _28138_ (.A(_06518_),
    .B(_06519_),
    .Y(_06520_));
 sky130_vsdinv _28139_ (.A(_06338_),
    .Y(_06521_));
 sky130_fd_sc_hd__a21o_2 _28140_ (.A1(_06336_),
    .A2(_06382_),
    .B1(_06521_),
    .X(_06522_));
 sky130_fd_sc_hd__o21bai_2 _28141_ (.A1(_06517_),
    .A2(_06520_),
    .B1_N(_06522_),
    .Y(_06523_));
 sky130_fd_sc_hd__nand2_2 _28142_ (.A(_06519_),
    .B(_06518_),
    .Y(_06524_));
 sky130_fd_sc_hd__nand3b_2 _28143_ (.A_N(_06518_),
    .B(_06516_),
    .C(_06514_),
    .Y(_06525_));
 sky130_fd_sc_hd__nand3_2 _28144_ (.A(_06522_),
    .B(_06524_),
    .C(_06525_),
    .Y(_06526_));
 sky130_fd_sc_hd__nand2_2 _28145_ (.A(_06523_),
    .B(_06526_),
    .Y(_06527_));
 sky130_fd_sc_hd__and2_2 _28146_ (.A(_05896_),
    .B(_06232_),
    .X(_06528_));
 sky130_fd_sc_hd__nand2_2 _28147_ (.A(_06148_),
    .B(_05988_),
    .Y(_06529_));
 sky130_fd_sc_hd__nand2_2 _28148_ (.A(_18820_),
    .B(_05556_),
    .Y(_06530_));
 sky130_fd_sc_hd__xnor2_2 _28149_ (.A(_06529_),
    .B(_06530_),
    .Y(_06531_));
 sky130_fd_sc_hd__xor2_2 _28150_ (.A(_06528_),
    .B(_06531_),
    .X(_06532_));
 sky130_fd_sc_hd__buf_1 _28151_ (.A(\pcpi_mul.rs2[14] ),
    .X(_06533_));
 sky130_fd_sc_hd__buf_1 _28152_ (.A(_06533_),
    .X(_06534_));
 sky130_fd_sc_hd__buf_1 _28153_ (.A(_06534_),
    .X(_06535_));
 sky130_fd_sc_hd__buf_1 _28154_ (.A(\pcpi_mul.rs2[13] ),
    .X(_06536_));
 sky130_fd_sc_hd__buf_1 _28155_ (.A(_06536_),
    .X(_06537_));
 sky130_fd_sc_hd__buf_1 _28156_ (.A(_06537_),
    .X(_06538_));
 sky130_fd_sc_hd__a22oi_2 _28157_ (.A1(_06535_),
    .A2(_05567_),
    .B1(_06538_),
    .B2(_05425_),
    .Y(_06539_));
 sky130_fd_sc_hd__buf_1 _28158_ (.A(_18801_),
    .X(_06540_));
 sky130_fd_sc_hd__buf_1 _28159_ (.A(_06540_),
    .X(_06541_));
 sky130_fd_sc_hd__nand2_2 _28160_ (.A(_06541_),
    .B(_05402_),
    .Y(_06542_));
 sky130_fd_sc_hd__buf_1 _28161_ (.A(\pcpi_mul.rs2[14] ),
    .X(_06543_));
 sky130_fd_sc_hd__buf_1 _28162_ (.A(_06543_),
    .X(_06544_));
 sky130_fd_sc_hd__buf_1 _28163_ (.A(_06544_),
    .X(_06545_));
 sky130_fd_sc_hd__buf_1 _28164_ (.A(_05238_),
    .X(_06546_));
 sky130_fd_sc_hd__nand2_2 _28165_ (.A(_06545_),
    .B(_06546_),
    .Y(_06547_));
 sky130_fd_sc_hd__nor2_2 _28166_ (.A(_06542_),
    .B(_06547_),
    .Y(_06548_));
 sky130_vsdinv _28167_ (.A(_06548_),
    .Y(_06549_));
 sky130_fd_sc_hd__buf_1 _28168_ (.A(_18807_),
    .X(_06550_));
 sky130_fd_sc_hd__buf_1 _28169_ (.A(_06550_),
    .X(_06551_));
 sky130_fd_sc_hd__and2_2 _28170_ (.A(_06551_),
    .B(_05413_),
    .X(_06552_));
 sky130_fd_sc_hd__nand3b_2 _28171_ (.A_N(_06539_),
    .B(_06549_),
    .C(_06552_),
    .Y(_06553_));
 sky130_fd_sc_hd__o21bai_2 _28172_ (.A1(_06539_),
    .A2(_06548_),
    .B1_N(_06552_),
    .Y(_06554_));
 sky130_fd_sc_hd__nor2_2 _28173_ (.A(_06395_),
    .B(_06396_),
    .Y(_06555_));
 sky130_fd_sc_hd__a21oi_2 _28174_ (.A1(_06553_),
    .A2(_06554_),
    .B1(_06555_),
    .Y(_06556_));
 sky130_fd_sc_hd__nand3_2 _28175_ (.A(_06553_),
    .B(_06554_),
    .C(_06555_),
    .Y(_06557_));
 sky130_vsdinv _28176_ (.A(_06557_),
    .Y(_06558_));
 sky130_fd_sc_hd__nor2_2 _28177_ (.A(_06556_),
    .B(_06558_),
    .Y(_06559_));
 sky130_fd_sc_hd__xor2_2 _28178_ (.A(_06532_),
    .B(_06559_),
    .X(_06560_));
 sky130_fd_sc_hd__nand2_2 _28179_ (.A(_06527_),
    .B(_06560_),
    .Y(_06561_));
 sky130_fd_sc_hd__buf_1 _28180_ (.A(_06526_),
    .X(_06562_));
 sky130_fd_sc_hd__nand3b_2 _28181_ (.A_N(_06560_),
    .B(_06523_),
    .C(_06562_),
    .Y(_06563_));
 sky130_fd_sc_hd__a21oi_2 _28182_ (.A1(_06561_),
    .A2(_06563_),
    .B1(_06412_),
    .Y(_06564_));
 sky130_fd_sc_hd__nand3_2 _28183_ (.A(_06561_),
    .B(_06412_),
    .C(_06563_),
    .Y(_06565_));
 sky130_vsdinv _28184_ (.A(_06565_),
    .Y(_06566_));
 sky130_fd_sc_hd__nand2_2 _28185_ (.A(_06380_),
    .B(_06376_),
    .Y(_06567_));
 sky130_fd_sc_hd__xnor2_2 _28186_ (.A(_06567_),
    .B(_06391_),
    .Y(_06568_));
 sky130_vsdinv _28187_ (.A(_06568_),
    .Y(_06569_));
 sky130_fd_sc_hd__o21a_2 _28188_ (.A1(_06564_),
    .A2(_06566_),
    .B1(_06569_),
    .X(_06570_));
 sky130_fd_sc_hd__nor3b_2 _28189_ (.A(_06569_),
    .B(_06564_),
    .C_N(_06565_),
    .Y(_06571_));
 sky130_vsdinv _28190_ (.A(_06571_),
    .Y(_06572_));
 sky130_fd_sc_hd__o21ai_2 _28191_ (.A1(_06420_),
    .A2(_06421_),
    .B1(_06416_),
    .Y(_06573_));
 sky130_fd_sc_hd__nand3b_2 _28192_ (.A_N(_06570_),
    .B(_06572_),
    .C(_06573_),
    .Y(_06574_));
 sky130_fd_sc_hd__o21bai_2 _28193_ (.A1(_06571_),
    .A2(_06570_),
    .B1_N(_06573_),
    .Y(_06575_));
 sky130_fd_sc_hd__nor2_2 _28194_ (.A(_06417_),
    .B(_06263_),
    .Y(_06576_));
 sky130_fd_sc_hd__a21o_2 _28195_ (.A1(_06574_),
    .A2(_06575_),
    .B1(_06576_),
    .X(_06577_));
 sky130_fd_sc_hd__nand3_2 _28196_ (.A(_06574_),
    .B(_06576_),
    .C(_06575_),
    .Y(_06578_));
 sky130_fd_sc_hd__a21oi_2 _28197_ (.A1(_06425_),
    .A2(_06430_),
    .B1(_06434_),
    .Y(_06579_));
 sky130_fd_sc_hd__a21boi_2 _28198_ (.A1(_06577_),
    .A2(_06578_),
    .B1_N(_06579_),
    .Y(_06580_));
 sky130_fd_sc_hd__o211a_2 _28199_ (.A1(_06434_),
    .A2(_06435_),
    .B1(_06578_),
    .C1(_06577_),
    .X(_06581_));
 sky130_fd_sc_hd__nor2_2 _28200_ (.A(_06580_),
    .B(_06581_),
    .Y(_06582_));
 sky130_vsdinv _28201_ (.A(_06440_),
    .Y(_06583_));
 sky130_fd_sc_hd__o21bai_2 _28202_ (.A1(_06441_),
    .A2(_06442_),
    .B1_N(_06583_),
    .Y(_06584_));
 sky130_fd_sc_hd__xor2_2 _28203_ (.A(_06582_),
    .B(_06584_),
    .X(_02633_));
 sky130_fd_sc_hd__nand2_2 _28204_ (.A(_06578_),
    .B(_06574_),
    .Y(_06585_));
 sky130_fd_sc_hd__buf_1 _28205_ (.A(_05496_),
    .X(_06586_));
 sky130_fd_sc_hd__nand2_2 _28206_ (.A(_06586_),
    .B(_06064_),
    .Y(_06587_));
 sky130_fd_sc_hd__buf_1 _28207_ (.A(_06201_),
    .X(_06588_));
 sky130_fd_sc_hd__buf_1 _28208_ (.A(_06588_),
    .X(_06589_));
 sky130_fd_sc_hd__nand2_2 _28209_ (.A(_05732_),
    .B(_06589_),
    .Y(_06590_));
 sky130_fd_sc_hd__nand2_2 _28210_ (.A(_06587_),
    .B(_06590_),
    .Y(_06591_));
 sky130_fd_sc_hd__nor2_2 _28211_ (.A(_06587_),
    .B(_06590_),
    .Y(_06592_));
 sky130_vsdinv _28212_ (.A(_06592_),
    .Y(_06593_));
 sky130_fd_sc_hd__o2bb2ai_2 _28213_ (.A1_N(_06591_),
    .A2_N(_06593_),
    .B1(_18881_),
    .B2(_19228_),
    .Y(_06594_));
 sky130_fd_sc_hd__buf_1 _28214_ (.A(_19224_),
    .X(_06595_));
 sky130_fd_sc_hd__buf_1 _28215_ (.A(_06595_),
    .X(_06596_));
 sky130_fd_sc_hd__and2_2 _28216_ (.A(_06349_),
    .B(_06596_),
    .X(_06597_));
 sky130_fd_sc_hd__nand3b_2 _28217_ (.A_N(_06592_),
    .B(_06597_),
    .C(_06591_),
    .Y(_06598_));
 sky130_fd_sc_hd__nor2_2 _28218_ (.A(_06443_),
    .B(_06445_),
    .Y(_06599_));
 sky130_fd_sc_hd__a21oi_2 _28219_ (.A1(_06446_),
    .A2(_06455_),
    .B1(_06599_),
    .Y(_06600_));
 sky130_vsdinv _28220_ (.A(_06600_),
    .Y(_06601_));
 sky130_fd_sc_hd__a21o_2 _28221_ (.A1(_06594_),
    .A2(_06598_),
    .B1(_06601_),
    .X(_06602_));
 sky130_fd_sc_hd__nand3_2 _28222_ (.A(_06594_),
    .B(_06601_),
    .C(_06598_),
    .Y(_06603_));
 sky130_fd_sc_hd__and2_2 _28223_ (.A(_05460_),
    .B(_06479_),
    .X(_06604_));
 sky130_fd_sc_hd__nand2_2 _28224_ (.A(_05422_),
    .B(_06467_),
    .Y(_06605_));
 sky130_fd_sc_hd__buf_1 _28225_ (.A(_19230_),
    .X(_06606_));
 sky130_fd_sc_hd__buf_1 _28226_ (.A(_06606_),
    .X(_06607_));
 sky130_fd_sc_hd__buf_1 _28227_ (.A(_06607_),
    .X(_06608_));
 sky130_fd_sc_hd__nand2_2 _28228_ (.A(_06363_),
    .B(_06608_),
    .Y(_06609_));
 sky130_fd_sc_hd__xnor2_2 _28229_ (.A(_06605_),
    .B(_06609_),
    .Y(_06610_));
 sky130_fd_sc_hd__xnor2_2 _28230_ (.A(_06604_),
    .B(_06610_),
    .Y(_06611_));
 sky130_fd_sc_hd__a21o_2 _28231_ (.A1(_06602_),
    .A2(_06603_),
    .B1(_06611_),
    .X(_06612_));
 sky130_fd_sc_hd__nand3_2 _28232_ (.A(_06602_),
    .B(_06611_),
    .C(_06603_),
    .Y(_06613_));
 sky130_fd_sc_hd__nand2_2 _28233_ (.A(_06472_),
    .B(_06457_),
    .Y(_06614_));
 sky130_fd_sc_hd__a21o_2 _28234_ (.A1(_06612_),
    .A2(_06613_),
    .B1(_06614_),
    .X(_06615_));
 sky130_fd_sc_hd__buf_1 _28235_ (.A(_19237_),
    .X(_06616_));
 sky130_fd_sc_hd__buf_1 _28236_ (.A(_06616_),
    .X(_06617_));
 sky130_fd_sc_hd__nor3_2 _28237_ (.A(_05690_),
    .B(_19250_),
    .C(_06469_),
    .Y(_06618_));
 sky130_fd_sc_hd__a41oi_2 _28238_ (.A1(_18868_),
    .A2(_05408_),
    .A3(_06617_),
    .A4(_06479_),
    .B1(_06618_),
    .Y(_06619_));
 sky130_vsdinv _28239_ (.A(_06619_),
    .Y(_06620_));
 sky130_fd_sc_hd__nand3_2 _28240_ (.A(_06614_),
    .B(_06612_),
    .C(_06613_),
    .Y(_06621_));
 sky130_fd_sc_hd__nand3_2 _28241_ (.A(_06615_),
    .B(_06620_),
    .C(_06621_),
    .Y(_06622_));
 sky130_fd_sc_hd__a21o_2 _28242_ (.A1(_06615_),
    .A2(_06621_),
    .B1(_06620_),
    .X(_06623_));
 sky130_fd_sc_hd__nand2_2 _28243_ (.A(_05990_),
    .B(_05964_),
    .Y(_06624_));
 sky130_fd_sc_hd__nand2_2 _28244_ (.A(_06097_),
    .B(_05954_),
    .Y(_06625_));
 sky130_fd_sc_hd__nor2_2 _28245_ (.A(_06624_),
    .B(_06625_),
    .Y(_06626_));
 sky130_fd_sc_hd__and2_2 _28246_ (.A(_05779_),
    .B(_05951_),
    .X(_06627_));
 sky130_fd_sc_hd__nand2_2 _28247_ (.A(_06624_),
    .B(_06625_),
    .Y(_06628_));
 sky130_fd_sc_hd__nand3b_2 _28248_ (.A_N(_06626_),
    .B(_06627_),
    .C(_06628_),
    .Y(_06629_));
 sky130_fd_sc_hd__a22oi_2 _28249_ (.A1(_18830_),
    .A2(_06317_),
    .B1(_06238_),
    .B2(_05848_),
    .Y(_06630_));
 sky130_fd_sc_hd__o21bai_2 _28250_ (.A1(_06630_),
    .A2(_06626_),
    .B1_N(_06627_),
    .Y(_06631_));
 sky130_fd_sc_hd__nand2_2 _28251_ (.A(_06529_),
    .B(_06530_),
    .Y(_06632_));
 sky130_fd_sc_hd__nor2_2 _28252_ (.A(_06529_),
    .B(_06530_),
    .Y(_06633_));
 sky130_fd_sc_hd__a21oi_2 _28253_ (.A1(_06632_),
    .A2(_06528_),
    .B1(_06633_),
    .Y(_06634_));
 sky130_fd_sc_hd__a21bo_2 _28254_ (.A1(_06629_),
    .A2(_06631_),
    .B1_N(_06634_),
    .X(_06635_));
 sky130_fd_sc_hd__nand3b_2 _28255_ (.A_N(_06634_),
    .B(_06629_),
    .C(_06631_),
    .Y(_06636_));
 sky130_fd_sc_hd__nand2_2 _28256_ (.A(_06635_),
    .B(_06636_),
    .Y(_06637_));
 sky130_fd_sc_hd__a21boi_2 _28257_ (.A1(_06491_),
    .A2(_06488_),
    .B1_N(_06489_),
    .Y(_06638_));
 sky130_fd_sc_hd__nand2_2 _28258_ (.A(_06637_),
    .B(_06638_),
    .Y(_06639_));
 sky130_vsdinv _28259_ (.A(_06638_),
    .Y(_06640_));
 sky130_fd_sc_hd__nand3_2 _28260_ (.A(_06635_),
    .B(_06640_),
    .C(_06636_),
    .Y(_06641_));
 sky130_fd_sc_hd__o21bai_2 _28261_ (.A1(_06556_),
    .A2(_06532_),
    .B1_N(_06558_),
    .Y(_06642_));
 sky130_fd_sc_hd__a21o_2 _28262_ (.A1(_06639_),
    .A2(_06641_),
    .B1(_06642_),
    .X(_06643_));
 sky130_fd_sc_hd__nand3_2 _28263_ (.A(_06642_),
    .B(_06639_),
    .C(_06641_),
    .Y(_06644_));
 sky130_fd_sc_hd__nand2_2 _28264_ (.A(_06643_),
    .B(_06644_),
    .Y(_06645_));
 sky130_vsdinv _28265_ (.A(_06498_),
    .Y(_06646_));
 sky130_fd_sc_hd__a21oi_2 _28266_ (.A1(_06495_),
    .A2(_06497_),
    .B1(_06646_),
    .Y(_06647_));
 sky130_fd_sc_hd__nand2_2 _28267_ (.A(_06645_),
    .B(_06647_),
    .Y(_06648_));
 sky130_fd_sc_hd__nand3b_2 _28268_ (.A_N(_06647_),
    .B(_06643_),
    .C(_06644_),
    .Y(_06649_));
 sky130_fd_sc_hd__a21oi_2 _28269_ (.A1(_06500_),
    .A2(_06499_),
    .B1(_06504_),
    .Y(_06650_));
 sky130_fd_sc_hd__o21ai_2 _28270_ (.A1(_06507_),
    .A2(_06650_),
    .B1(_06505_),
    .Y(_06651_));
 sky130_fd_sc_hd__a21o_2 _28271_ (.A1(_06648_),
    .A2(_06649_),
    .B1(_06651_),
    .X(_06652_));
 sky130_fd_sc_hd__nand3_2 _28272_ (.A(_06648_),
    .B(_06651_),
    .C(_06649_),
    .Y(_06653_));
 sky130_fd_sc_hd__a22oi_2 _28273_ (.A1(_06622_),
    .A2(_06623_),
    .B1(_06652_),
    .B2(_06653_),
    .Y(_06654_));
 sky130_fd_sc_hd__nand2_2 _28274_ (.A(_06623_),
    .B(_06622_),
    .Y(_06655_));
 sky130_fd_sc_hd__nand2_2 _28275_ (.A(_06652_),
    .B(_06653_),
    .Y(_06656_));
 sky130_fd_sc_hd__nor2_2 _28276_ (.A(_06655_),
    .B(_06656_),
    .Y(_06657_));
 sky130_fd_sc_hd__a21oi_2 _28277_ (.A1(_06515_),
    .A2(_06510_),
    .B1(_06513_),
    .Y(_06658_));
 sky130_fd_sc_hd__o21ai_2 _28278_ (.A1(_06518_),
    .A2(_06658_),
    .B1(_06516_),
    .Y(_06659_));
 sky130_fd_sc_hd__o21bai_2 _28279_ (.A1(_06654_),
    .A2(_06657_),
    .B1_N(_06659_),
    .Y(_06660_));
 sky130_fd_sc_hd__nand3b_2 _28280_ (.A_N(_06655_),
    .B(_06652_),
    .C(_06653_),
    .Y(_06661_));
 sky130_fd_sc_hd__nand2_2 _28281_ (.A(_06656_),
    .B(_06655_),
    .Y(_06662_));
 sky130_fd_sc_hd__nand3_2 _28282_ (.A(_06659_),
    .B(_06661_),
    .C(_06662_),
    .Y(_06663_));
 sky130_fd_sc_hd__buf_1 _28283_ (.A(_06663_),
    .X(_06664_));
 sky130_fd_sc_hd__buf_1 _28284_ (.A(\pcpi_mul.rs2[15] ),
    .X(_06665_));
 sky130_fd_sc_hd__buf_1 _28285_ (.A(_06665_),
    .X(_06666_));
 sky130_fd_sc_hd__buf_1 _28286_ (.A(_06666_),
    .X(_06667_));
 sky130_fd_sc_hd__buf_1 _28287_ (.A(_06667_),
    .X(_06668_));
 sky130_fd_sc_hd__and2_2 _28288_ (.A(_06668_),
    .B(_05589_),
    .X(_06669_));
 sky130_fd_sc_hd__buf_1 _28289_ (.A(_18813_),
    .X(_06670_));
 sky130_fd_sc_hd__buf_1 _28290_ (.A(_06670_),
    .X(_06671_));
 sky130_fd_sc_hd__nand2_2 _28291_ (.A(_06671_),
    .B(_05733_),
    .Y(_06672_));
 sky130_fd_sc_hd__buf_1 _28292_ (.A(_06140_),
    .X(_06673_));
 sky130_fd_sc_hd__buf_1 _28293_ (.A(_06673_),
    .X(_06674_));
 sky130_fd_sc_hd__nand2_2 _28294_ (.A(_06674_),
    .B(_05746_),
    .Y(_06675_));
 sky130_fd_sc_hd__nand2_2 _28295_ (.A(_06672_),
    .B(_06675_),
    .Y(_06676_));
 sky130_fd_sc_hd__nor2_2 _28296_ (.A(_06672_),
    .B(_06675_),
    .Y(_06677_));
 sky130_vsdinv _28297_ (.A(_06677_),
    .Y(_06678_));
 sky130_fd_sc_hd__o2bb2ai_2 _28298_ (.A1_N(_06676_),
    .A2_N(_06678_),
    .B1(_18825_),
    .B2(_19275_),
    .Y(_06679_));
 sky130_fd_sc_hd__buf_1 _28299_ (.A(_18822_),
    .X(_06680_));
 sky130_fd_sc_hd__and2_2 _28300_ (.A(_06680_),
    .B(_19273_),
    .X(_06681_));
 sky130_fd_sc_hd__nand3b_2 _28301_ (.A_N(_06677_),
    .B(_06681_),
    .C(_06676_),
    .Y(_06682_));
 sky130_fd_sc_hd__nand2_2 _28302_ (.A(_06679_),
    .B(_06682_),
    .Y(_06683_));
 sky130_fd_sc_hd__nand2_2 _28303_ (.A(_06545_),
    .B(_06144_),
    .Y(_06684_));
 sky130_fd_sc_hd__nand2_2 _28304_ (.A(_06541_),
    .B(_05413_),
    .Y(_06685_));
 sky130_fd_sc_hd__nor2_2 _28305_ (.A(_06684_),
    .B(_06685_),
    .Y(_06686_));
 sky130_fd_sc_hd__nand2_2 _28306_ (.A(_06684_),
    .B(_06685_),
    .Y(_06687_));
 sky130_vsdinv _28307_ (.A(_06687_),
    .Y(_06688_));
 sky130_fd_sc_hd__and2_2 _28308_ (.A(_06551_),
    .B(_05552_),
    .X(_06689_));
 sky130_fd_sc_hd__o21bai_2 _28309_ (.A1(_06686_),
    .A2(_06688_),
    .B1_N(_06689_),
    .Y(_06690_));
 sky130_fd_sc_hd__nand3b_2 _28310_ (.A_N(_06686_),
    .B(_06689_),
    .C(_06687_),
    .Y(_06691_));
 sky130_fd_sc_hd__buf_1 _28311_ (.A(_18809_),
    .X(_06692_));
 sky130_fd_sc_hd__o31ai_2 _28312_ (.A1(_06692_),
    .A2(_19295_),
    .A3(_06539_),
    .B1(_06549_),
    .Y(_06693_));
 sky130_fd_sc_hd__a21oi_2 _28313_ (.A1(_06690_),
    .A2(_06691_),
    .B1(_06693_),
    .Y(_06694_));
 sky130_fd_sc_hd__nand3_2 _28314_ (.A(_06693_),
    .B(_06690_),
    .C(_06691_),
    .Y(_06695_));
 sky130_fd_sc_hd__nor3b_2 _28315_ (.A(_06683_),
    .B(_06694_),
    .C_N(_06695_),
    .Y(_06696_));
 sky130_vsdinv _28316_ (.A(_06695_),
    .Y(_06697_));
 sky130_fd_sc_hd__o21ai_2 _28317_ (.A1(_06694_),
    .A2(_06697_),
    .B1(_06683_),
    .Y(_06698_));
 sky130_fd_sc_hd__and2b_2 _28318_ (.A_N(_06696_),
    .B(_06698_),
    .X(_06699_));
 sky130_fd_sc_hd__xnor2_2 _28319_ (.A(_06669_),
    .B(_06699_),
    .Y(_06700_));
 sky130_fd_sc_hd__buf_1 _28320_ (.A(_06700_),
    .X(_06701_));
 sky130_fd_sc_hd__a21boi_2 _28321_ (.A1(_06660_),
    .A2(_06664_),
    .B1_N(_06701_),
    .Y(_06702_));
 sky130_fd_sc_hd__a21oi_2 _28322_ (.A1(_06661_),
    .A2(_06662_),
    .B1(_06659_),
    .Y(_06703_));
 sky130_fd_sc_hd__nor3b_2 _28323_ (.A(_06701_),
    .B(_06703_),
    .C_N(_06663_),
    .Y(_06704_));
 sky130_fd_sc_hd__o22ai_2 _28324_ (.A1(_06560_),
    .A2(_06527_),
    .B1(_06702_),
    .B2(_06704_),
    .Y(_06705_));
 sky130_fd_sc_hd__a21oi_2 _28325_ (.A1(_06524_),
    .A2(_06525_),
    .B1(_06522_),
    .Y(_06706_));
 sky130_fd_sc_hd__nor3b_2 _28326_ (.A(_06560_),
    .B(_06706_),
    .C_N(_06526_),
    .Y(_06707_));
 sky130_fd_sc_hd__nand2_2 _28327_ (.A(_06660_),
    .B(_06663_),
    .Y(_06708_));
 sky130_fd_sc_hd__nand2_2 _28328_ (.A(_06708_),
    .B(_06701_),
    .Y(_06709_));
 sky130_fd_sc_hd__nand3b_2 _28329_ (.A_N(_06700_),
    .B(_06660_),
    .C(_06664_),
    .Y(_06710_));
 sky130_fd_sc_hd__nand3_2 _28330_ (.A(_06707_),
    .B(_06709_),
    .C(_06710_),
    .Y(_06711_));
 sky130_fd_sc_hd__a21boi_2 _28331_ (.A1(_06482_),
    .A2(_06476_),
    .B1_N(_06474_),
    .Y(_06712_));
 sky130_fd_sc_hd__xor2_2 _28332_ (.A(_06712_),
    .B(_06562_),
    .X(_06713_));
 sky130_fd_sc_hd__a21oi_2 _28333_ (.A1(_06705_),
    .A2(_06711_),
    .B1(_06713_),
    .Y(_06714_));
 sky130_fd_sc_hd__nand3_2 _28334_ (.A(_06705_),
    .B(_06713_),
    .C(_06711_),
    .Y(_06715_));
 sky130_vsdinv _28335_ (.A(_06715_),
    .Y(_06716_));
 sky130_fd_sc_hd__o21ai_2 _28336_ (.A1(_06569_),
    .A2(_06564_),
    .B1(_06565_),
    .Y(_06717_));
 sky130_fd_sc_hd__o21bai_2 _28337_ (.A1(_06714_),
    .A2(_06716_),
    .B1_N(_06717_),
    .Y(_06718_));
 sky130_fd_sc_hd__a21o_2 _28338_ (.A1(_06705_),
    .A2(_06711_),
    .B1(_06713_),
    .X(_06719_));
 sky130_fd_sc_hd__nand3_2 _28339_ (.A(_06719_),
    .B(_06717_),
    .C(_06715_),
    .Y(_06720_));
 sky130_fd_sc_hd__o2111a_2 _28340_ (.A1(_06386_),
    .A2(_06265_),
    .B1(_06384_),
    .C1(_06567_),
    .D1(_06390_),
    .X(_06721_));
 sky130_fd_sc_hd__a21oi_2 _28341_ (.A1(_06718_),
    .A2(_06720_),
    .B1(_06721_),
    .Y(_06722_));
 sky130_fd_sc_hd__and3_2 _28342_ (.A(_06718_),
    .B(_06721_),
    .C(_06720_),
    .X(_06723_));
 sky130_fd_sc_hd__nor2_2 _28343_ (.A(_06722_),
    .B(_06723_),
    .Y(_06724_));
 sky130_fd_sc_hd__xnor2_2 _28344_ (.A(_06585_),
    .B(_06724_),
    .Y(_06725_));
 sky130_fd_sc_hd__a21oi_2 _28345_ (.A1(_06584_),
    .A2(_06582_),
    .B1(_06581_),
    .Y(_06726_));
 sky130_fd_sc_hd__xor2_2 _28346_ (.A(_06725_),
    .B(_06726_),
    .X(_02634_));
 sky130_fd_sc_hd__nand2_2 _28347_ (.A(_05492_),
    .B(_06589_),
    .Y(_06727_));
 sky130_fd_sc_hd__buf_1 _28348_ (.A(_06462_),
    .X(_06728_));
 sky130_fd_sc_hd__buf_1 _28349_ (.A(_06728_),
    .X(_06729_));
 sky130_fd_sc_hd__nand2_2 _28350_ (.A(_05652_),
    .B(_06729_),
    .Y(_06730_));
 sky130_fd_sc_hd__nor2_2 _28351_ (.A(_06727_),
    .B(_06730_),
    .Y(_06731_));
 sky130_fd_sc_hd__buf_1 _28352_ (.A(_18877_),
    .X(_06732_));
 sky130_fd_sc_hd__buf_1 _28353_ (.A(\pcpi_mul.rs1[16] ),
    .X(_06733_));
 sky130_fd_sc_hd__buf_1 _28354_ (.A(_06733_),
    .X(_06734_));
 sky130_fd_sc_hd__buf_1 _28355_ (.A(_06734_),
    .X(_06735_));
 sky130_fd_sc_hd__and2_2 _28356_ (.A(_06732_),
    .B(_06735_),
    .X(_06736_));
 sky130_fd_sc_hd__nand2_2 _28357_ (.A(_06727_),
    .B(_06730_),
    .Y(_06737_));
 sky130_fd_sc_hd__nand3b_2 _28358_ (.A_N(_06731_),
    .B(_06736_),
    .C(_06737_),
    .Y(_06738_));
 sky130_fd_sc_hd__a22oi_2 _28359_ (.A1(_05566_),
    .A2(_06361_),
    .B1(_05940_),
    .B2(_06366_),
    .Y(_06739_));
 sky130_fd_sc_hd__o21bai_2 _28360_ (.A1(_06739_),
    .A2(_06731_),
    .B1_N(_06736_),
    .Y(_06740_));
 sky130_fd_sc_hd__a21oi_2 _28361_ (.A1(_06591_),
    .A2(_06597_),
    .B1(_06592_),
    .Y(_06741_));
 sky130_fd_sc_hd__a21boi_2 _28362_ (.A1(_06738_),
    .A2(_06740_),
    .B1_N(_06741_),
    .Y(_06742_));
 sky130_fd_sc_hd__nand2_2 _28363_ (.A(_05550_),
    .B(_06454_),
    .Y(_06743_));
 sky130_fd_sc_hd__buf_1 _28364_ (.A(\pcpi_mul.rs1[15] ),
    .X(_06744_));
 sky130_fd_sc_hd__buf_1 _28365_ (.A(_06744_),
    .X(_06745_));
 sky130_fd_sc_hd__buf_1 _28366_ (.A(_06745_),
    .X(_06746_));
 sky130_fd_sc_hd__nand2_2 _28367_ (.A(_05429_),
    .B(_06746_),
    .Y(_06747_));
 sky130_fd_sc_hd__xor2_2 _28368_ (.A(_06743_),
    .B(_06747_),
    .X(_06748_));
 sky130_fd_sc_hd__and2_2 _28369_ (.A(_05460_),
    .B(_06617_),
    .X(_06749_));
 sky130_fd_sc_hd__nand2_2 _28370_ (.A(_06748_),
    .B(_06749_),
    .Y(_06750_));
 sky130_fd_sc_hd__xnor2_2 _28371_ (.A(_06743_),
    .B(_06747_),
    .Y(_06751_));
 sky130_fd_sc_hd__o21ai_2 _28372_ (.A1(_18858_),
    .A2(_19239_),
    .B1(_06751_),
    .Y(_06752_));
 sky130_fd_sc_hd__nand2_2 _28373_ (.A(_06750_),
    .B(_06752_),
    .Y(_06753_));
 sky130_fd_sc_hd__nand3b_2 _28374_ (.A_N(_06741_),
    .B(_06738_),
    .C(_06740_),
    .Y(_06754_));
 sky130_vsdinv _28375_ (.A(_06754_),
    .Y(_06755_));
 sky130_fd_sc_hd__nor3_2 _28376_ (.A(_06742_),
    .B(_06753_),
    .C(_06755_),
    .Y(_06756_));
 sky130_fd_sc_hd__o21a_2 _28377_ (.A1(_06742_),
    .A2(_06755_),
    .B1(_06753_),
    .X(_06757_));
 sky130_fd_sc_hd__o211ai_2 _28378_ (.A1(_06756_),
    .A2(_06757_),
    .B1(_06603_),
    .C1(_06613_),
    .Y(_06758_));
 sky130_fd_sc_hd__nand2_2 _28379_ (.A(_06613_),
    .B(_06603_),
    .Y(_06759_));
 sky130_vsdinv _28380_ (.A(_06756_),
    .Y(_06760_));
 sky130_fd_sc_hd__nand3b_2 _28381_ (.A_N(_06757_),
    .B(_06759_),
    .C(_06760_),
    .Y(_06761_));
 sky130_fd_sc_hd__nor3_2 _28382_ (.A(_18859_),
    .B(_19244_),
    .C(_06610_),
    .Y(_06762_));
 sky130_fd_sc_hd__a41oi_2 _28383_ (.A1(_18869_),
    .A2(_05408_),
    .A3(_06608_),
    .A4(_06617_),
    .B1(_06762_),
    .Y(_06763_));
 sky130_vsdinv _28384_ (.A(_06763_),
    .Y(_06764_));
 sky130_fd_sc_hd__nand3_2 _28385_ (.A(_06758_),
    .B(_06761_),
    .C(_06764_),
    .Y(_06765_));
 sky130_fd_sc_hd__a21o_2 _28386_ (.A1(_06758_),
    .A2(_06761_),
    .B1(_06764_),
    .X(_06766_));
 sky130_fd_sc_hd__a22oi_2 _28387_ (.A1(_06311_),
    .A2(_05842_),
    .B1(_05769_),
    .B2(_06344_),
    .Y(_06767_));
 sky130_fd_sc_hd__nand2_2 _28388_ (.A(_05982_),
    .B(_06181_),
    .Y(_06768_));
 sky130_fd_sc_hd__nand2_2 _28389_ (.A(_06237_),
    .B(_05959_),
    .Y(_06769_));
 sky130_fd_sc_hd__nor2_2 _28390_ (.A(_06768_),
    .B(_06769_),
    .Y(_06770_));
 sky130_fd_sc_hd__buf_1 _28391_ (.A(_06100_),
    .X(_06771_));
 sky130_fd_sc_hd__and2_2 _28392_ (.A(_06771_),
    .B(_06069_),
    .X(_06772_));
 sky130_fd_sc_hd__o21bai_2 _28393_ (.A1(_06767_),
    .A2(_06770_),
    .B1_N(_06772_),
    .Y(_06773_));
 sky130_fd_sc_hd__nand3b_2 _28394_ (.A_N(_06768_),
    .B(_06231_),
    .C(_06344_),
    .Y(_06774_));
 sky130_fd_sc_hd__nand2_2 _28395_ (.A(_06768_),
    .B(_06769_),
    .Y(_06775_));
 sky130_fd_sc_hd__nand3_2 _28396_ (.A(_06774_),
    .B(_06772_),
    .C(_06775_),
    .Y(_06776_));
 sky130_fd_sc_hd__nand2_2 _28397_ (.A(_06773_),
    .B(_06776_),
    .Y(_06777_));
 sky130_fd_sc_hd__a21oi_2 _28398_ (.A1(_06676_),
    .A2(_06681_),
    .B1(_06677_),
    .Y(_06778_));
 sky130_fd_sc_hd__nand2_2 _28399_ (.A(_06777_),
    .B(_06778_),
    .Y(_06779_));
 sky130_fd_sc_hd__nand3b_2 _28400_ (.A_N(_06778_),
    .B(_06776_),
    .C(_06773_),
    .Y(_06780_));
 sky130_fd_sc_hd__nand2_2 _28401_ (.A(_06779_),
    .B(_06780_),
    .Y(_06781_));
 sky130_fd_sc_hd__a21oi_2 _28402_ (.A1(_06628_),
    .A2(_06627_),
    .B1(_06626_),
    .Y(_06782_));
 sky130_fd_sc_hd__nand2_2 _28403_ (.A(_06781_),
    .B(_06782_),
    .Y(_06783_));
 sky130_vsdinv _28404_ (.A(_06782_),
    .Y(_06784_));
 sky130_fd_sc_hd__nand3_2 _28405_ (.A(_06779_),
    .B(_06784_),
    .C(_06780_),
    .Y(_06785_));
 sky130_fd_sc_hd__o21ai_2 _28406_ (.A1(_06683_),
    .A2(_06694_),
    .B1(_06695_),
    .Y(_06786_));
 sky130_fd_sc_hd__a21oi_2 _28407_ (.A1(_06783_),
    .A2(_06785_),
    .B1(_06786_),
    .Y(_06787_));
 sky130_fd_sc_hd__nand3_2 _28408_ (.A(_06786_),
    .B(_06783_),
    .C(_06785_),
    .Y(_06788_));
 sky130_vsdinv _28409_ (.A(_06788_),
    .Y(_06789_));
 sky130_vsdinv _28410_ (.A(_06636_),
    .Y(_06790_));
 sky130_fd_sc_hd__a21oi_2 _28411_ (.A1(_06635_),
    .A2(_06640_),
    .B1(_06790_),
    .Y(_06791_));
 sky130_vsdinv _28412_ (.A(_06791_),
    .Y(_06792_));
 sky130_fd_sc_hd__o21bai_2 _28413_ (.A1(_06787_),
    .A2(_06789_),
    .B1_N(_06792_),
    .Y(_06793_));
 sky130_fd_sc_hd__a21o_2 _28414_ (.A1(_06783_),
    .A2(_06785_),
    .B1(_06786_),
    .X(_06794_));
 sky130_fd_sc_hd__nand3b_2 _28415_ (.A_N(_06791_),
    .B(_06794_),
    .C(_06788_),
    .Y(_06795_));
 sky130_fd_sc_hd__a21oi_2 _28416_ (.A1(_06639_),
    .A2(_06641_),
    .B1(_06642_),
    .Y(_06796_));
 sky130_fd_sc_hd__o21ai_2 _28417_ (.A1(_06647_),
    .A2(_06796_),
    .B1(_06644_),
    .Y(_06797_));
 sky130_fd_sc_hd__a21o_2 _28418_ (.A1(_06793_),
    .A2(_06795_),
    .B1(_06797_),
    .X(_06798_));
 sky130_fd_sc_hd__nand3_2 _28419_ (.A(_06793_),
    .B(_06797_),
    .C(_06795_),
    .Y(_06799_));
 sky130_fd_sc_hd__a22oi_2 _28420_ (.A1(_06765_),
    .A2(_06766_),
    .B1(_06798_),
    .B2(_06799_),
    .Y(_06800_));
 sky130_fd_sc_hd__nand2_2 _28421_ (.A(_06766_),
    .B(_06765_),
    .Y(_06801_));
 sky130_fd_sc_hd__nand2_2 _28422_ (.A(_06798_),
    .B(_06799_),
    .Y(_06802_));
 sky130_fd_sc_hd__nor2_2 _28423_ (.A(_06801_),
    .B(_06802_),
    .Y(_06803_));
 sky130_fd_sc_hd__a21oi_2 _28424_ (.A1(_06648_),
    .A2(_06649_),
    .B1(_06651_),
    .Y(_06804_));
 sky130_fd_sc_hd__o21ai_2 _28425_ (.A1(_06804_),
    .A2(_06655_),
    .B1(_06653_),
    .Y(_06805_));
 sky130_fd_sc_hd__o21bai_2 _28426_ (.A1(_06800_),
    .A2(_06803_),
    .B1_N(_06805_),
    .Y(_06806_));
 sky130_fd_sc_hd__nand3b_2 _28427_ (.A_N(_06801_),
    .B(_06799_),
    .C(_06798_),
    .Y(_06807_));
 sky130_fd_sc_hd__nand3b_2 _28428_ (.A_N(_06800_),
    .B(_06805_),
    .C(_06807_),
    .Y(_06808_));
 sky130_fd_sc_hd__and3b_2 _28429_ (.A_N(_06696_),
    .B(_06698_),
    .C(_06669_),
    .X(_06809_));
 sky130_fd_sc_hd__buf_1 _28430_ (.A(\pcpi_mul.rs2[11] ),
    .X(_06810_));
 sky130_fd_sc_hd__buf_1 _28431_ (.A(_06810_),
    .X(_06811_));
 sky130_fd_sc_hd__buf_1 _28432_ (.A(_06673_),
    .X(_06812_));
 sky130_fd_sc_hd__a22oi_2 _28433_ (.A1(_06811_),
    .A2(_06102_),
    .B1(_06812_),
    .B2(_06052_),
    .Y(_06813_));
 sky130_fd_sc_hd__and4_2 _28434_ (.A(_18815_),
    .B(_18820_),
    .C(_05941_),
    .D(_06232_),
    .X(_06814_));
 sky130_fd_sc_hd__buf_1 _28435_ (.A(\pcpi_mul.rs2[9] ),
    .X(_06815_));
 sky130_fd_sc_hd__buf_1 _28436_ (.A(_06815_),
    .X(_06816_));
 sky130_fd_sc_hd__nand2_2 _28437_ (.A(_06816_),
    .B(_06486_),
    .Y(_06817_));
 sky130_vsdinv _28438_ (.A(_06817_),
    .Y(_06818_));
 sky130_fd_sc_hd__o21bai_2 _28439_ (.A1(_06813_),
    .A2(_06814_),
    .B1_N(_06818_),
    .Y(_06819_));
 sky130_fd_sc_hd__buf_1 _28440_ (.A(_05668_),
    .X(_06820_));
 sky130_fd_sc_hd__nand2_2 _28441_ (.A(_18814_),
    .B(_06820_),
    .Y(_06821_));
 sky130_fd_sc_hd__nand3b_2 _28442_ (.A_N(_06821_),
    .B(_06142_),
    .C(_05852_),
    .Y(_06822_));
 sky130_fd_sc_hd__nand3b_2 _28443_ (.A_N(_06813_),
    .B(_06822_),
    .C(_06818_),
    .Y(_06823_));
 sky130_fd_sc_hd__nand2_2 _28444_ (.A(_06819_),
    .B(_06823_),
    .Y(_06824_));
 sky130_fd_sc_hd__nand2_2 _28445_ (.A(_06534_),
    .B(_05636_),
    .Y(_06825_));
 sky130_fd_sc_hd__buf_1 _28446_ (.A(_05443_),
    .X(_06826_));
 sky130_fd_sc_hd__buf_1 _28447_ (.A(_06826_),
    .X(_06827_));
 sky130_fd_sc_hd__nand2_2 _28448_ (.A(_06537_),
    .B(_06827_),
    .Y(_06828_));
 sky130_fd_sc_hd__nor2_2 _28449_ (.A(_06825_),
    .B(_06828_),
    .Y(_06829_));
 sky130_fd_sc_hd__and2_2 _28450_ (.A(_06550_),
    .B(_05470_),
    .X(_06830_));
 sky130_fd_sc_hd__nand2_2 _28451_ (.A(_06825_),
    .B(_06828_),
    .Y(_06831_));
 sky130_fd_sc_hd__nand3b_2 _28452_ (.A_N(_06829_),
    .B(_06830_),
    .C(_06831_),
    .Y(_06832_));
 sky130_fd_sc_hd__a22oi_2 _28453_ (.A1(_18799_),
    .A2(_05432_),
    .B1(_06394_),
    .B2(_05446_),
    .Y(_06833_));
 sky130_fd_sc_hd__o21bai_2 _28454_ (.A1(_06833_),
    .A2(_06829_),
    .B1_N(_06830_),
    .Y(_06834_));
 sky130_fd_sc_hd__a21oi_2 _28455_ (.A1(_06687_),
    .A2(_06689_),
    .B1(_06686_),
    .Y(_06835_));
 sky130_fd_sc_hd__a21boi_2 _28456_ (.A1(_06832_),
    .A2(_06834_),
    .B1_N(_06835_),
    .Y(_06836_));
 sky130_fd_sc_hd__nand3b_2 _28457_ (.A_N(_06835_),
    .B(_06832_),
    .C(_06834_),
    .Y(_06837_));
 sky130_fd_sc_hd__nor3b_2 _28458_ (.A(_06824_),
    .B(_06836_),
    .C_N(_06837_),
    .Y(_06838_));
 sky130_vsdinv _28459_ (.A(_06838_),
    .Y(_06839_));
 sky130_vsdinv _28460_ (.A(_06837_),
    .Y(_06840_));
 sky130_fd_sc_hd__o21ai_2 _28461_ (.A1(_06836_),
    .A2(_06840_),
    .B1(_06824_),
    .Y(_06841_));
 sky130_fd_sc_hd__nand2_2 _28462_ (.A(_18787_),
    .B(_05466_),
    .Y(_06842_));
 sky130_fd_sc_hd__nand2_2 _28463_ (.A(_06667_),
    .B(_05403_),
    .Y(_06843_));
 sky130_fd_sc_hd__xor2_2 _28464_ (.A(_06842_),
    .B(_06843_),
    .X(_06844_));
 sky130_fd_sc_hd__a21oi_2 _28465_ (.A1(_06839_),
    .A2(_06841_),
    .B1(_06844_),
    .Y(_06845_));
 sky130_fd_sc_hd__nand3b_2 _28466_ (.A_N(_06838_),
    .B(_06844_),
    .C(_06841_),
    .Y(_06846_));
 sky130_fd_sc_hd__or2b_2 _28467_ (.A(_06845_),
    .B_N(_06846_),
    .X(_06847_));
 sky130_fd_sc_hd__xnor2_2 _28468_ (.A(_06809_),
    .B(_06847_),
    .Y(_06848_));
 sky130_fd_sc_hd__a21oi_2 _28469_ (.A1(_06806_),
    .A2(_06808_),
    .B1(_06848_),
    .Y(_06849_));
 sky130_fd_sc_hd__nand3_2 _28470_ (.A(_06806_),
    .B(_06848_),
    .C(_06808_),
    .Y(_06850_));
 sky130_vsdinv _28471_ (.A(_06850_),
    .Y(_06851_));
 sky130_fd_sc_hd__o22ai_2 _28472_ (.A1(_06701_),
    .A2(_06708_),
    .B1(_06849_),
    .B2(_06851_),
    .Y(_06852_));
 sky130_fd_sc_hd__buf_1 _28473_ (.A(_06808_),
    .X(_06853_));
 sky130_fd_sc_hd__a21o_2 _28474_ (.A1(_06806_),
    .A2(_06853_),
    .B1(_06848_),
    .X(_06854_));
 sky130_fd_sc_hd__nand3_2 _28475_ (.A(_06704_),
    .B(_06854_),
    .C(_06850_),
    .Y(_06855_));
 sky130_fd_sc_hd__a21boi_2 _28476_ (.A1(_06615_),
    .A2(_06620_),
    .B1_N(_06621_),
    .Y(_06856_));
 sky130_fd_sc_hd__xor2_2 _28477_ (.A(_06856_),
    .B(_06664_),
    .X(_06857_));
 sky130_fd_sc_hd__a21oi_2 _28478_ (.A1(_06852_),
    .A2(_06855_),
    .B1(_06857_),
    .Y(_06858_));
 sky130_fd_sc_hd__nand3_2 _28479_ (.A(_06852_),
    .B(_06855_),
    .C(_06857_),
    .Y(_06859_));
 sky130_vsdinv _28480_ (.A(_06713_),
    .Y(_06860_));
 sky130_fd_sc_hd__a21boi_2 _28481_ (.A1(_06709_),
    .A2(_06710_),
    .B1_N(_06563_),
    .Y(_06861_));
 sky130_fd_sc_hd__o21ai_2 _28482_ (.A1(_06860_),
    .A2(_06861_),
    .B1(_06711_),
    .Y(_06862_));
 sky130_fd_sc_hd__nand3b_2 _28483_ (.A_N(_06858_),
    .B(_06859_),
    .C(_06862_),
    .Y(_06863_));
 sky130_vsdinv _28484_ (.A(_06859_),
    .Y(_06864_));
 sky130_fd_sc_hd__o21bai_2 _28485_ (.A1(_06858_),
    .A2(_06864_),
    .B1_N(_06862_),
    .Y(_06865_));
 sky130_fd_sc_hd__o2bb2ai_2 _28486_ (.A1_N(_06863_),
    .A2_N(_06865_),
    .B1(_06562_),
    .B2(_06712_),
    .Y(_06866_));
 sky130_fd_sc_hd__nor2_2 _28487_ (.A(_06712_),
    .B(_06562_),
    .Y(_06867_));
 sky130_fd_sc_hd__nand3_2 _28488_ (.A(_06865_),
    .B(_06863_),
    .C(_06867_),
    .Y(_06868_));
 sky130_fd_sc_hd__nand2_2 _28489_ (.A(_06866_),
    .B(_06868_),
    .Y(_06869_));
 sky130_fd_sc_hd__a21boi_2 _28490_ (.A1(_06718_),
    .A2(_06721_),
    .B1_N(_06720_),
    .Y(_06870_));
 sky130_fd_sc_hd__nand2_2 _28491_ (.A(_06869_),
    .B(_06870_),
    .Y(_06871_));
 sky130_fd_sc_hd__a21bo_2 _28492_ (.A1(_06718_),
    .A2(_06721_),
    .B1_N(_06720_),
    .X(_06872_));
 sky130_fd_sc_hd__nand3_2 _28493_ (.A(_06872_),
    .B(_06868_),
    .C(_06866_),
    .Y(_06873_));
 sky130_fd_sc_hd__and2_2 _28494_ (.A(_06871_),
    .B(_06873_),
    .X(_06874_));
 sky130_fd_sc_hd__nor2_2 _28495_ (.A(_06585_),
    .B(_06724_),
    .Y(_06875_));
 sky130_fd_sc_hd__a211oi_2 _28496_ (.A1(_06578_),
    .A2(_06574_),
    .B1(_06722_),
    .C1(_06723_),
    .Y(_06876_));
 sky130_fd_sc_hd__o21bai_2 _28497_ (.A1(_06875_),
    .A2(_06726_),
    .B1_N(_06876_),
    .Y(_06877_));
 sky130_fd_sc_hd__buf_1 _28498_ (.A(_06877_),
    .X(_06878_));
 sky130_fd_sc_hd__xor2_2 _28499_ (.A(_06874_),
    .B(_06878_),
    .X(_02635_));
 sky130_fd_sc_hd__a22oi_2 _28500_ (.A1(_05870_),
    .A2(_06061_),
    .B1(_06237_),
    .B2(_06064_),
    .Y(_06879_));
 sky130_fd_sc_hd__buf_1 _28501_ (.A(\pcpi_mul.rs2[8] ),
    .X(_06880_));
 sky130_fd_sc_hd__buf_1 _28502_ (.A(_06880_),
    .X(_06881_));
 sky130_fd_sc_hd__nand2_2 _28503_ (.A(_06881_),
    .B(_06060_),
    .Y(_06882_));
 sky130_fd_sc_hd__buf_1 _28504_ (.A(_05934_),
    .X(_06883_));
 sky130_fd_sc_hd__nand2_2 _28505_ (.A(_06226_),
    .B(_06883_),
    .Y(_06884_));
 sky130_fd_sc_hd__nor2_2 _28506_ (.A(_06882_),
    .B(_06884_),
    .Y(_06885_));
 sky130_fd_sc_hd__buf_1 _28507_ (.A(_06046_),
    .X(_06886_));
 sky130_fd_sc_hd__and2_2 _28508_ (.A(_05778_),
    .B(_06886_),
    .X(_06887_));
 sky130_fd_sc_hd__o21bai_2 _28509_ (.A1(_06879_),
    .A2(_06885_),
    .B1_N(_06887_),
    .Y(_06888_));
 sky130_fd_sc_hd__buf_1 _28510_ (.A(_06095_),
    .X(_06889_));
 sky130_fd_sc_hd__buf_1 _28511_ (.A(_06889_),
    .X(_06890_));
 sky130_fd_sc_hd__nand3b_2 _28512_ (.A_N(_06882_),
    .B(_06890_),
    .C(_06444_),
    .Y(_06891_));
 sky130_fd_sc_hd__nand2_2 _28513_ (.A(_06882_),
    .B(_06884_),
    .Y(_06892_));
 sky130_fd_sc_hd__nand3_2 _28514_ (.A(_06891_),
    .B(_06887_),
    .C(_06892_),
    .Y(_06893_));
 sky130_fd_sc_hd__nand2_2 _28515_ (.A(_06888_),
    .B(_06893_),
    .Y(_06894_));
 sky130_fd_sc_hd__o21ai_2 _28516_ (.A1(_06817_),
    .A2(_06813_),
    .B1(_06822_),
    .Y(_06895_));
 sky130_vsdinv _28517_ (.A(_06895_),
    .Y(_06896_));
 sky130_fd_sc_hd__nand2_2 _28518_ (.A(_06894_),
    .B(_06896_),
    .Y(_06897_));
 sky130_fd_sc_hd__nand3_2 _28519_ (.A(_06888_),
    .B(_06895_),
    .C(_06893_),
    .Y(_06898_));
 sky130_fd_sc_hd__a21oi_2 _28520_ (.A1(_06775_),
    .A2(_06772_),
    .B1(_06770_),
    .Y(_06899_));
 sky130_vsdinv _28521_ (.A(_06899_),
    .Y(_06900_));
 sky130_fd_sc_hd__a21oi_2 _28522_ (.A1(_06897_),
    .A2(_06898_),
    .B1(_06900_),
    .Y(_06901_));
 sky130_fd_sc_hd__a21oi_2 _28523_ (.A1(_06888_),
    .A2(_06893_),
    .B1(_06895_),
    .Y(_06902_));
 sky130_vsdinv _28524_ (.A(_06898_),
    .Y(_06903_));
 sky130_fd_sc_hd__nor3_2 _28525_ (.A(_06899_),
    .B(_06902_),
    .C(_06903_),
    .Y(_06904_));
 sky130_fd_sc_hd__o21ai_2 _28526_ (.A1(_06824_),
    .A2(_06836_),
    .B1(_06837_),
    .Y(_06905_));
 sky130_fd_sc_hd__o21bai_2 _28527_ (.A1(_06901_),
    .A2(_06904_),
    .B1_N(_06905_),
    .Y(_06906_));
 sky130_fd_sc_hd__o21bai_2 _28528_ (.A1(_06902_),
    .A2(_06903_),
    .B1_N(_06900_),
    .Y(_06907_));
 sky130_fd_sc_hd__nand3_2 _28529_ (.A(_06897_),
    .B(_06900_),
    .C(_06898_),
    .Y(_06908_));
 sky130_fd_sc_hd__nand3_2 _28530_ (.A(_06907_),
    .B(_06905_),
    .C(_06908_),
    .Y(_06909_));
 sky130_fd_sc_hd__buf_1 _28531_ (.A(_06909_),
    .X(_06910_));
 sky130_fd_sc_hd__a21boi_2 _28532_ (.A1(_06779_),
    .A2(_06784_),
    .B1_N(_06780_),
    .Y(_06911_));
 sky130_vsdinv _28533_ (.A(_06911_),
    .Y(_06912_));
 sky130_fd_sc_hd__a21oi_2 _28534_ (.A1(_06906_),
    .A2(_06910_),
    .B1(_06912_),
    .Y(_06913_));
 sky130_vsdinv _28535_ (.A(_06780_),
    .Y(_06914_));
 sky130_vsdinv _28536_ (.A(_06785_),
    .Y(_06915_));
 sky130_fd_sc_hd__o211a_2 _28537_ (.A1(_06914_),
    .A2(_06915_),
    .B1(_06910_),
    .C1(_06906_),
    .X(_06916_));
 sky130_fd_sc_hd__o21ai_2 _28538_ (.A1(_06791_),
    .A2(_06787_),
    .B1(_06788_),
    .Y(_06917_));
 sky130_fd_sc_hd__o21bai_2 _28539_ (.A1(_06913_),
    .A2(_06916_),
    .B1_N(_06917_),
    .Y(_06918_));
 sky130_fd_sc_hd__nand2_2 _28540_ (.A(_06906_),
    .B(_06910_),
    .Y(_06919_));
 sky130_fd_sc_hd__nand2_2 _28541_ (.A(_06919_),
    .B(_06911_),
    .Y(_06920_));
 sky130_fd_sc_hd__nand3_2 _28542_ (.A(_06906_),
    .B(_06912_),
    .C(_06910_),
    .Y(_06921_));
 sky130_fd_sc_hd__nand3_2 _28543_ (.A(_06920_),
    .B(_06921_),
    .C(_06917_),
    .Y(_06922_));
 sky130_fd_sc_hd__buf_1 _28544_ (.A(_18856_),
    .X(_06923_));
 sky130_fd_sc_hd__buf_1 _28545_ (.A(_19225_),
    .X(_06924_));
 sky130_fd_sc_hd__nand2_2 _28546_ (.A(_05953_),
    .B(_06924_),
    .Y(_06925_));
 sky130_fd_sc_hd__nand2_2 _28547_ (.A(_05956_),
    .B(_06735_),
    .Y(_06926_));
 sky130_fd_sc_hd__xnor2_2 _28548_ (.A(_06925_),
    .B(_06926_),
    .Y(_06927_));
 sky130_fd_sc_hd__o21ai_2 _28549_ (.A1(_06923_),
    .A2(_19234_),
    .B1(_06927_),
    .Y(_06928_));
 sky130_fd_sc_hd__xor2_2 _28550_ (.A(_06925_),
    .B(_06926_),
    .X(_06929_));
 sky130_fd_sc_hd__and2_2 _28551_ (.A(_06460_),
    .B(_06608_),
    .X(_06930_));
 sky130_fd_sc_hd__nand2_2 _28552_ (.A(_06929_),
    .B(_06930_),
    .Y(_06931_));
 sky130_fd_sc_hd__nand2_2 _28553_ (.A(_06586_),
    .B(_06729_),
    .Y(_06932_));
 sky130_fd_sc_hd__nand2_2 _28554_ (.A(_18850_),
    .B(_06351_),
    .Y(_06933_));
 sky130_fd_sc_hd__nor2_2 _28555_ (.A(_06932_),
    .B(_06933_),
    .Y(_06934_));
 sky130_fd_sc_hd__buf_1 _28556_ (.A(\pcpi_mul.rs1[17] ),
    .X(_06935_));
 sky130_fd_sc_hd__buf_1 _28557_ (.A(_06935_),
    .X(_06936_));
 sky130_fd_sc_hd__buf_1 _28558_ (.A(_06936_),
    .X(_06937_));
 sky130_fd_sc_hd__and2_2 _28559_ (.A(_06349_),
    .B(_06937_),
    .X(_06938_));
 sky130_fd_sc_hd__nand2_2 _28560_ (.A(_06932_),
    .B(_06933_),
    .Y(_06939_));
 sky130_fd_sc_hd__nand3b_2 _28561_ (.A_N(_06934_),
    .B(_06938_),
    .C(_06939_),
    .Y(_06940_));
 sky130_fd_sc_hd__a22oi_2 _28562_ (.A1(_18845_),
    .A2(_06479_),
    .B1(_05464_),
    .B2(_06617_),
    .Y(_06941_));
 sky130_fd_sc_hd__o21bai_2 _28563_ (.A1(_06941_),
    .A2(_06934_),
    .B1_N(_06938_),
    .Y(_06942_));
 sky130_fd_sc_hd__nand2_2 _28564_ (.A(_06940_),
    .B(_06942_),
    .Y(_06943_));
 sky130_fd_sc_hd__a21oi_2 _28565_ (.A1(_06737_),
    .A2(_06736_),
    .B1(_06731_),
    .Y(_06944_));
 sky130_fd_sc_hd__nand2_2 _28566_ (.A(_06943_),
    .B(_06944_),
    .Y(_06945_));
 sky130_fd_sc_hd__nand3b_2 _28567_ (.A_N(_06944_),
    .B(_06940_),
    .C(_06942_),
    .Y(_06946_));
 sky130_fd_sc_hd__a22oi_2 _28568_ (.A1(_06928_),
    .A2(_06931_),
    .B1(_06945_),
    .B2(_06946_),
    .Y(_06947_));
 sky130_fd_sc_hd__a21boi_2 _28569_ (.A1(_06940_),
    .A2(_06942_),
    .B1_N(_06944_),
    .Y(_06948_));
 sky130_fd_sc_hd__nand2_2 _28570_ (.A(_06931_),
    .B(_06928_),
    .Y(_06949_));
 sky130_fd_sc_hd__nor3b_2 _28571_ (.A(_06948_),
    .B(_06949_),
    .C_N(_06946_),
    .Y(_06950_));
 sky130_fd_sc_hd__o21ai_2 _28572_ (.A1(_06742_),
    .A2(_06753_),
    .B1(_06754_),
    .Y(_06951_));
 sky130_fd_sc_hd__o21bai_2 _28573_ (.A1(_06947_),
    .A2(_06950_),
    .B1_N(_06951_),
    .Y(_06952_));
 sky130_fd_sc_hd__nand3b_2 _28574_ (.A_N(_06949_),
    .B(_06946_),
    .C(_06945_),
    .Y(_06953_));
 sky130_fd_sc_hd__nand3b_2 _28575_ (.A_N(_06947_),
    .B(_06953_),
    .C(_06951_),
    .Y(_06954_));
 sky130_fd_sc_hd__nand2_2 _28576_ (.A(_06952_),
    .B(_06954_),
    .Y(_06955_));
 sky130_fd_sc_hd__nor2_2 _28577_ (.A(_06743_),
    .B(_06747_),
    .Y(_06956_));
 sky130_fd_sc_hd__a21oi_2 _28578_ (.A1(_06748_),
    .A2(_06749_),
    .B1(_06956_),
    .Y(_06957_));
 sky130_fd_sc_hd__nand2_2 _28579_ (.A(_06955_),
    .B(_06957_),
    .Y(_06958_));
 sky130_vsdinv _28580_ (.A(_06957_),
    .Y(_06959_));
 sky130_fd_sc_hd__nand3_2 _28581_ (.A(_06952_),
    .B(_06954_),
    .C(_06959_),
    .Y(_06960_));
 sky130_fd_sc_hd__and2_2 _28582_ (.A(_06958_),
    .B(_06960_),
    .X(_06961_));
 sky130_fd_sc_hd__a21oi_2 _28583_ (.A1(_06918_),
    .A2(_06922_),
    .B1(_06961_),
    .Y(_06962_));
 sky130_fd_sc_hd__nand2_2 _28584_ (.A(_06958_),
    .B(_06960_),
    .Y(_06963_));
 sky130_fd_sc_hd__a21oi_2 _28585_ (.A1(_06920_),
    .A2(_06921_),
    .B1(_06917_),
    .Y(_06964_));
 sky130_vsdinv _28586_ (.A(_06922_),
    .Y(_06965_));
 sky130_fd_sc_hd__nor3_2 _28587_ (.A(_06963_),
    .B(_06964_),
    .C(_06965_),
    .Y(_06966_));
 sky130_fd_sc_hd__nand3b_2 _28588_ (.A_N(_06845_),
    .B(_06809_),
    .C(_06846_),
    .Y(_06967_));
 sky130_vsdinv _28589_ (.A(_06967_),
    .Y(_06968_));
 sky130_fd_sc_hd__o21bai_2 _28590_ (.A1(_06962_),
    .A2(_06966_),
    .B1_N(_06968_),
    .Y(_06969_));
 sky130_fd_sc_hd__nand2_2 _28591_ (.A(_06918_),
    .B(_06922_),
    .Y(_06970_));
 sky130_fd_sc_hd__nand2_2 _28592_ (.A(_06970_),
    .B(_06963_),
    .Y(_06971_));
 sky130_fd_sc_hd__nand3_2 _28593_ (.A(_06961_),
    .B(_06918_),
    .C(_06922_),
    .Y(_06972_));
 sky130_fd_sc_hd__nand3_2 _28594_ (.A(_06971_),
    .B(_06968_),
    .C(_06972_),
    .Y(_06973_));
 sky130_vsdinv _28595_ (.A(_06799_),
    .Y(_06974_));
 sky130_fd_sc_hd__a31o_2 _28596_ (.A1(_06798_),
    .A2(_06765_),
    .A3(_06766_),
    .B1(_06974_),
    .X(_06975_));
 sky130_fd_sc_hd__a21oi_2 _28597_ (.A1(_06969_),
    .A2(_06973_),
    .B1(_06975_),
    .Y(_06976_));
 sky130_fd_sc_hd__o211a_2 _28598_ (.A1(_06974_),
    .A2(_06803_),
    .B1(_06973_),
    .C1(_06969_),
    .X(_06977_));
 sky130_fd_sc_hd__nand2_2 _28599_ (.A(_06146_),
    .B(_05930_),
    .Y(_06978_));
 sky130_fd_sc_hd__buf_1 _28600_ (.A(_05836_),
    .X(_06979_));
 sky130_fd_sc_hd__nand2_2 _28601_ (.A(_18818_),
    .B(_06979_),
    .Y(_06980_));
 sky130_fd_sc_hd__nor2_2 _28602_ (.A(_06978_),
    .B(_06980_),
    .Y(_06981_));
 sky130_fd_sc_hd__nand2_2 _28603_ (.A(_06978_),
    .B(_06980_),
    .Y(_06982_));
 sky130_vsdinv _28604_ (.A(_06982_),
    .Y(_06983_));
 sky130_fd_sc_hd__and2_2 _28605_ (.A(_05894_),
    .B(_19261_),
    .X(_06984_));
 sky130_fd_sc_hd__o21bai_2 _28606_ (.A1(_06981_),
    .A2(_06983_),
    .B1_N(_06984_),
    .Y(_06985_));
 sky130_fd_sc_hd__nand3b_2 _28607_ (.A_N(_06981_),
    .B(_06984_),
    .C(_06982_),
    .Y(_06986_));
 sky130_fd_sc_hd__nand2_2 _28608_ (.A(_06985_),
    .B(_06986_),
    .Y(_06987_));
 sky130_fd_sc_hd__nand2_2 _28609_ (.A(_06544_),
    .B(_05644_),
    .Y(_06988_));
 sky130_fd_sc_hd__nand2_2 _28610_ (.A(_06540_),
    .B(_05533_),
    .Y(_06989_));
 sky130_fd_sc_hd__nor2_2 _28611_ (.A(_06988_),
    .B(_06989_),
    .Y(_06990_));
 sky130_fd_sc_hd__buf_1 _28612_ (.A(_05517_),
    .X(_06991_));
 sky130_fd_sc_hd__and2_2 _28613_ (.A(_18808_),
    .B(_06991_),
    .X(_06992_));
 sky130_fd_sc_hd__nand2_2 _28614_ (.A(_06988_),
    .B(_06989_),
    .Y(_06993_));
 sky130_fd_sc_hd__nand3b_2 _28615_ (.A_N(_06990_),
    .B(_06992_),
    .C(_06993_),
    .Y(_06994_));
 sky130_fd_sc_hd__a22oi_2 _28616_ (.A1(_06545_),
    .A2(_05445_),
    .B1(_06541_),
    .B2(_05997_),
    .Y(_06995_));
 sky130_fd_sc_hd__o21bai_2 _28617_ (.A1(_06995_),
    .A2(_06990_),
    .B1_N(_06992_),
    .Y(_06996_));
 sky130_fd_sc_hd__a21oi_2 _28618_ (.A1(_06831_),
    .A2(_06830_),
    .B1(_06829_),
    .Y(_06997_));
 sky130_fd_sc_hd__a21boi_2 _28619_ (.A1(_06994_),
    .A2(_06996_),
    .B1_N(_06997_),
    .Y(_06998_));
 sky130_fd_sc_hd__nand3b_2 _28620_ (.A_N(_06997_),
    .B(_06994_),
    .C(_06996_),
    .Y(_06999_));
 sky130_fd_sc_hd__nor3b_2 _28621_ (.A(_06987_),
    .B(_06998_),
    .C_N(_06999_),
    .Y(_07000_));
 sky130_vsdinv _28622_ (.A(_06998_),
    .Y(_07001_));
 sky130_fd_sc_hd__a21boi_2 _28623_ (.A1(_07001_),
    .A2(_06999_),
    .B1_N(_06987_),
    .Y(_07002_));
 sky130_fd_sc_hd__nor2_2 _28624_ (.A(_06842_),
    .B(_06843_),
    .Y(_07003_));
 sky130_fd_sc_hd__buf_1 _28625_ (.A(_18784_),
    .X(_07004_));
 sky130_fd_sc_hd__nand2_2 _28626_ (.A(_07004_),
    .B(_19297_),
    .Y(_07005_));
 sky130_fd_sc_hd__buf_1 _28627_ (.A(_18779_),
    .X(_07006_));
 sky130_fd_sc_hd__nand2_2 _28628_ (.A(_07006_),
    .B(_19300_),
    .Y(_07007_));
 sky130_fd_sc_hd__nand2_2 _28629_ (.A(_07005_),
    .B(_07007_),
    .Y(_07008_));
 sky130_fd_sc_hd__nor2_2 _28630_ (.A(_07005_),
    .B(_07007_),
    .Y(_07009_));
 sky130_vsdinv _28631_ (.A(_07009_),
    .Y(_07010_));
 sky130_fd_sc_hd__o2bb2ai_2 _28632_ (.A1_N(_07008_),
    .A2_N(_07010_),
    .B1(_18793_),
    .B2(_19294_),
    .Y(_07011_));
 sky130_fd_sc_hd__buf_1 _28633_ (.A(_18789_),
    .X(_07012_));
 sky130_fd_sc_hd__buf_1 _28634_ (.A(_19292_),
    .X(_07013_));
 sky130_fd_sc_hd__and2_2 _28635_ (.A(_07012_),
    .B(_07013_),
    .X(_07014_));
 sky130_fd_sc_hd__nand3b_2 _28636_ (.A_N(_07009_),
    .B(_07014_),
    .C(_07008_),
    .Y(_07015_));
 sky130_fd_sc_hd__nand2_2 _28637_ (.A(_07011_),
    .B(_07015_),
    .Y(_07016_));
 sky130_fd_sc_hd__xnor2_2 _28638_ (.A(_07003_),
    .B(_07016_),
    .Y(_07017_));
 sky130_fd_sc_hd__nor3b_2 _28639_ (.A(_07000_),
    .B(_07002_),
    .C_N(_07017_),
    .Y(_07018_));
 sky130_fd_sc_hd__o21ba_2 _28640_ (.A1(_07000_),
    .A2(_07002_),
    .B1_N(_07017_),
    .X(_07019_));
 sky130_fd_sc_hd__or2_2 _28641_ (.A(_07018_),
    .B(_07019_),
    .X(_07020_));
 sky130_fd_sc_hd__xor2_2 _28642_ (.A(_06846_),
    .B(_07020_),
    .X(_07021_));
 sky130_fd_sc_hd__o21bai_2 _28643_ (.A1(_06976_),
    .A2(_06977_),
    .B1_N(_07021_),
    .Y(_07022_));
 sky130_fd_sc_hd__a21oi_2 _28644_ (.A1(_06971_),
    .A2(_06972_),
    .B1(_06968_),
    .Y(_07023_));
 sky130_fd_sc_hd__nor3_2 _28645_ (.A(_06967_),
    .B(_06962_),
    .C(_06966_),
    .Y(_07024_));
 sky130_fd_sc_hd__o21bai_2 _28646_ (.A1(_07023_),
    .A2(_07024_),
    .B1_N(_06975_),
    .Y(_07025_));
 sky130_fd_sc_hd__nand3_2 _28647_ (.A(_06969_),
    .B(_06975_),
    .C(_06973_),
    .Y(_07026_));
 sky130_fd_sc_hd__nand3_2 _28648_ (.A(_07025_),
    .B(_07021_),
    .C(_07026_),
    .Y(_07027_));
 sky130_fd_sc_hd__buf_1 _28649_ (.A(_06851_),
    .X(_07028_));
 sky130_fd_sc_hd__a21oi_2 _28650_ (.A1(_07022_),
    .A2(_07027_),
    .B1(_07028_),
    .Y(_07029_));
 sky130_fd_sc_hd__a21oi_2 _28651_ (.A1(_07025_),
    .A2(_07026_),
    .B1(_07021_),
    .Y(_07030_));
 sky130_vsdinv _28652_ (.A(_07021_),
    .Y(_07031_));
 sky130_fd_sc_hd__nor3_2 _28653_ (.A(_07031_),
    .B(_06976_),
    .C(_06977_),
    .Y(_07032_));
 sky130_fd_sc_hd__nor3_2 _28654_ (.A(_06850_),
    .B(_07030_),
    .C(_07032_),
    .Y(_07033_));
 sky130_fd_sc_hd__a21boi_2 _28655_ (.A1(_06758_),
    .A2(_06764_),
    .B1_N(_06761_),
    .Y(_07034_));
 sky130_fd_sc_hd__xor2_2 _28656_ (.A(_07034_),
    .B(_06853_),
    .X(_07035_));
 sky130_fd_sc_hd__o21bai_2 _28657_ (.A1(_07029_),
    .A2(_07033_),
    .B1_N(_07035_),
    .Y(_07036_));
 sky130_fd_sc_hd__o21bai_2 _28658_ (.A1(_07030_),
    .A2(_07032_),
    .B1_N(_07028_),
    .Y(_07037_));
 sky130_fd_sc_hd__nand3_2 _28659_ (.A(_07022_),
    .B(_07028_),
    .C(_07027_),
    .Y(_07038_));
 sky130_fd_sc_hd__nand3_2 _28660_ (.A(_07037_),
    .B(_07035_),
    .C(_07038_),
    .Y(_07039_));
 sky130_fd_sc_hd__nor3_2 _28661_ (.A(_06710_),
    .B(_06849_),
    .C(_07028_),
    .Y(_07040_));
 sky130_fd_sc_hd__a21oi_2 _28662_ (.A1(_06852_),
    .A2(_06857_),
    .B1(_07040_),
    .Y(_07041_));
 sky130_vsdinv _28663_ (.A(_07041_),
    .Y(_07042_));
 sky130_fd_sc_hd__a21oi_2 _28664_ (.A1(_07036_),
    .A2(_07039_),
    .B1(_07042_),
    .Y(_07043_));
 sky130_fd_sc_hd__a21oi_2 _28665_ (.A1(_07037_),
    .A2(_07038_),
    .B1(_07035_),
    .Y(_07044_));
 sky130_vsdinv _28666_ (.A(_07039_),
    .Y(_07045_));
 sky130_fd_sc_hd__nor3_2 _28667_ (.A(_07041_),
    .B(_07044_),
    .C(_07045_),
    .Y(_07046_));
 sky130_fd_sc_hd__nor2_2 _28668_ (.A(_06856_),
    .B(_06664_),
    .Y(_07047_));
 sky130_fd_sc_hd__o21bai_2 _28669_ (.A1(_07043_),
    .A2(_07046_),
    .B1_N(_07047_),
    .Y(_07048_));
 sky130_fd_sc_hd__o21bai_2 _28670_ (.A1(_07044_),
    .A2(_07045_),
    .B1_N(_07042_),
    .Y(_07049_));
 sky130_fd_sc_hd__nand3_2 _28671_ (.A(_07036_),
    .B(_07042_),
    .C(_07039_),
    .Y(_07050_));
 sky130_fd_sc_hd__nand3_2 _28672_ (.A(_07049_),
    .B(_07047_),
    .C(_07050_),
    .Y(_07051_));
 sky130_fd_sc_hd__nand2_2 _28673_ (.A(_06868_),
    .B(_06863_),
    .Y(_07052_));
 sky130_fd_sc_hd__a21oi_2 _28674_ (.A1(_07048_),
    .A2(_07051_),
    .B1(_07052_),
    .Y(_07053_));
 sky130_vsdinv _28675_ (.A(_07053_),
    .Y(_07054_));
 sky130_fd_sc_hd__nand3_2 _28676_ (.A(_07048_),
    .B(_07051_),
    .C(_07052_),
    .Y(_07055_));
 sky130_fd_sc_hd__nand2_2 _28677_ (.A(_07054_),
    .B(_07055_),
    .Y(_07056_));
 sky130_fd_sc_hd__a21boi_2 _28678_ (.A1(_06878_),
    .A2(_06871_),
    .B1_N(_06873_),
    .Y(_07057_));
 sky130_fd_sc_hd__xor2_2 _28679_ (.A(_07056_),
    .B(_07057_),
    .X(_02636_));
 sky130_fd_sc_hd__buf_1 _28680_ (.A(\pcpi_mul.rs2[8] ),
    .X(_07058_));
 sky130_fd_sc_hd__buf_1 _28681_ (.A(_07058_),
    .X(_07059_));
 sky130_fd_sc_hd__buf_1 _28682_ (.A(_06046_),
    .X(_07060_));
 sky130_fd_sc_hd__a22oi_2 _28683_ (.A1(_07059_),
    .A2(_06063_),
    .B1(_06096_),
    .B2(_07060_),
    .Y(_07061_));
 sky130_fd_sc_hd__nand2_2 _28684_ (.A(_07058_),
    .B(_06062_),
    .Y(_07062_));
 sky130_fd_sc_hd__nand2_2 _28685_ (.A(_05767_),
    .B(_06202_),
    .Y(_07063_));
 sky130_fd_sc_hd__nor2_2 _28686_ (.A(_07062_),
    .B(_07063_),
    .Y(_07064_));
 sky130_fd_sc_hd__and2_2 _28687_ (.A(_18838_),
    .B(_06364_),
    .X(_07065_));
 sky130_fd_sc_hd__o21bai_2 _28688_ (.A1(_07061_),
    .A2(_07064_),
    .B1_N(_07065_),
    .Y(_07066_));
 sky130_fd_sc_hd__nand3b_2 _28689_ (.A_N(_07062_),
    .B(_06889_),
    .C(_06047_),
    .Y(_07067_));
 sky130_fd_sc_hd__nand2_2 _28690_ (.A(_07062_),
    .B(_07063_),
    .Y(_07068_));
 sky130_fd_sc_hd__nand3_2 _28691_ (.A(_07067_),
    .B(_07065_),
    .C(_07068_),
    .Y(_07069_));
 sky130_fd_sc_hd__nand2_2 _28692_ (.A(_07066_),
    .B(_07069_),
    .Y(_07070_));
 sky130_fd_sc_hd__a21oi_2 _28693_ (.A1(_06982_),
    .A2(_06984_),
    .B1(_06981_),
    .Y(_07071_));
 sky130_fd_sc_hd__nand2_2 _28694_ (.A(_07070_),
    .B(_07071_),
    .Y(_07072_));
 sky130_fd_sc_hd__buf_1 _28695_ (.A(_07072_),
    .X(_07073_));
 sky130_fd_sc_hd__nand3b_2 _28696_ (.A_N(_07071_),
    .B(_07069_),
    .C(_07066_),
    .Y(_07074_));
 sky130_fd_sc_hd__buf_1 _28697_ (.A(_07074_),
    .X(_07075_));
 sky130_fd_sc_hd__a21oi_2 _28698_ (.A1(_06892_),
    .A2(_06887_),
    .B1(_06885_),
    .Y(_07076_));
 sky130_vsdinv _28699_ (.A(_07076_),
    .Y(_07077_));
 sky130_fd_sc_hd__a21oi_2 _28700_ (.A1(_07073_),
    .A2(_07075_),
    .B1(_07077_),
    .Y(_07078_));
 sky130_vsdinv _28701_ (.A(_06893_),
    .Y(_07079_));
 sky130_fd_sc_hd__o211a_2 _28702_ (.A1(_06885_),
    .A2(_07079_),
    .B1(_07075_),
    .C1(_07073_),
    .X(_07080_));
 sky130_fd_sc_hd__o21ai_2 _28703_ (.A1(_06987_),
    .A2(_06998_),
    .B1(_06999_),
    .Y(_07081_));
 sky130_fd_sc_hd__o21bai_2 _28704_ (.A1(_07078_),
    .A2(_07080_),
    .B1_N(_07081_),
    .Y(_07082_));
 sky130_fd_sc_hd__a21o_2 _28705_ (.A1(_07072_),
    .A2(_07074_),
    .B1(_07077_),
    .X(_07083_));
 sky130_fd_sc_hd__nand3_2 _28706_ (.A(_07073_),
    .B(_07077_),
    .C(_07075_),
    .Y(_07084_));
 sky130_fd_sc_hd__nand3_2 _28707_ (.A(_07083_),
    .B(_07081_),
    .C(_07084_),
    .Y(_07085_));
 sky130_fd_sc_hd__buf_1 _28708_ (.A(_07085_),
    .X(_07086_));
 sky130_fd_sc_hd__a21oi_2 _28709_ (.A1(_06897_),
    .A2(_06900_),
    .B1(_06903_),
    .Y(_07087_));
 sky130_vsdinv _28710_ (.A(_07087_),
    .Y(_07088_));
 sky130_fd_sc_hd__a21oi_2 _28711_ (.A1(_07082_),
    .A2(_07086_),
    .B1(_07088_),
    .Y(_07089_));
 sky130_fd_sc_hd__o211a_2 _28712_ (.A1(_06903_),
    .A2(_06904_),
    .B1(_07086_),
    .C1(_07082_),
    .X(_07090_));
 sky130_fd_sc_hd__a21oi_2 _28713_ (.A1(_06907_),
    .A2(_06908_),
    .B1(_06905_),
    .Y(_07091_));
 sky130_fd_sc_hd__o21ai_2 _28714_ (.A1(_06911_),
    .A2(_07091_),
    .B1(_06909_),
    .Y(_07092_));
 sky130_fd_sc_hd__o21bai_2 _28715_ (.A1(_07089_),
    .A2(_07090_),
    .B1_N(_07092_),
    .Y(_07093_));
 sky130_fd_sc_hd__nand2_2 _28716_ (.A(_07082_),
    .B(_07085_),
    .Y(_07094_));
 sky130_fd_sc_hd__nand2_2 _28717_ (.A(_07094_),
    .B(_07087_),
    .Y(_07095_));
 sky130_fd_sc_hd__nand3_2 _28718_ (.A(_07082_),
    .B(_07088_),
    .C(_07086_),
    .Y(_07096_));
 sky130_fd_sc_hd__nand3_2 _28719_ (.A(_07095_),
    .B(_07096_),
    .C(_07092_),
    .Y(_07097_));
 sky130_fd_sc_hd__buf_1 _28720_ (.A(\pcpi_mul.rs1[13] ),
    .X(_07098_));
 sky130_fd_sc_hd__buf_1 _28721_ (.A(_07098_),
    .X(_07099_));
 sky130_fd_sc_hd__buf_1 _28722_ (.A(_07099_),
    .X(_07100_));
 sky130_fd_sc_hd__nand2_2 _28723_ (.A(_05813_),
    .B(_07100_),
    .Y(_07101_));
 sky130_fd_sc_hd__buf_1 _28724_ (.A(_06606_),
    .X(_07102_));
 sky130_fd_sc_hd__nand2_2 _28725_ (.A(_05816_),
    .B(_07102_),
    .Y(_07103_));
 sky130_fd_sc_hd__nor2_2 _28726_ (.A(_07101_),
    .B(_07103_),
    .Y(_07104_));
 sky130_fd_sc_hd__buf_1 _28727_ (.A(\pcpi_mul.rs1[18] ),
    .X(_07105_));
 sky130_fd_sc_hd__buf_1 _28728_ (.A(_07105_),
    .X(_07106_));
 sky130_fd_sc_hd__and2_2 _28729_ (.A(_18878_),
    .B(_07106_),
    .X(_07107_));
 sky130_fd_sc_hd__nand2_2 _28730_ (.A(_07101_),
    .B(_07103_),
    .Y(_07108_));
 sky130_fd_sc_hd__nand3b_2 _28731_ (.A_N(_07104_),
    .B(_07107_),
    .C(_07108_),
    .Y(_07109_));
 sky130_fd_sc_hd__a22oi_2 _28732_ (.A1(_05825_),
    .A2(_06467_),
    .B1(_05940_),
    .B2(_06608_),
    .Y(_07110_));
 sky130_fd_sc_hd__o21bai_2 _28733_ (.A1(_07110_),
    .A2(_07104_),
    .B1_N(_07107_),
    .Y(_07111_));
 sky130_fd_sc_hd__a21o_2 _28734_ (.A1(_06939_),
    .A2(_06938_),
    .B1(_06934_),
    .X(_07112_));
 sky130_fd_sc_hd__a21o_2 _28735_ (.A1(_07109_),
    .A2(_07111_),
    .B1(_07112_),
    .X(_07113_));
 sky130_fd_sc_hd__nand3_2 _28736_ (.A(_07109_),
    .B(_07111_),
    .C(_07112_),
    .Y(_07114_));
 sky130_fd_sc_hd__buf_1 _28737_ (.A(_06733_),
    .X(_07115_));
 sky130_fd_sc_hd__buf_1 _28738_ (.A(_07115_),
    .X(_07116_));
 sky130_fd_sc_hd__nand2_2 _28739_ (.A(_05421_),
    .B(_07116_),
    .Y(_07117_));
 sky130_fd_sc_hd__buf_1 _28740_ (.A(_19211_),
    .X(_07118_));
 sky130_fd_sc_hd__nand2_2 _28741_ (.A(_05428_),
    .B(_07118_),
    .Y(_07119_));
 sky130_fd_sc_hd__xor2_2 _28742_ (.A(_07117_),
    .B(_07119_),
    .X(_07120_));
 sky130_fd_sc_hd__buf_1 _28743_ (.A(_06073_),
    .X(_07121_));
 sky130_fd_sc_hd__and2_2 _28744_ (.A(_07121_),
    .B(_06746_),
    .X(_07122_));
 sky130_fd_sc_hd__nand2_2 _28745_ (.A(_07120_),
    .B(_07122_),
    .Y(_07123_));
 sky130_fd_sc_hd__xnor2_2 _28746_ (.A(_07117_),
    .B(_07119_),
    .Y(_07124_));
 sky130_fd_sc_hd__o21ai_2 _28747_ (.A1(_18857_),
    .A2(_19228_),
    .B1(_07124_),
    .Y(_07125_));
 sky130_fd_sc_hd__nand2_2 _28748_ (.A(_07123_),
    .B(_07125_),
    .Y(_07126_));
 sky130_fd_sc_hd__a21boi_2 _28749_ (.A1(_07113_),
    .A2(_07114_),
    .B1_N(_07126_),
    .Y(_07127_));
 sky130_fd_sc_hd__a21oi_2 _28750_ (.A1(_07109_),
    .A2(_07111_),
    .B1(_07112_),
    .Y(_07128_));
 sky130_fd_sc_hd__nor3b_2 _28751_ (.A(_07128_),
    .B(_07126_),
    .C_N(_07114_),
    .Y(_07129_));
 sky130_fd_sc_hd__o21ai_2 _28752_ (.A1(_06948_),
    .A2(_06949_),
    .B1(_06946_),
    .Y(_07130_));
 sky130_fd_sc_hd__o21bai_2 _28753_ (.A1(_07127_),
    .A2(_07129_),
    .B1_N(_07130_),
    .Y(_07131_));
 sky130_fd_sc_hd__nand3b_2 _28754_ (.A_N(_07126_),
    .B(_07114_),
    .C(_07113_),
    .Y(_07132_));
 sky130_fd_sc_hd__nand3b_2 _28755_ (.A_N(_07127_),
    .B(_07132_),
    .C(_07130_),
    .Y(_07133_));
 sky130_fd_sc_hd__nor2_2 _28756_ (.A(_06925_),
    .B(_06926_),
    .Y(_07134_));
 sky130_fd_sc_hd__a21oi_2 _28757_ (.A1(_06929_),
    .A2(_06930_),
    .B1(_07134_),
    .Y(_07135_));
 sky130_vsdinv _28758_ (.A(_07135_),
    .Y(_07136_));
 sky130_fd_sc_hd__a21oi_2 _28759_ (.A1(_07131_),
    .A2(_07133_),
    .B1(_07136_),
    .Y(_07137_));
 sky130_fd_sc_hd__nand3_2 _28760_ (.A(_07131_),
    .B(_07133_),
    .C(_07136_),
    .Y(_07138_));
 sky130_vsdinv _28761_ (.A(_07138_),
    .Y(_07139_));
 sky130_fd_sc_hd__nor2_2 _28762_ (.A(_07137_),
    .B(_07139_),
    .Y(_07140_));
 sky130_fd_sc_hd__a21oi_2 _28763_ (.A1(_07093_),
    .A2(_07097_),
    .B1(_07140_),
    .Y(_07141_));
 sky130_fd_sc_hd__nand2_2 _28764_ (.A(_07131_),
    .B(_07133_),
    .Y(_07142_));
 sky130_fd_sc_hd__nand2_2 _28765_ (.A(_07142_),
    .B(_07135_),
    .Y(_07143_));
 sky130_fd_sc_hd__nand2_2 _28766_ (.A(_07143_),
    .B(_07138_),
    .Y(_07144_));
 sky130_fd_sc_hd__a21oi_2 _28767_ (.A1(_07095_),
    .A2(_07096_),
    .B1(_07092_),
    .Y(_07145_));
 sky130_vsdinv _28768_ (.A(_07097_),
    .Y(_07146_));
 sky130_fd_sc_hd__nor3_2 _28769_ (.A(_07144_),
    .B(_07145_),
    .C(_07146_),
    .Y(_07147_));
 sky130_fd_sc_hd__nor3_2 _28770_ (.A(_06846_),
    .B(_07018_),
    .C(_07019_),
    .Y(_07148_));
 sky130_fd_sc_hd__o21bai_2 _28771_ (.A1(_07141_),
    .A2(_07147_),
    .B1_N(_07148_),
    .Y(_07149_));
 sky130_fd_sc_hd__nand2_2 _28772_ (.A(_07093_),
    .B(_07097_),
    .Y(_07150_));
 sky130_fd_sc_hd__nand2_2 _28773_ (.A(_07150_),
    .B(_07144_),
    .Y(_07151_));
 sky130_fd_sc_hd__nand3_2 _28774_ (.A(_07140_),
    .B(_07093_),
    .C(_07097_),
    .Y(_07152_));
 sky130_fd_sc_hd__nand3_2 _28775_ (.A(_07151_),
    .B(_07148_),
    .C(_07152_),
    .Y(_07153_));
 sky130_fd_sc_hd__a21oi_2 _28776_ (.A1(_06961_),
    .A2(_06918_),
    .B1(_06965_),
    .Y(_07154_));
 sky130_vsdinv _28777_ (.A(_07154_),
    .Y(_07155_));
 sky130_fd_sc_hd__a21oi_2 _28778_ (.A1(_07149_),
    .A2(_07153_),
    .B1(_07155_),
    .Y(_07156_));
 sky130_fd_sc_hd__a21oi_2 _28779_ (.A1(_07151_),
    .A2(_07152_),
    .B1(_07148_),
    .Y(_07157_));
 sky130_vsdinv _28780_ (.A(_07148_),
    .Y(_07158_));
 sky130_fd_sc_hd__nor3_2 _28781_ (.A(_07158_),
    .B(_07141_),
    .C(_07147_),
    .Y(_07159_));
 sky130_fd_sc_hd__nor3_2 _28782_ (.A(_07154_),
    .B(_07157_),
    .C(_07159_),
    .Y(_07160_));
 sky130_fd_sc_hd__buf_1 _28783_ (.A(_18775_),
    .X(_07161_));
 sky130_fd_sc_hd__buf_1 _28784_ (.A(_07161_),
    .X(_07162_));
 sky130_fd_sc_hd__and2_2 _28785_ (.A(_07162_),
    .B(_05243_),
    .X(_07163_));
 sky130_fd_sc_hd__buf_1 _28786_ (.A(\pcpi_mul.rs2[17] ),
    .X(_07164_));
 sky130_fd_sc_hd__buf_1 _28787_ (.A(_07164_),
    .X(_07165_));
 sky130_fd_sc_hd__nand2_2 _28788_ (.A(_07165_),
    .B(_05401_),
    .Y(_07166_));
 sky130_fd_sc_hd__buf_1 _28789_ (.A(\pcpi_mul.rs2[16] ),
    .X(_07167_));
 sky130_fd_sc_hd__buf_1 _28790_ (.A(_07167_),
    .X(_07168_));
 sky130_fd_sc_hd__nand2_2 _28791_ (.A(_07168_),
    .B(_05635_),
    .Y(_07169_));
 sky130_fd_sc_hd__nor2_2 _28792_ (.A(_07166_),
    .B(_07169_),
    .Y(_07170_));
 sky130_fd_sc_hd__buf_1 _28793_ (.A(_05443_),
    .X(_07171_));
 sky130_fd_sc_hd__and2_2 _28794_ (.A(_18790_),
    .B(_07171_),
    .X(_07172_));
 sky130_vsdinv _28795_ (.A(_07172_),
    .Y(_07173_));
 sky130_fd_sc_hd__nand2_2 _28796_ (.A(_07166_),
    .B(_07169_),
    .Y(_07174_));
 sky130_fd_sc_hd__nor3b_2 _28797_ (.A(_07170_),
    .B(_07173_),
    .C_N(_07174_),
    .Y(_07175_));
 sky130_vsdinv _28798_ (.A(_07175_),
    .Y(_07176_));
 sky130_vsdinv _28799_ (.A(_07170_),
    .Y(_07177_));
 sky130_fd_sc_hd__buf_1 _28800_ (.A(_18791_),
    .X(_07178_));
 sky130_fd_sc_hd__o2bb2ai_2 _28801_ (.A1_N(_07174_),
    .A2_N(_07177_),
    .B1(_07178_),
    .B2(_19289_),
    .Y(_07179_));
 sky130_fd_sc_hd__a21oi_2 _28802_ (.A1(_07008_),
    .A2(_07014_),
    .B1(_07009_),
    .Y(_07180_));
 sky130_vsdinv _28803_ (.A(_07180_),
    .Y(_07181_));
 sky130_fd_sc_hd__a21o_2 _28804_ (.A1(_07176_),
    .A2(_07179_),
    .B1(_07181_),
    .X(_07182_));
 sky130_fd_sc_hd__nand3b_2 _28805_ (.A_N(_07175_),
    .B(_07179_),
    .C(_07181_),
    .Y(_07183_));
 sky130_fd_sc_hd__buf_1 _28806_ (.A(_07183_),
    .X(_07184_));
 sky130_fd_sc_hd__nand3_2 _28807_ (.A(_07011_),
    .B(_07003_),
    .C(_07015_),
    .Y(_07185_));
 sky130_vsdinv _28808_ (.A(_07185_),
    .Y(_07186_));
 sky130_fd_sc_hd__a21oi_2 _28809_ (.A1(_07182_),
    .A2(_07184_),
    .B1(_07186_),
    .Y(_07187_));
 sky130_fd_sc_hd__nand3_2 _28810_ (.A(_07182_),
    .B(_07186_),
    .C(_07184_),
    .Y(_07188_));
 sky130_vsdinv _28811_ (.A(_07188_),
    .Y(_07189_));
 sky130_fd_sc_hd__buf_1 _28812_ (.A(_06543_),
    .X(_07190_));
 sky130_fd_sc_hd__nand2_2 _28813_ (.A(_07190_),
    .B(_05674_),
    .Y(_07191_));
 sky130_fd_sc_hd__buf_1 _28814_ (.A(\pcpi_mul.rs2[13] ),
    .X(_07192_));
 sky130_fd_sc_hd__nand2_2 _28815_ (.A(_07192_),
    .B(_05745_),
    .Y(_07193_));
 sky130_fd_sc_hd__nor2_2 _28816_ (.A(_07191_),
    .B(_07193_),
    .Y(_07194_));
 sky130_fd_sc_hd__buf_1 _28817_ (.A(_18807_),
    .X(_07195_));
 sky130_fd_sc_hd__and2_2 _28818_ (.A(_07195_),
    .B(_05500_),
    .X(_07196_));
 sky130_fd_sc_hd__nand2_2 _28819_ (.A(_07191_),
    .B(_07193_),
    .Y(_07197_));
 sky130_fd_sc_hd__nand3b_2 _28820_ (.A_N(_07194_),
    .B(_07196_),
    .C(_07197_),
    .Y(_07198_));
 sky130_fd_sc_hd__buf_1 _28821_ (.A(_06533_),
    .X(_07199_));
 sky130_fd_sc_hd__buf_1 _28822_ (.A(\pcpi_mul.rs2[13] ),
    .X(_07200_));
 sky130_fd_sc_hd__buf_1 _28823_ (.A(_07200_),
    .X(_07201_));
 sky130_fd_sc_hd__a22oi_2 _28824_ (.A1(_07199_),
    .A2(_05470_),
    .B1(_07201_),
    .B2(_05529_),
    .Y(_07202_));
 sky130_fd_sc_hd__o21bai_2 _28825_ (.A1(_07202_),
    .A2(_07194_),
    .B1_N(_07196_),
    .Y(_07203_));
 sky130_fd_sc_hd__a21oi_2 _28826_ (.A1(_06993_),
    .A2(_06992_),
    .B1(_06990_),
    .Y(_07204_));
 sky130_fd_sc_hd__a21boi_2 _28827_ (.A1(_07198_),
    .A2(_07203_),
    .B1_N(_07204_),
    .Y(_07205_));
 sky130_fd_sc_hd__nand3b_2 _28828_ (.A_N(_07204_),
    .B(_07198_),
    .C(_07203_),
    .Y(_07206_));
 sky130_vsdinv _28829_ (.A(_07206_),
    .Y(_07207_));
 sky130_fd_sc_hd__buf_1 _28830_ (.A(_05836_),
    .X(_07208_));
 sky130_fd_sc_hd__nand2_2 _28831_ (.A(_06146_),
    .B(_07208_),
    .Y(_07209_));
 sky130_fd_sc_hd__nand2_2 _28832_ (.A(_18818_),
    .B(_05840_),
    .Y(_07210_));
 sky130_fd_sc_hd__nand2_2 _28833_ (.A(_07209_),
    .B(_07210_),
    .Y(_07211_));
 sky130_fd_sc_hd__nor2_2 _28834_ (.A(_07209_),
    .B(_07210_),
    .Y(_07212_));
 sky130_vsdinv _28835_ (.A(_07212_),
    .Y(_07213_));
 sky130_fd_sc_hd__buf_1 _28836_ (.A(_18823_),
    .X(_07214_));
 sky130_fd_sc_hd__o2bb2ai_2 _28837_ (.A1_N(_07211_),
    .A2_N(_07213_),
    .B1(_07214_),
    .B2(_19259_),
    .Y(_07215_));
 sky130_fd_sc_hd__buf_1 _28838_ (.A(_19256_),
    .X(_07216_));
 sky130_fd_sc_hd__and2_2 _28839_ (.A(_05894_),
    .B(_07216_),
    .X(_07217_));
 sky130_fd_sc_hd__nand3b_2 _28840_ (.A_N(_07212_),
    .B(_07217_),
    .C(_07211_),
    .Y(_07218_));
 sky130_fd_sc_hd__nand2_2 _28841_ (.A(_07215_),
    .B(_07218_),
    .Y(_07219_));
 sky130_fd_sc_hd__o21ai_2 _28842_ (.A1(_07205_),
    .A2(_07207_),
    .B1(_07219_),
    .Y(_07220_));
 sky130_fd_sc_hd__and2_2 _28843_ (.A(_07215_),
    .B(_07218_),
    .X(_07221_));
 sky130_fd_sc_hd__nand3b_2 _28844_ (.A_N(_07205_),
    .B(_07221_),
    .C(_07206_),
    .Y(_07222_));
 sky130_fd_sc_hd__nand2_2 _28845_ (.A(_07220_),
    .B(_07222_),
    .Y(_07223_));
 sky130_fd_sc_hd__o21ai_2 _28846_ (.A1(_07187_),
    .A2(_07189_),
    .B1(_07223_),
    .Y(_07224_));
 sky130_fd_sc_hd__a21o_2 _28847_ (.A1(_07182_),
    .A2(_07184_),
    .B1(_07186_),
    .X(_07225_));
 sky130_fd_sc_hd__nand3b_2 _28848_ (.A_N(_07223_),
    .B(_07225_),
    .C(_07188_),
    .Y(_07226_));
 sky130_fd_sc_hd__a21o_2 _28849_ (.A1(_07224_),
    .A2(_07226_),
    .B1(_07018_),
    .X(_07227_));
 sky130_fd_sc_hd__nand3_2 _28850_ (.A(_07224_),
    .B(_07018_),
    .C(_07226_),
    .Y(_07228_));
 sky130_fd_sc_hd__nand2_2 _28851_ (.A(_07227_),
    .B(_07228_),
    .Y(_07229_));
 sky130_fd_sc_hd__xnor2_2 _28852_ (.A(_07163_),
    .B(_07229_),
    .Y(_07230_));
 sky130_fd_sc_hd__o21bai_2 _28853_ (.A1(_07156_),
    .A2(_07160_),
    .B1_N(_07230_),
    .Y(_07231_));
 sky130_fd_sc_hd__o21bai_2 _28854_ (.A1(_07157_),
    .A2(_07159_),
    .B1_N(_07155_),
    .Y(_07232_));
 sky130_fd_sc_hd__nand3_2 _28855_ (.A(_07149_),
    .B(_07155_),
    .C(_07153_),
    .Y(_07233_));
 sky130_fd_sc_hd__nand3_2 _28856_ (.A(_07232_),
    .B(_07230_),
    .C(_07233_),
    .Y(_07234_));
 sky130_fd_sc_hd__a21oi_2 _28857_ (.A1(_07231_),
    .A2(_07234_),
    .B1(_07032_),
    .Y(_07235_));
 sky130_fd_sc_hd__a21oi_2 _28858_ (.A1(_07232_),
    .A2(_07233_),
    .B1(_07230_),
    .Y(_07236_));
 sky130_vsdinv _28859_ (.A(_07230_),
    .Y(_07237_));
 sky130_fd_sc_hd__nor3_2 _28860_ (.A(_07237_),
    .B(_07156_),
    .C(_07160_),
    .Y(_07238_));
 sky130_fd_sc_hd__nor3_2 _28861_ (.A(_07027_),
    .B(_07236_),
    .C(_07238_),
    .Y(_07239_));
 sky130_fd_sc_hd__a21boi_2 _28862_ (.A1(_06952_),
    .A2(_06959_),
    .B1_N(_06954_),
    .Y(_07240_));
 sky130_fd_sc_hd__a21o_2 _28863_ (.A1(_06969_),
    .A2(_06975_),
    .B1(_07024_),
    .X(_07241_));
 sky130_fd_sc_hd__xnor2_2 _28864_ (.A(_07240_),
    .B(_07241_),
    .Y(_07242_));
 sky130_fd_sc_hd__o21bai_2 _28865_ (.A1(_07235_),
    .A2(_07239_),
    .B1_N(_07242_),
    .Y(_07243_));
 sky130_fd_sc_hd__o21ai_2 _28866_ (.A1(_07236_),
    .A2(_07238_),
    .B1(_07027_),
    .Y(_07244_));
 sky130_fd_sc_hd__nand3_2 _28867_ (.A(_07032_),
    .B(_07231_),
    .C(_07234_),
    .Y(_07245_));
 sky130_fd_sc_hd__nand3_2 _28868_ (.A(_07244_),
    .B(_07242_),
    .C(_07245_),
    .Y(_07246_));
 sky130_vsdinv _28869_ (.A(_07035_),
    .Y(_07247_));
 sky130_fd_sc_hd__o21ai_2 _28870_ (.A1(_07247_),
    .A2(_07029_),
    .B1(_07038_),
    .Y(_07248_));
 sky130_fd_sc_hd__nand3_2 _28871_ (.A(_07243_),
    .B(_07246_),
    .C(_07248_),
    .Y(_07249_));
 sky130_fd_sc_hd__a21oi_2 _28872_ (.A1(_07244_),
    .A2(_07245_),
    .B1(_07242_),
    .Y(_07250_));
 sky130_fd_sc_hd__xor2_2 _28873_ (.A(_07240_),
    .B(_07241_),
    .X(_07251_));
 sky130_fd_sc_hd__nor3_2 _28874_ (.A(_07251_),
    .B(_07235_),
    .C(_07239_),
    .Y(_07252_));
 sky130_fd_sc_hd__o21bai_2 _28875_ (.A1(_07250_),
    .A2(_07252_),
    .B1_N(_07248_),
    .Y(_07253_));
 sky130_fd_sc_hd__o2bb2ai_2 _28876_ (.A1_N(_07249_),
    .A2_N(_07253_),
    .B1(_06853_),
    .B2(_07034_),
    .Y(_07254_));
 sky130_fd_sc_hd__nor2_2 _28877_ (.A(_07034_),
    .B(_06853_),
    .Y(_07255_));
 sky130_fd_sc_hd__nand3_2 _28878_ (.A(_07253_),
    .B(_07255_),
    .C(_07249_),
    .Y(_07256_));
 sky130_fd_sc_hd__a21o_2 _28879_ (.A1(_07049_),
    .A2(_07047_),
    .B1(_07046_),
    .X(_07257_));
 sky130_fd_sc_hd__a21oi_2 _28880_ (.A1(_07254_),
    .A2(_07256_),
    .B1(_07257_),
    .Y(_07258_));
 sky130_fd_sc_hd__nand3_2 _28881_ (.A(_07257_),
    .B(_07254_),
    .C(_07256_),
    .Y(_07259_));
 sky130_vsdinv _28882_ (.A(_07259_),
    .Y(_07260_));
 sky130_fd_sc_hd__nor2_2 _28883_ (.A(_07258_),
    .B(_07260_),
    .Y(_07261_));
 sky130_fd_sc_hd__a21oi_2 _28884_ (.A1(_06873_),
    .A2(_07055_),
    .B1(_07053_),
    .Y(_07262_));
 sky130_fd_sc_hd__a41oi_2 _28885_ (.A1(_06874_),
    .A2(_06878_),
    .A3(_07055_),
    .A4(_07054_),
    .B1(_07262_),
    .Y(_07263_));
 sky130_fd_sc_hd__xnor2_2 _28886_ (.A(_07261_),
    .B(_07263_),
    .Y(_02637_));
 sky130_fd_sc_hd__buf_1 _28887_ (.A(_06462_),
    .X(_07264_));
 sky130_fd_sc_hd__a22oi_2 _28888_ (.A1(_05869_),
    .A2(_06588_),
    .B1(_05992_),
    .B2(_07264_),
    .Y(_07265_));
 sky130_fd_sc_hd__nand2_2 _28889_ (.A(_06880_),
    .B(_06046_),
    .Y(_07266_));
 sky130_fd_sc_hd__nand2_2 _28890_ (.A(_18832_),
    .B(_19242_),
    .Y(_07267_));
 sky130_fd_sc_hd__nor2_2 _28891_ (.A(_07266_),
    .B(_07267_),
    .Y(_07268_));
 sky130_fd_sc_hd__and2_2 _28892_ (.A(_05585_),
    .B(_19236_),
    .X(_07269_));
 sky130_fd_sc_hd__o21bai_2 _28893_ (.A1(_07265_),
    .A2(_07268_),
    .B1_N(_07269_),
    .Y(_07270_));
 sky130_fd_sc_hd__buf_1 _28894_ (.A(_06095_),
    .X(_07271_));
 sky130_fd_sc_hd__nand3b_2 _28895_ (.A_N(_07266_),
    .B(_07271_),
    .C(_06463_),
    .Y(_07272_));
 sky130_fd_sc_hd__nand2_2 _28896_ (.A(_07266_),
    .B(_07267_),
    .Y(_07273_));
 sky130_fd_sc_hd__nand3_2 _28897_ (.A(_07272_),
    .B(_07269_),
    .C(_07273_),
    .Y(_07274_));
 sky130_fd_sc_hd__nand2_2 _28898_ (.A(_07270_),
    .B(_07274_),
    .Y(_07275_));
 sky130_fd_sc_hd__a21oi_2 _28899_ (.A1(_07211_),
    .A2(_07217_),
    .B1(_07212_),
    .Y(_07276_));
 sky130_fd_sc_hd__nand2_2 _28900_ (.A(_07275_),
    .B(_07276_),
    .Y(_07277_));
 sky130_fd_sc_hd__a21o_2 _28901_ (.A1(_07211_),
    .A2(_07217_),
    .B1(_07212_),
    .X(_07278_));
 sky130_fd_sc_hd__nand3_2 _28902_ (.A(_07270_),
    .B(_07278_),
    .C(_07274_),
    .Y(_07279_));
 sky130_fd_sc_hd__nand2_2 _28903_ (.A(_07277_),
    .B(_07279_),
    .Y(_07280_));
 sky130_fd_sc_hd__a21oi_2 _28904_ (.A1(_07068_),
    .A2(_07065_),
    .B1(_07064_),
    .Y(_07281_));
 sky130_fd_sc_hd__nand2_2 _28905_ (.A(_07280_),
    .B(_07281_),
    .Y(_07282_));
 sky130_vsdinv _28906_ (.A(_07281_),
    .Y(_07283_));
 sky130_fd_sc_hd__nand3_2 _28907_ (.A(_07277_),
    .B(_07283_),
    .C(_07279_),
    .Y(_07284_));
 sky130_fd_sc_hd__nand2_2 _28908_ (.A(_07282_),
    .B(_07284_),
    .Y(_07285_));
 sky130_fd_sc_hd__o21a_2 _28909_ (.A1(_07219_),
    .A2(_07205_),
    .B1(_07206_),
    .X(_07286_));
 sky130_fd_sc_hd__nand2_2 _28910_ (.A(_07285_),
    .B(_07286_),
    .Y(_07287_));
 sky130_fd_sc_hd__o21ai_2 _28911_ (.A1(_07219_),
    .A2(_07205_),
    .B1(_07206_),
    .Y(_07288_));
 sky130_fd_sc_hd__nand3_2 _28912_ (.A(_07288_),
    .B(_07282_),
    .C(_07284_),
    .Y(_07289_));
 sky130_fd_sc_hd__buf_1 _28913_ (.A(_07289_),
    .X(_07290_));
 sky130_fd_sc_hd__a21boi_2 _28914_ (.A1(_07073_),
    .A2(_07077_),
    .B1_N(_07075_),
    .Y(_07291_));
 sky130_vsdinv _28915_ (.A(_07291_),
    .Y(_07292_));
 sky130_fd_sc_hd__a21oi_2 _28916_ (.A1(_07287_),
    .A2(_07290_),
    .B1(_07292_),
    .Y(_07293_));
 sky130_fd_sc_hd__a21oi_2 _28917_ (.A1(_07282_),
    .A2(_07284_),
    .B1(_07288_),
    .Y(_07294_));
 sky130_fd_sc_hd__nor3b_2 _28918_ (.A(_07291_),
    .B(_07294_),
    .C_N(_07290_),
    .Y(_07295_));
 sky130_fd_sc_hd__a21oi_2 _28919_ (.A1(_07083_),
    .A2(_07084_),
    .B1(_07081_),
    .Y(_07296_));
 sky130_fd_sc_hd__o21ai_2 _28920_ (.A1(_07087_),
    .A2(_07296_),
    .B1(_07086_),
    .Y(_07297_));
 sky130_fd_sc_hd__o21bai_2 _28921_ (.A1(_07293_),
    .A2(_07295_),
    .B1_N(_07297_),
    .Y(_07298_));
 sky130_fd_sc_hd__nand2_2 _28922_ (.A(_07287_),
    .B(_07289_),
    .Y(_07299_));
 sky130_fd_sc_hd__nand2_2 _28923_ (.A(_07299_),
    .B(_07291_),
    .Y(_07300_));
 sky130_fd_sc_hd__nand3_2 _28924_ (.A(_07287_),
    .B(_07292_),
    .C(_07290_),
    .Y(_07301_));
 sky130_fd_sc_hd__nand3_2 _28925_ (.A(_07300_),
    .B(_07297_),
    .C(_07301_),
    .Y(_07302_));
 sky130_fd_sc_hd__buf_1 _28926_ (.A(_07302_),
    .X(_07303_));
 sky130_fd_sc_hd__buf_1 _28927_ (.A(_06452_),
    .X(_07304_));
 sky130_fd_sc_hd__nand2_2 _28928_ (.A(_05724_),
    .B(_07304_),
    .Y(_07305_));
 sky130_fd_sc_hd__buf_1 _28929_ (.A(_19224_),
    .X(_07306_));
 sky130_fd_sc_hd__nand2_2 _28930_ (.A(_05643_),
    .B(_07306_),
    .Y(_07307_));
 sky130_fd_sc_hd__nor2_2 _28931_ (.A(_07305_),
    .B(_07307_),
    .Y(_07308_));
 sky130_fd_sc_hd__buf_1 _28932_ (.A(\pcpi_mul.rs1[19] ),
    .X(_07309_));
 sky130_fd_sc_hd__buf_1 _28933_ (.A(_07309_),
    .X(_07310_));
 sky130_fd_sc_hd__and2_2 _28934_ (.A(_05516_),
    .B(_07310_),
    .X(_07311_));
 sky130_fd_sc_hd__nand2_2 _28935_ (.A(_07305_),
    .B(_07307_),
    .Y(_07312_));
 sky130_fd_sc_hd__nand3b_2 _28936_ (.A_N(_07308_),
    .B(_07311_),
    .C(_07312_),
    .Y(_07313_));
 sky130_fd_sc_hd__buf_1 _28937_ (.A(_19231_),
    .X(_07314_));
 sky130_fd_sc_hd__a22oi_2 _28938_ (.A1(_06586_),
    .A2(_07314_),
    .B1(_05504_),
    .B2(_06924_),
    .Y(_07315_));
 sky130_fd_sc_hd__o21bai_2 _28939_ (.A1(_07315_),
    .A2(_07308_),
    .B1_N(_07311_),
    .Y(_07316_));
 sky130_fd_sc_hd__a21oi_2 _28940_ (.A1(_07108_),
    .A2(_07107_),
    .B1(_07104_),
    .Y(_07317_));
 sky130_fd_sc_hd__a21bo_2 _28941_ (.A1(_07313_),
    .A2(_07316_),
    .B1_N(_07317_),
    .X(_07318_));
 sky130_fd_sc_hd__nand3b_2 _28942_ (.A_N(_07317_),
    .B(_07313_),
    .C(_07316_),
    .Y(_07319_));
 sky130_fd_sc_hd__nand2_2 _28943_ (.A(_07318_),
    .B(_07319_),
    .Y(_07320_));
 sky130_fd_sc_hd__buf_1 _28944_ (.A(_06935_),
    .X(_07321_));
 sky130_fd_sc_hd__nand2_2 _28945_ (.A(_05531_),
    .B(_07321_),
    .Y(_07322_));
 sky130_fd_sc_hd__buf_1 _28946_ (.A(_05427_),
    .X(_07323_));
 sky130_fd_sc_hd__buf_1 _28947_ (.A(\pcpi_mul.rs1[18] ),
    .X(_07324_));
 sky130_fd_sc_hd__buf_1 _28948_ (.A(_07324_),
    .X(_07325_));
 sky130_fd_sc_hd__nand2_2 _28949_ (.A(_07323_),
    .B(_07325_),
    .Y(_07326_));
 sky130_fd_sc_hd__xor2_2 _28950_ (.A(_07322_),
    .B(_07326_),
    .X(_07327_));
 sky130_fd_sc_hd__buf_1 _28951_ (.A(_06733_),
    .X(_07328_));
 sky130_fd_sc_hd__buf_1 _28952_ (.A(_07328_),
    .X(_07329_));
 sky130_fd_sc_hd__and2_2 _28953_ (.A(_05459_),
    .B(_07329_),
    .X(_07330_));
 sky130_fd_sc_hd__nand2_2 _28954_ (.A(_07327_),
    .B(_07330_),
    .Y(_07331_));
 sky130_fd_sc_hd__buf_1 _28955_ (.A(_18855_),
    .X(_07332_));
 sky130_fd_sc_hd__xnor2_2 _28956_ (.A(_07322_),
    .B(_07326_),
    .Y(_07333_));
 sky130_fd_sc_hd__o21ai_2 _28957_ (.A1(_07332_),
    .A2(_19218_),
    .B1(_07333_),
    .Y(_07334_));
 sky130_fd_sc_hd__nand2_2 _28958_ (.A(_07331_),
    .B(_07334_),
    .Y(_07335_));
 sky130_fd_sc_hd__nand2_2 _28959_ (.A(_07320_),
    .B(_07335_),
    .Y(_07336_));
 sky130_fd_sc_hd__nand3b_2 _28960_ (.A_N(_07335_),
    .B(_07319_),
    .C(_07318_),
    .Y(_07337_));
 sky130_fd_sc_hd__o21ai_2 _28961_ (.A1(_07128_),
    .A2(_07126_),
    .B1(_07114_),
    .Y(_07338_));
 sky130_fd_sc_hd__a21o_2 _28962_ (.A1(_07336_),
    .A2(_07337_),
    .B1(_07338_),
    .X(_07339_));
 sky130_fd_sc_hd__nand3_2 _28963_ (.A(_07336_),
    .B(_07337_),
    .C(_07338_),
    .Y(_07340_));
 sky130_fd_sc_hd__nand2_2 _28964_ (.A(_07339_),
    .B(_07340_),
    .Y(_07341_));
 sky130_fd_sc_hd__nor2_2 _28965_ (.A(_07117_),
    .B(_07119_),
    .Y(_07342_));
 sky130_fd_sc_hd__a21oi_2 _28966_ (.A1(_07120_),
    .A2(_07122_),
    .B1(_07342_),
    .Y(_07343_));
 sky130_fd_sc_hd__nand2_2 _28967_ (.A(_07341_),
    .B(_07343_),
    .Y(_07344_));
 sky130_vsdinv _28968_ (.A(_07343_),
    .Y(_07345_));
 sky130_fd_sc_hd__nand3_2 _28969_ (.A(_07339_),
    .B(_07345_),
    .C(_07340_),
    .Y(_07346_));
 sky130_fd_sc_hd__nand2_2 _28970_ (.A(_07344_),
    .B(_07346_),
    .Y(_07347_));
 sky130_fd_sc_hd__buf_1 _28971_ (.A(_07347_),
    .X(_07348_));
 sky130_fd_sc_hd__a21boi_2 _28972_ (.A1(_07298_),
    .A2(_07303_),
    .B1_N(_07348_),
    .Y(_07349_));
 sky130_fd_sc_hd__a21oi_2 _28973_ (.A1(_07300_),
    .A2(_07301_),
    .B1(_07297_),
    .Y(_07350_));
 sky130_fd_sc_hd__nor3b_2 _28974_ (.A(_07348_),
    .B(_07350_),
    .C_N(_07303_),
    .Y(_07351_));
 sky130_vsdinv _28975_ (.A(_07228_),
    .Y(_07352_));
 sky130_fd_sc_hd__o21bai_2 _28976_ (.A1(_07349_),
    .A2(_07351_),
    .B1_N(_07352_),
    .Y(_07353_));
 sky130_fd_sc_hd__nand2_2 _28977_ (.A(_07298_),
    .B(_07303_),
    .Y(_07354_));
 sky130_fd_sc_hd__nand2_2 _28978_ (.A(_07354_),
    .B(_07348_),
    .Y(_07355_));
 sky130_fd_sc_hd__nand3b_2 _28979_ (.A_N(_07347_),
    .B(_07303_),
    .C(_07298_),
    .Y(_07356_));
 sky130_fd_sc_hd__nand3_2 _28980_ (.A(_07355_),
    .B(_07356_),
    .C(_07352_),
    .Y(_07357_));
 sky130_fd_sc_hd__a21oi_2 _28981_ (.A1(_07140_),
    .A2(_07093_),
    .B1(_07146_),
    .Y(_07358_));
 sky130_vsdinv _28982_ (.A(_07358_),
    .Y(_07359_));
 sky130_fd_sc_hd__a21oi_2 _28983_ (.A1(_07353_),
    .A2(_07357_),
    .B1(_07359_),
    .Y(_07360_));
 sky130_fd_sc_hd__a21oi_2 _28984_ (.A1(_07355_),
    .A2(_07356_),
    .B1(_07352_),
    .Y(_07361_));
 sky130_fd_sc_hd__nor3_2 _28985_ (.A(_07228_),
    .B(_07349_),
    .C(_07351_),
    .Y(_07362_));
 sky130_fd_sc_hd__nor3_2 _28986_ (.A(_07358_),
    .B(_07361_),
    .C(_07362_),
    .Y(_07363_));
 sky130_fd_sc_hd__nand2_2 _28987_ (.A(_18797_),
    .B(_05528_),
    .Y(_07364_));
 sky130_fd_sc_hd__buf_1 _28988_ (.A(_19271_),
    .X(_07365_));
 sky130_fd_sc_hd__nand2_2 _28989_ (.A(_07192_),
    .B(_07365_),
    .Y(_07366_));
 sky130_fd_sc_hd__nor2_2 _28990_ (.A(_07364_),
    .B(_07366_),
    .Y(_07367_));
 sky130_fd_sc_hd__and2_2 _28991_ (.A(_06274_),
    .B(_05837_),
    .X(_07368_));
 sky130_fd_sc_hd__nand2_2 _28992_ (.A(_07364_),
    .B(_07366_),
    .Y(_07369_));
 sky130_fd_sc_hd__nand3b_2 _28993_ (.A_N(_07367_),
    .B(_07368_),
    .C(_07369_),
    .Y(_07370_));
 sky130_fd_sc_hd__a22oi_2 _28994_ (.A1(_07199_),
    .A2(_05669_),
    .B1(_06537_),
    .B2(_05671_),
    .Y(_07371_));
 sky130_fd_sc_hd__o21bai_2 _28995_ (.A1(_07371_),
    .A2(_07367_),
    .B1_N(_07368_),
    .Y(_07372_));
 sky130_fd_sc_hd__a21oi_2 _28996_ (.A1(_07197_),
    .A2(_07196_),
    .B1(_07194_),
    .Y(_07373_));
 sky130_fd_sc_hd__a21boi_2 _28997_ (.A1(_07370_),
    .A2(_07372_),
    .B1_N(_07373_),
    .Y(_07374_));
 sky130_fd_sc_hd__buf_1 _28998_ (.A(_05845_),
    .X(_07375_));
 sky130_fd_sc_hd__nand2_2 _28999_ (.A(_06146_),
    .B(_07375_),
    .Y(_07376_));
 sky130_fd_sc_hd__buf_1 _29000_ (.A(_06140_),
    .X(_07377_));
 sky130_fd_sc_hd__nand2_2 _29001_ (.A(_07377_),
    .B(_05821_),
    .Y(_07378_));
 sky130_fd_sc_hd__nor2_2 _29002_ (.A(_07376_),
    .B(_07378_),
    .Y(_07379_));
 sky130_fd_sc_hd__nand2_2 _29003_ (.A(_07376_),
    .B(_07378_),
    .Y(_07380_));
 sky130_vsdinv _29004_ (.A(_07380_),
    .Y(_07381_));
 sky130_fd_sc_hd__buf_1 _29005_ (.A(_06067_),
    .X(_07382_));
 sky130_fd_sc_hd__and2_2 _29006_ (.A(_05894_),
    .B(_07382_),
    .X(_07383_));
 sky130_fd_sc_hd__o21bai_2 _29007_ (.A1(_07379_),
    .A2(_07381_),
    .B1_N(_07383_),
    .Y(_07384_));
 sky130_fd_sc_hd__nand3b_2 _29008_ (.A_N(_07379_),
    .B(_07383_),
    .C(_07380_),
    .Y(_07385_));
 sky130_fd_sc_hd__nand2_2 _29009_ (.A(_07384_),
    .B(_07385_),
    .Y(_07386_));
 sky130_vsdinv _29010_ (.A(_07386_),
    .Y(_07387_));
 sky130_fd_sc_hd__nand3b_2 _29011_ (.A_N(_07373_),
    .B(_07370_),
    .C(_07372_),
    .Y(_07388_));
 sky130_fd_sc_hd__nand3b_2 _29012_ (.A_N(_07374_),
    .B(_07387_),
    .C(_07388_),
    .Y(_07389_));
 sky130_vsdinv _29013_ (.A(_07388_),
    .Y(_07390_));
 sky130_fd_sc_hd__o21bai_2 _29014_ (.A1(_07374_),
    .A2(_07390_),
    .B1_N(_07387_),
    .Y(_07391_));
 sky130_fd_sc_hd__buf_1 _29015_ (.A(_07165_),
    .X(_07392_));
 sky130_fd_sc_hd__nand2_2 _29016_ (.A(_07392_),
    .B(_05874_),
    .Y(_07393_));
 sky130_fd_sc_hd__buf_1 _29017_ (.A(_07167_),
    .X(_07394_));
 sky130_fd_sc_hd__buf_1 _29018_ (.A(_07394_),
    .X(_07395_));
 sky130_fd_sc_hd__nand2_2 _29019_ (.A(_07395_),
    .B(_06827_),
    .Y(_07396_));
 sky130_fd_sc_hd__nand2_2 _29020_ (.A(_07393_),
    .B(_07396_),
    .Y(_07397_));
 sky130_fd_sc_hd__nor2_2 _29021_ (.A(_07393_),
    .B(_07396_),
    .Y(_07398_));
 sky130_vsdinv _29022_ (.A(_07398_),
    .Y(_07399_));
 sky130_fd_sc_hd__buf_1 _29023_ (.A(_18792_),
    .X(_07400_));
 sky130_fd_sc_hd__o2bb2ai_2 _29024_ (.A1_N(_07397_),
    .A2_N(_07399_),
    .B1(_07400_),
    .B2(_19283_),
    .Y(_07401_));
 sky130_fd_sc_hd__buf_1 _29025_ (.A(_07012_),
    .X(_07402_));
 sky130_fd_sc_hd__buf_1 _29026_ (.A(_05469_),
    .X(_07403_));
 sky130_fd_sc_hd__and2_2 _29027_ (.A(_07402_),
    .B(_07403_),
    .X(_07404_));
 sky130_fd_sc_hd__nand3b_2 _29028_ (.A_N(_07398_),
    .B(_07404_),
    .C(_07397_),
    .Y(_07405_));
 sky130_fd_sc_hd__a21oi_2 _29029_ (.A1(_07174_),
    .A2(_07172_),
    .B1(_07170_),
    .Y(_07406_));
 sky130_vsdinv _29030_ (.A(_07406_),
    .Y(_07407_));
 sky130_fd_sc_hd__a21o_2 _29031_ (.A1(_07401_),
    .A2(_07405_),
    .B1(_07407_),
    .X(_07408_));
 sky130_fd_sc_hd__nand3_2 _29032_ (.A(_07401_),
    .B(_07405_),
    .C(_07407_),
    .Y(_07409_));
 sky130_fd_sc_hd__a21bo_2 _29033_ (.A1(_07408_),
    .A2(_07409_),
    .B1_N(_07184_),
    .X(_07410_));
 sky130_fd_sc_hd__nand3b_2 _29034_ (.A_N(_07183_),
    .B(_07408_),
    .C(_07409_),
    .Y(_07411_));
 sky130_fd_sc_hd__a22oi_2 _29035_ (.A1(_07389_),
    .A2(_07391_),
    .B1(_07410_),
    .B2(_07411_),
    .Y(_07412_));
 sky130_fd_sc_hd__nand2_2 _29036_ (.A(_07391_),
    .B(_07389_),
    .Y(_07413_));
 sky130_fd_sc_hd__nand2_2 _29037_ (.A(_07410_),
    .B(_07411_),
    .Y(_07414_));
 sky130_fd_sc_hd__nor2_2 _29038_ (.A(_07413_),
    .B(_07414_),
    .Y(_07415_));
 sky130_fd_sc_hd__o21ai_2 _29039_ (.A1(_07223_),
    .A2(_07187_),
    .B1(_07188_),
    .Y(_07416_));
 sky130_fd_sc_hd__o21bai_2 _29040_ (.A1(_07412_),
    .A2(_07415_),
    .B1_N(_07416_),
    .Y(_07417_));
 sky130_fd_sc_hd__nand3b_2 _29041_ (.A_N(_07413_),
    .B(_07411_),
    .C(_07410_),
    .Y(_07418_));
 sky130_fd_sc_hd__nand3b_2 _29042_ (.A_N(_07412_),
    .B(_07418_),
    .C(_07416_),
    .Y(_07419_));
 sky130_fd_sc_hd__nand2_2 _29043_ (.A(_18771_),
    .B(_06546_),
    .Y(_07420_));
 sky130_fd_sc_hd__buf_1 _29044_ (.A(_18775_),
    .X(_07421_));
 sky130_fd_sc_hd__nand2_2 _29045_ (.A(_07421_),
    .B(_05402_),
    .Y(_07422_));
 sky130_fd_sc_hd__xor2_2 _29046_ (.A(_07420_),
    .B(_07422_),
    .X(_07423_));
 sky130_fd_sc_hd__a21oi_2 _29047_ (.A1(_07417_),
    .A2(_07419_),
    .B1(_07423_),
    .Y(_07424_));
 sky130_fd_sc_hd__nand3_2 _29048_ (.A(_07417_),
    .B(_07419_),
    .C(_07423_),
    .Y(_07425_));
 sky130_vsdinv _29049_ (.A(_07425_),
    .Y(_07426_));
 sky130_fd_sc_hd__nand3_2 _29050_ (.A(_07227_),
    .B(_07163_),
    .C(_07228_),
    .Y(_07427_));
 sky130_fd_sc_hd__o21ai_2 _29051_ (.A1(_07424_),
    .A2(_07426_),
    .B1(_07427_),
    .Y(_07428_));
 sky130_fd_sc_hd__a21o_2 _29052_ (.A1(_07417_),
    .A2(_07419_),
    .B1(_07423_),
    .X(_07429_));
 sky130_fd_sc_hd__nand3b_2 _29053_ (.A_N(_07427_),
    .B(_07429_),
    .C(_07425_),
    .Y(_07430_));
 sky130_fd_sc_hd__nand2_2 _29054_ (.A(_07428_),
    .B(_07430_),
    .Y(_07431_));
 sky130_vsdinv _29055_ (.A(_07431_),
    .Y(_07432_));
 sky130_fd_sc_hd__o21bai_2 _29056_ (.A1(_07360_),
    .A2(_07363_),
    .B1_N(_07432_),
    .Y(_07433_));
 sky130_fd_sc_hd__o21bai_2 _29057_ (.A1(_07361_),
    .A2(_07362_),
    .B1_N(_07359_),
    .Y(_07434_));
 sky130_fd_sc_hd__nand3_2 _29058_ (.A(_07353_),
    .B(_07359_),
    .C(_07357_),
    .Y(_07435_));
 sky130_fd_sc_hd__nand3_2 _29059_ (.A(_07434_),
    .B(_07432_),
    .C(_07435_),
    .Y(_07436_));
 sky130_fd_sc_hd__a21oi_2 _29060_ (.A1(_07433_),
    .A2(_07436_),
    .B1(_07238_),
    .Y(_07437_));
 sky130_fd_sc_hd__a21oi_2 _29061_ (.A1(_07434_),
    .A2(_07435_),
    .B1(_07432_),
    .Y(_07438_));
 sky130_fd_sc_hd__nor3_2 _29062_ (.A(_07431_),
    .B(_07360_),
    .C(_07363_),
    .Y(_07439_));
 sky130_fd_sc_hd__nor3_2 _29063_ (.A(_07234_),
    .B(_07438_),
    .C(_07439_),
    .Y(_07440_));
 sky130_fd_sc_hd__a21boi_2 _29064_ (.A1(_07136_),
    .A2(_07131_),
    .B1_N(_07133_),
    .Y(_07441_));
 sky130_fd_sc_hd__o21ai_2 _29065_ (.A1(_07154_),
    .A2(_07157_),
    .B1(_07153_),
    .Y(_07442_));
 sky130_fd_sc_hd__xor2_2 _29066_ (.A(_07441_),
    .B(_07442_),
    .X(_07443_));
 sky130_vsdinv _29067_ (.A(_07443_),
    .Y(_07444_));
 sky130_fd_sc_hd__o21bai_2 _29068_ (.A1(_07437_),
    .A2(_07440_),
    .B1_N(_07444_),
    .Y(_07445_));
 sky130_fd_sc_hd__o21ai_2 _29069_ (.A1(_07438_),
    .A2(_07439_),
    .B1(_07234_),
    .Y(_07446_));
 sky130_fd_sc_hd__nand3_2 _29070_ (.A(_07238_),
    .B(_07433_),
    .C(_07436_),
    .Y(_07447_));
 sky130_fd_sc_hd__nand3_2 _29071_ (.A(_07446_),
    .B(_07444_),
    .C(_07447_),
    .Y(_07448_));
 sky130_fd_sc_hd__o21ai_2 _29072_ (.A1(_07251_),
    .A2(_07235_),
    .B1(_07245_),
    .Y(_07449_));
 sky130_fd_sc_hd__a21oi_2 _29073_ (.A1(_07445_),
    .A2(_07448_),
    .B1(_07449_),
    .Y(_07450_));
 sky130_fd_sc_hd__nand3_2 _29074_ (.A(_07445_),
    .B(_07448_),
    .C(_07449_),
    .Y(_07451_));
 sky130_vsdinv _29075_ (.A(_07451_),
    .Y(_07452_));
 sky130_fd_sc_hd__a21oi_2 _29076_ (.A1(_07026_),
    .A2(_06973_),
    .B1(_07240_),
    .Y(_07453_));
 sky130_fd_sc_hd__o21bai_2 _29077_ (.A1(_07450_),
    .A2(_07452_),
    .B1_N(_07453_),
    .Y(_07454_));
 sky130_fd_sc_hd__a21oi_2 _29078_ (.A1(_07446_),
    .A2(_07447_),
    .B1(_07444_),
    .Y(_07455_));
 sky130_fd_sc_hd__nor3_2 _29079_ (.A(_07443_),
    .B(_07437_),
    .C(_07440_),
    .Y(_07456_));
 sky130_fd_sc_hd__o21bai_2 _29080_ (.A1(_07455_),
    .A2(_07456_),
    .B1_N(_07449_),
    .Y(_07457_));
 sky130_fd_sc_hd__nand3_2 _29081_ (.A(_07457_),
    .B(_07453_),
    .C(_07451_),
    .Y(_07458_));
 sky130_vsdinv _29082_ (.A(_07249_),
    .Y(_07459_));
 sky130_fd_sc_hd__a21o_2 _29083_ (.A1(_07253_),
    .A2(_07255_),
    .B1(_07459_),
    .X(_07460_));
 sky130_fd_sc_hd__a21oi_2 _29084_ (.A1(_07454_),
    .A2(_07458_),
    .B1(_07460_),
    .Y(_07461_));
 sky130_fd_sc_hd__a21oi_2 _29085_ (.A1(_07253_),
    .A2(_07255_),
    .B1(_07459_),
    .Y(_07462_));
 sky130_fd_sc_hd__a21oi_2 _29086_ (.A1(_07457_),
    .A2(_07451_),
    .B1(_07453_),
    .Y(_07463_));
 sky130_vsdinv _29087_ (.A(_07458_),
    .Y(_07464_));
 sky130_fd_sc_hd__nor3_2 _29088_ (.A(_07462_),
    .B(_07463_),
    .C(_07464_),
    .Y(_07465_));
 sky130_fd_sc_hd__nor2_2 _29089_ (.A(_07461_),
    .B(_07465_),
    .Y(_07466_));
 sky130_fd_sc_hd__o21bai_2 _29090_ (.A1(_07258_),
    .A2(_07263_),
    .B1_N(_07260_),
    .Y(_07467_));
 sky130_fd_sc_hd__xor2_2 _29091_ (.A(_07466_),
    .B(_07467_),
    .X(_02638_));
 sky130_fd_sc_hd__buf_1 _29092_ (.A(\pcpi_mul.rs2[17] ),
    .X(_07468_));
 sky130_fd_sc_hd__buf_1 _29093_ (.A(_07468_),
    .X(_07469_));
 sky130_fd_sc_hd__buf_1 _29094_ (.A(_07394_),
    .X(_07470_));
 sky130_fd_sc_hd__a22oi_2 _29095_ (.A1(_07469_),
    .A2(_05540_),
    .B1(_07470_),
    .B2(_05814_),
    .Y(_07471_));
 sky130_fd_sc_hd__buf_1 _29096_ (.A(_07164_),
    .X(_07472_));
 sky130_fd_sc_hd__nand2_2 _29097_ (.A(_07472_),
    .B(_05444_),
    .Y(_07473_));
 sky130_fd_sc_hd__buf_1 _29098_ (.A(_07168_),
    .X(_07474_));
 sky130_fd_sc_hd__nand2_2 _29099_ (.A(_07474_),
    .B(_07403_),
    .Y(_07475_));
 sky130_fd_sc_hd__nor2_2 _29100_ (.A(_07473_),
    .B(_07475_),
    .Y(_07476_));
 sky130_fd_sc_hd__buf_1 _29101_ (.A(_06665_),
    .X(_07477_));
 sky130_fd_sc_hd__and2_2 _29102_ (.A(_07477_),
    .B(_06991_),
    .X(_07478_));
 sky130_fd_sc_hd__o21bai_2 _29103_ (.A1(_07471_),
    .A2(_07476_),
    .B1_N(_07478_),
    .Y(_07479_));
 sky130_fd_sc_hd__buf_1 _29104_ (.A(_07004_),
    .X(_07480_));
 sky130_fd_sc_hd__nand3b_2 _29105_ (.A_N(_07473_),
    .B(_07480_),
    .C(_05733_),
    .Y(_07481_));
 sky130_fd_sc_hd__nand3b_2 _29106_ (.A_N(_07471_),
    .B(_07481_),
    .C(_07478_),
    .Y(_07482_));
 sky130_fd_sc_hd__nor2_2 _29107_ (.A(_07420_),
    .B(_07422_),
    .Y(_07483_));
 sky130_fd_sc_hd__a21oi_2 _29108_ (.A1(_07479_),
    .A2(_07482_),
    .B1(_07483_),
    .Y(_07484_));
 sky130_fd_sc_hd__nand3_2 _29109_ (.A(_07479_),
    .B(_07482_),
    .C(_07483_),
    .Y(_07485_));
 sky130_vsdinv _29110_ (.A(_07485_),
    .Y(_07486_));
 sky130_fd_sc_hd__a21oi_2 _29111_ (.A1(_07397_),
    .A2(_07404_),
    .B1(_07398_),
    .Y(_07487_));
 sky130_vsdinv _29112_ (.A(_07487_),
    .Y(_07488_));
 sky130_fd_sc_hd__o21bai_2 _29113_ (.A1(_07484_),
    .A2(_07486_),
    .B1_N(_07488_),
    .Y(_07489_));
 sky130_fd_sc_hd__o2bb2ai_2 _29114_ (.A1_N(_07482_),
    .A2_N(_07479_),
    .B1(_07420_),
    .B2(_07422_),
    .Y(_07490_));
 sky130_fd_sc_hd__nand3_2 _29115_ (.A(_07490_),
    .B(_07488_),
    .C(_07485_),
    .Y(_07491_));
 sky130_vsdinv _29116_ (.A(_07409_),
    .Y(_07492_));
 sky130_fd_sc_hd__a21o_2 _29117_ (.A1(_07489_),
    .A2(_07491_),
    .B1(_07492_),
    .X(_07493_));
 sky130_fd_sc_hd__nand3_2 _29118_ (.A(_07489_),
    .B(_07492_),
    .C(_07491_),
    .Y(_07494_));
 sky130_fd_sc_hd__buf_1 _29119_ (.A(\pcpi_mul.rs2[14] ),
    .X(_07495_));
 sky130_fd_sc_hd__nand2_2 _29120_ (.A(_07495_),
    .B(_05739_),
    .Y(_07496_));
 sky130_fd_sc_hd__nand2_2 _29121_ (.A(_07200_),
    .B(_05741_),
    .Y(_07497_));
 sky130_fd_sc_hd__nor2_2 _29122_ (.A(_07496_),
    .B(_07497_),
    .Y(_07498_));
 sky130_fd_sc_hd__buf_1 _29123_ (.A(_05727_),
    .X(_07499_));
 sky130_fd_sc_hd__and2_2 _29124_ (.A(_07195_),
    .B(_07499_),
    .X(_07500_));
 sky130_fd_sc_hd__nand2_2 _29125_ (.A(_07496_),
    .B(_07497_),
    .Y(_07501_));
 sky130_fd_sc_hd__nand3b_2 _29126_ (.A_N(_07498_),
    .B(_07500_),
    .C(_07501_),
    .Y(_07502_));
 sky130_fd_sc_hd__buf_1 _29127_ (.A(_07495_),
    .X(_07503_));
 sky130_fd_sc_hd__a22oi_2 _29128_ (.A1(_07503_),
    .A2(_05666_),
    .B1(_07201_),
    .B2(_05838_),
    .Y(_07504_));
 sky130_fd_sc_hd__o21bai_2 _29129_ (.A1(_07504_),
    .A2(_07498_),
    .B1_N(_07500_),
    .Y(_07505_));
 sky130_fd_sc_hd__nand2_2 _29130_ (.A(_07502_),
    .B(_07505_),
    .Y(_07506_));
 sky130_fd_sc_hd__a21oi_2 _29131_ (.A1(_07369_),
    .A2(_07368_),
    .B1(_07367_),
    .Y(_07507_));
 sky130_fd_sc_hd__nand2_2 _29132_ (.A(_07506_),
    .B(_07507_),
    .Y(_07508_));
 sky130_fd_sc_hd__nand3b_2 _29133_ (.A_N(_07507_),
    .B(_07502_),
    .C(_07505_),
    .Y(_07509_));
 sky130_fd_sc_hd__nand2_2 _29134_ (.A(_06810_),
    .B(_07216_),
    .Y(_07510_));
 sky130_fd_sc_hd__nand2_2 _29135_ (.A(_07377_),
    .B(_06068_),
    .Y(_07511_));
 sky130_fd_sc_hd__nor2_2 _29136_ (.A(_07510_),
    .B(_07511_),
    .Y(_07512_));
 sky130_vsdinv _29137_ (.A(_07512_),
    .Y(_07513_));
 sky130_fd_sc_hd__nand2_2 _29138_ (.A(_07510_),
    .B(_07511_),
    .Y(_07514_));
 sky130_fd_sc_hd__buf_1 _29139_ (.A(_06201_),
    .X(_07515_));
 sky130_fd_sc_hd__and2_2 _29140_ (.A(_18822_),
    .B(_07515_),
    .X(_07516_));
 sky130_fd_sc_hd__a21oi_2 _29141_ (.A1(_07513_),
    .A2(_07514_),
    .B1(_07516_),
    .Y(_07517_));
 sky130_fd_sc_hd__nand3b_2 _29142_ (.A_N(_07512_),
    .B(_07516_),
    .C(_07514_),
    .Y(_07518_));
 sky130_vsdinv _29143_ (.A(_07518_),
    .Y(_07519_));
 sky130_fd_sc_hd__nor2_2 _29144_ (.A(_07517_),
    .B(_07519_),
    .Y(_07520_));
 sky130_fd_sc_hd__a21oi_2 _29145_ (.A1(_07508_),
    .A2(_07509_),
    .B1(_07520_),
    .Y(_07521_));
 sky130_fd_sc_hd__nand3_2 _29146_ (.A(_07520_),
    .B(_07508_),
    .C(_07509_),
    .Y(_07522_));
 sky130_fd_sc_hd__and2b_2 _29147_ (.A_N(_07521_),
    .B(_07522_),
    .X(_07523_));
 sky130_fd_sc_hd__a21oi_2 _29148_ (.A1(_07493_),
    .A2(_07494_),
    .B1(_07523_),
    .Y(_07524_));
 sky130_fd_sc_hd__nand3_2 _29149_ (.A(_07493_),
    .B(_07523_),
    .C(_07494_),
    .Y(_07525_));
 sky130_vsdinv _29150_ (.A(_07525_),
    .Y(_07526_));
 sky130_fd_sc_hd__nand2_2 _29151_ (.A(_07418_),
    .B(_07411_),
    .Y(_07527_));
 sky130_fd_sc_hd__o21bai_2 _29152_ (.A1(_07524_),
    .A2(_07526_),
    .B1_N(_07527_),
    .Y(_07528_));
 sky130_fd_sc_hd__a21o_2 _29153_ (.A1(_07493_),
    .A2(_07494_),
    .B1(_07523_),
    .X(_07529_));
 sky130_fd_sc_hd__nand3_2 _29154_ (.A(_07529_),
    .B(_07527_),
    .C(_07525_),
    .Y(_07530_));
 sky130_fd_sc_hd__nand2_2 _29155_ (.A(_07528_),
    .B(_07530_),
    .Y(_07531_));
 sky130_fd_sc_hd__buf_1 _29156_ (.A(\pcpi_mul.rs2[18] ),
    .X(_07532_));
 sky130_fd_sc_hd__buf_1 _29157_ (.A(_07532_),
    .X(_07533_));
 sky130_fd_sc_hd__and2_2 _29158_ (.A(_07533_),
    .B(_05984_),
    .X(_07534_));
 sky130_fd_sc_hd__buf_1 _29159_ (.A(_18769_),
    .X(_07535_));
 sky130_fd_sc_hd__nand2_2 _29160_ (.A(_07535_),
    .B(_05510_),
    .Y(_07536_));
 sky130_fd_sc_hd__buf_1 _29161_ (.A(_18763_),
    .X(_07537_));
 sky130_fd_sc_hd__nand2_2 _29162_ (.A(_07537_),
    .B(_05238_),
    .Y(_07538_));
 sky130_fd_sc_hd__xnor2_2 _29163_ (.A(_07536_),
    .B(_07538_),
    .Y(_07539_));
 sky130_fd_sc_hd__xnor2_2 _29164_ (.A(_07534_),
    .B(_07539_),
    .Y(_07540_));
 sky130_vsdinv _29165_ (.A(_07540_),
    .Y(_07541_));
 sky130_fd_sc_hd__nand2_2 _29166_ (.A(_07531_),
    .B(_07541_),
    .Y(_07542_));
 sky130_fd_sc_hd__nand3_2 _29167_ (.A(_07528_),
    .B(_07540_),
    .C(_07530_),
    .Y(_07543_));
 sky130_fd_sc_hd__a21oi_2 _29168_ (.A1(_07542_),
    .A2(_07543_),
    .B1(_07426_),
    .Y(_07544_));
 sky130_fd_sc_hd__a21oi_2 _29169_ (.A1(_07528_),
    .A2(_07530_),
    .B1(_07540_),
    .Y(_07545_));
 sky130_vsdinv _29170_ (.A(_07543_),
    .Y(_07546_));
 sky130_fd_sc_hd__nor3_2 _29171_ (.A(_07425_),
    .B(_07545_),
    .C(_07546_),
    .Y(_07547_));
 sky130_fd_sc_hd__buf_1 _29172_ (.A(_06880_),
    .X(_07548_));
 sky130_fd_sc_hd__a22oi_2 _29173_ (.A1(_07548_),
    .A2(_06463_),
    .B1(_06889_),
    .B2(_07100_),
    .Y(_07549_));
 sky130_fd_sc_hd__nand2_2 _29174_ (.A(_07058_),
    .B(_06186_),
    .Y(_07550_));
 sky130_fd_sc_hd__buf_1 _29175_ (.A(_07098_),
    .X(_07551_));
 sky130_fd_sc_hd__nand2_2 _29176_ (.A(_05767_),
    .B(_07551_),
    .Y(_07552_));
 sky130_fd_sc_hd__nor2_2 _29177_ (.A(_07550_),
    .B(_07552_),
    .Y(_07553_));
 sky130_fd_sc_hd__and2_2 _29178_ (.A(_18838_),
    .B(_06606_),
    .X(_07554_));
 sky130_fd_sc_hd__o21bai_2 _29179_ (.A1(_07549_),
    .A2(_07553_),
    .B1_N(_07554_),
    .Y(_07555_));
 sky130_fd_sc_hd__buf_1 _29180_ (.A(_18832_),
    .X(_07556_));
 sky130_fd_sc_hd__buf_1 _29181_ (.A(_07551_),
    .X(_07557_));
 sky130_fd_sc_hd__nand3b_2 _29182_ (.A_N(_07550_),
    .B(_07556_),
    .C(_07557_),
    .Y(_07558_));
 sky130_fd_sc_hd__nand2_2 _29183_ (.A(_07550_),
    .B(_07552_),
    .Y(_07559_));
 sky130_fd_sc_hd__nand3_2 _29184_ (.A(_07558_),
    .B(_07554_),
    .C(_07559_),
    .Y(_07560_));
 sky130_fd_sc_hd__nand2_2 _29185_ (.A(_07555_),
    .B(_07560_),
    .Y(_07561_));
 sky130_fd_sc_hd__a21oi_2 _29186_ (.A1(_07380_),
    .A2(_07383_),
    .B1(_07379_),
    .Y(_07562_));
 sky130_fd_sc_hd__nand2_2 _29187_ (.A(_07561_),
    .B(_07562_),
    .Y(_07563_));
 sky130_fd_sc_hd__nand3b_2 _29188_ (.A_N(_07562_),
    .B(_07560_),
    .C(_07555_),
    .Y(_07564_));
 sky130_fd_sc_hd__a21oi_2 _29189_ (.A1(_07273_),
    .A2(_07269_),
    .B1(_07268_),
    .Y(_07565_));
 sky130_vsdinv _29190_ (.A(_07565_),
    .Y(_07566_));
 sky130_fd_sc_hd__a21oi_2 _29191_ (.A1(_07563_),
    .A2(_07564_),
    .B1(_07566_),
    .Y(_07567_));
 sky130_fd_sc_hd__nand3_2 _29192_ (.A(_07563_),
    .B(_07566_),
    .C(_07564_),
    .Y(_07568_));
 sky130_vsdinv _29193_ (.A(_07568_),
    .Y(_07569_));
 sky130_fd_sc_hd__o21ai_2 _29194_ (.A1(_07386_),
    .A2(_07374_),
    .B1(_07388_),
    .Y(_07570_));
 sky130_fd_sc_hd__o21bai_2 _29195_ (.A1(_07567_),
    .A2(_07569_),
    .B1_N(_07570_),
    .Y(_07571_));
 sky130_fd_sc_hd__a21o_2 _29196_ (.A1(_07563_),
    .A2(_07564_),
    .B1(_07566_),
    .X(_07572_));
 sky130_fd_sc_hd__nand3_2 _29197_ (.A(_07572_),
    .B(_07570_),
    .C(_07568_),
    .Y(_07573_));
 sky130_fd_sc_hd__buf_1 _29198_ (.A(_07573_),
    .X(_07574_));
 sky130_fd_sc_hd__a21boi_2 _29199_ (.A1(_07277_),
    .A2(_07283_),
    .B1_N(_07279_),
    .Y(_07575_));
 sky130_vsdinv _29200_ (.A(_07575_),
    .Y(_07576_));
 sky130_fd_sc_hd__a21oi_2 _29201_ (.A1(_07571_),
    .A2(_07574_),
    .B1(_07576_),
    .Y(_07577_));
 sky130_vsdinv _29202_ (.A(_07279_),
    .Y(_07578_));
 sky130_vsdinv _29203_ (.A(_07284_),
    .Y(_07579_));
 sky130_fd_sc_hd__o211a_2 _29204_ (.A1(_07578_),
    .A2(_07579_),
    .B1(_07574_),
    .C1(_07571_),
    .X(_07580_));
 sky130_fd_sc_hd__o21ai_2 _29205_ (.A1(_07291_),
    .A2(_07294_),
    .B1(_07290_),
    .Y(_07581_));
 sky130_fd_sc_hd__o21bai_2 _29206_ (.A1(_07577_),
    .A2(_07580_),
    .B1_N(_07581_),
    .Y(_07582_));
 sky130_fd_sc_hd__nand2_2 _29207_ (.A(_07571_),
    .B(_07573_),
    .Y(_07583_));
 sky130_fd_sc_hd__nand2_2 _29208_ (.A(_07583_),
    .B(_07575_),
    .Y(_07584_));
 sky130_fd_sc_hd__nand3_2 _29209_ (.A(_07571_),
    .B(_07576_),
    .C(_07574_),
    .Y(_07585_));
 sky130_fd_sc_hd__nand3_2 _29210_ (.A(_07584_),
    .B(_07585_),
    .C(_07581_),
    .Y(_07586_));
 sky130_fd_sc_hd__buf_1 _29211_ (.A(_07586_),
    .X(_07587_));
 sky130_fd_sc_hd__nand2_2 _29212_ (.A(_06040_),
    .B(_07306_),
    .Y(_07588_));
 sky130_fd_sc_hd__nand2_2 _29213_ (.A(_05643_),
    .B(_19216_),
    .Y(_07589_));
 sky130_fd_sc_hd__nor2_2 _29214_ (.A(_07588_),
    .B(_07589_),
    .Y(_07590_));
 sky130_fd_sc_hd__buf_1 _29215_ (.A(_19195_),
    .X(_07591_));
 sky130_fd_sc_hd__and2_2 _29216_ (.A(_05516_),
    .B(_07591_),
    .X(_07592_));
 sky130_fd_sc_hd__nand2_2 _29217_ (.A(_07588_),
    .B(_07589_),
    .Y(_07593_));
 sky130_fd_sc_hd__nand3b_2 _29218_ (.A_N(_07590_),
    .B(_07592_),
    .C(_07593_),
    .Y(_07594_));
 sky130_fd_sc_hd__buf_1 _29219_ (.A(_05491_),
    .X(_07595_));
 sky130_fd_sc_hd__a22oi_2 _29220_ (.A1(_07595_),
    .A2(_06924_),
    .B1(_05826_),
    .B2(_06735_),
    .Y(_07596_));
 sky130_fd_sc_hd__o21bai_2 _29221_ (.A1(_07596_),
    .A2(_07590_),
    .B1_N(_07592_),
    .Y(_07597_));
 sky130_fd_sc_hd__a21oi_2 _29222_ (.A1(_07312_),
    .A2(_07311_),
    .B1(_07308_),
    .Y(_07598_));
 sky130_fd_sc_hd__a21bo_2 _29223_ (.A1(_07594_),
    .A2(_07597_),
    .B1_N(_07598_),
    .X(_07599_));
 sky130_fd_sc_hd__nand3b_2 _29224_ (.A_N(_07598_),
    .B(_07594_),
    .C(_07597_),
    .Y(_07600_));
 sky130_fd_sc_hd__nand2_2 _29225_ (.A(_07599_),
    .B(_07600_),
    .Y(_07601_));
 sky130_fd_sc_hd__nand2_2 _29226_ (.A(_05531_),
    .B(_07325_),
    .Y(_07602_));
 sky130_fd_sc_hd__nand2_2 _29227_ (.A(_07323_),
    .B(_07310_),
    .Y(_07603_));
 sky130_fd_sc_hd__xor2_2 _29228_ (.A(_07602_),
    .B(_07603_),
    .X(_07604_));
 sky130_fd_sc_hd__buf_1 _29229_ (.A(_06935_),
    .X(_07605_));
 sky130_fd_sc_hd__buf_1 _29230_ (.A(_07605_),
    .X(_07606_));
 sky130_fd_sc_hd__and2_2 _29231_ (.A(_05459_),
    .B(_07606_),
    .X(_07607_));
 sky130_fd_sc_hd__nand2_2 _29232_ (.A(_07604_),
    .B(_07607_),
    .Y(_07608_));
 sky130_fd_sc_hd__xnor2_2 _29233_ (.A(_07602_),
    .B(_07603_),
    .Y(_07609_));
 sky130_fd_sc_hd__o21ai_2 _29234_ (.A1(_07332_),
    .A2(_19213_),
    .B1(_07609_),
    .Y(_07610_));
 sky130_fd_sc_hd__nand2_2 _29235_ (.A(_07608_),
    .B(_07610_),
    .Y(_07611_));
 sky130_fd_sc_hd__nand2_2 _29236_ (.A(_07601_),
    .B(_07611_),
    .Y(_07612_));
 sky130_fd_sc_hd__nand3b_2 _29237_ (.A_N(_07611_),
    .B(_07600_),
    .C(_07599_),
    .Y(_07613_));
 sky130_fd_sc_hd__a21boi_2 _29238_ (.A1(_07313_),
    .A2(_07316_),
    .B1_N(_07317_),
    .Y(_07614_));
 sky130_fd_sc_hd__o21ai_2 _29239_ (.A1(_07614_),
    .A2(_07335_),
    .B1(_07319_),
    .Y(_07615_));
 sky130_fd_sc_hd__a21o_2 _29240_ (.A1(_07612_),
    .A2(_07613_),
    .B1(_07615_),
    .X(_07616_));
 sky130_fd_sc_hd__nand3_2 _29241_ (.A(_07612_),
    .B(_07613_),
    .C(_07615_),
    .Y(_07617_));
 sky130_fd_sc_hd__nand2_2 _29242_ (.A(_07616_),
    .B(_07617_),
    .Y(_07618_));
 sky130_fd_sc_hd__nor2_2 _29243_ (.A(_07322_),
    .B(_07326_),
    .Y(_07619_));
 sky130_fd_sc_hd__a21oi_2 _29244_ (.A1(_07327_),
    .A2(_07330_),
    .B1(_07619_),
    .Y(_07620_));
 sky130_fd_sc_hd__nand2_2 _29245_ (.A(_07618_),
    .B(_07620_),
    .Y(_07621_));
 sky130_vsdinv _29246_ (.A(_07620_),
    .Y(_07622_));
 sky130_fd_sc_hd__nand3_2 _29247_ (.A(_07616_),
    .B(_07622_),
    .C(_07617_),
    .Y(_07623_));
 sky130_fd_sc_hd__nand2_2 _29248_ (.A(_07621_),
    .B(_07623_),
    .Y(_07624_));
 sky130_fd_sc_hd__buf_1 _29249_ (.A(_07624_),
    .X(_07625_));
 sky130_fd_sc_hd__a21boi_2 _29250_ (.A1(_07582_),
    .A2(_07587_),
    .B1_N(_07625_),
    .Y(_07626_));
 sky130_fd_sc_hd__a21oi_2 _29251_ (.A1(_07584_),
    .A2(_07585_),
    .B1(_07581_),
    .Y(_07627_));
 sky130_vsdinv _29252_ (.A(_07587_),
    .Y(_07628_));
 sky130_fd_sc_hd__nor3_2 _29253_ (.A(_07625_),
    .B(_07627_),
    .C(_07628_),
    .Y(_07629_));
 sky130_vsdinv _29254_ (.A(_07419_),
    .Y(_07630_));
 sky130_fd_sc_hd__o21bai_2 _29255_ (.A1(_07626_),
    .A2(_07629_),
    .B1_N(_07630_),
    .Y(_07631_));
 sky130_fd_sc_hd__nand2_2 _29256_ (.A(_07582_),
    .B(_07586_),
    .Y(_07632_));
 sky130_fd_sc_hd__nand2_2 _29257_ (.A(_07632_),
    .B(_07625_),
    .Y(_07633_));
 sky130_fd_sc_hd__nand3b_2 _29258_ (.A_N(_07624_),
    .B(_07587_),
    .C(_07582_),
    .Y(_07634_));
 sky130_fd_sc_hd__nand3_2 _29259_ (.A(_07633_),
    .B(_07634_),
    .C(_07630_),
    .Y(_07635_));
 sky130_fd_sc_hd__buf_1 _29260_ (.A(_07635_),
    .X(_07636_));
 sky130_fd_sc_hd__o21a_2 _29261_ (.A1(_07348_),
    .A2(_07350_),
    .B1(_07302_),
    .X(_07637_));
 sky130_vsdinv _29262_ (.A(_07637_),
    .Y(_07638_));
 sky130_fd_sc_hd__a21oi_2 _29263_ (.A1(_07631_),
    .A2(_07636_),
    .B1(_07638_),
    .Y(_07639_));
 sky130_fd_sc_hd__a21oi_2 _29264_ (.A1(_07633_),
    .A2(_07634_),
    .B1(_07630_),
    .Y(_07640_));
 sky130_vsdinv _29265_ (.A(_07635_),
    .Y(_07641_));
 sky130_fd_sc_hd__nor3_2 _29266_ (.A(_07637_),
    .B(_07640_),
    .C(_07641_),
    .Y(_07642_));
 sky130_fd_sc_hd__o22ai_2 _29267_ (.A1(_07544_),
    .A2(_07547_),
    .B1(_07639_),
    .B2(_07642_),
    .Y(_07643_));
 sky130_fd_sc_hd__o21bai_2 _29268_ (.A1(_07640_),
    .A2(_07641_),
    .B1_N(_07638_),
    .Y(_07644_));
 sky130_fd_sc_hd__nor2_2 _29269_ (.A(_07544_),
    .B(_07547_),
    .Y(_07645_));
 sky130_fd_sc_hd__nand3_2 _29270_ (.A(_07631_),
    .B(_07638_),
    .C(_07636_),
    .Y(_07646_));
 sky130_fd_sc_hd__nand3_2 _29271_ (.A(_07644_),
    .B(_07645_),
    .C(_07646_),
    .Y(_07647_));
 sky130_fd_sc_hd__nand2_2 _29272_ (.A(_07643_),
    .B(_07647_),
    .Y(_07648_));
 sky130_vsdinv _29273_ (.A(_07430_),
    .Y(_07649_));
 sky130_fd_sc_hd__a31oi_2 _29274_ (.A1(_07434_),
    .A2(_07428_),
    .A3(_07435_),
    .B1(_07649_),
    .Y(_07650_));
 sky130_fd_sc_hd__nand2_2 _29275_ (.A(_07648_),
    .B(_07650_),
    .Y(_07651_));
 sky130_fd_sc_hd__nand2_2 _29276_ (.A(_07436_),
    .B(_07430_),
    .Y(_07652_));
 sky130_fd_sc_hd__nand3_2 _29277_ (.A(_07652_),
    .B(_07647_),
    .C(_07643_),
    .Y(_07653_));
 sky130_fd_sc_hd__buf_1 _29278_ (.A(_07653_),
    .X(_07654_));
 sky130_fd_sc_hd__a21boi_2 _29279_ (.A1(_07339_),
    .A2(_07345_),
    .B1_N(_07340_),
    .Y(_07655_));
 sky130_fd_sc_hd__o21ai_2 _29280_ (.A1(_07358_),
    .A2(_07361_),
    .B1(_07357_),
    .Y(_07656_));
 sky130_fd_sc_hd__xor2_2 _29281_ (.A(_07655_),
    .B(_07656_),
    .X(_07657_));
 sky130_vsdinv _29282_ (.A(_07657_),
    .Y(_07658_));
 sky130_fd_sc_hd__a21oi_2 _29283_ (.A1(_07651_),
    .A2(_07654_),
    .B1(_07658_),
    .Y(_07659_));
 sky130_fd_sc_hd__a21oi_2 _29284_ (.A1(_07643_),
    .A2(_07647_),
    .B1(_07652_),
    .Y(_07660_));
 sky130_fd_sc_hd__nor3b_2 _29285_ (.A(_07657_),
    .B(_07660_),
    .C_N(_07654_),
    .Y(_07661_));
 sky130_fd_sc_hd__o21ai_2 _29286_ (.A1(_07443_),
    .A2(_07437_),
    .B1(_07447_),
    .Y(_07662_));
 sky130_fd_sc_hd__o21bai_2 _29287_ (.A1(_07659_),
    .A2(_07661_),
    .B1_N(_07662_),
    .Y(_07663_));
 sky130_fd_sc_hd__nand2_2 _29288_ (.A(_07651_),
    .B(_07653_),
    .Y(_07664_));
 sky130_fd_sc_hd__nand2_2 _29289_ (.A(_07664_),
    .B(_07657_),
    .Y(_07665_));
 sky130_fd_sc_hd__nand3_2 _29290_ (.A(_07651_),
    .B(_07658_),
    .C(_07654_),
    .Y(_07666_));
 sky130_fd_sc_hd__nand3_2 _29291_ (.A(_07665_),
    .B(_07666_),
    .C(_07662_),
    .Y(_07667_));
 sky130_fd_sc_hd__a21oi_2 _29292_ (.A1(_07233_),
    .A2(_07153_),
    .B1(_07441_),
    .Y(_07668_));
 sky130_fd_sc_hd__a21oi_2 _29293_ (.A1(_07663_),
    .A2(_07667_),
    .B1(_07668_),
    .Y(_07669_));
 sky130_vsdinv _29294_ (.A(_07668_),
    .Y(_07670_));
 sky130_fd_sc_hd__a21oi_2 _29295_ (.A1(_07665_),
    .A2(_07666_),
    .B1(_07662_),
    .Y(_07671_));
 sky130_vsdinv _29296_ (.A(_07667_),
    .Y(_07672_));
 sky130_fd_sc_hd__nor3_2 _29297_ (.A(_07670_),
    .B(_07671_),
    .C(_07672_),
    .Y(_07673_));
 sky130_vsdinv _29298_ (.A(_07453_),
    .Y(_07674_));
 sky130_fd_sc_hd__o21ai_2 _29299_ (.A1(_07674_),
    .A2(_07450_),
    .B1(_07451_),
    .Y(_07675_));
 sky130_fd_sc_hd__o21bai_2 _29300_ (.A1(_07669_),
    .A2(_07673_),
    .B1_N(_07675_),
    .Y(_07676_));
 sky130_fd_sc_hd__o21bai_2 _29301_ (.A1(_07671_),
    .A2(_07672_),
    .B1_N(_07668_),
    .Y(_07677_));
 sky130_fd_sc_hd__nand3_2 _29302_ (.A(_07663_),
    .B(_07668_),
    .C(_07667_),
    .Y(_07678_));
 sky130_fd_sc_hd__nand3_2 _29303_ (.A(_07677_),
    .B(_07678_),
    .C(_07675_),
    .Y(_07679_));
 sky130_fd_sc_hd__nand2_2 _29304_ (.A(_07676_),
    .B(_07679_),
    .Y(_07680_));
 sky130_fd_sc_hd__nand3_2 _29305_ (.A(_06874_),
    .B(_07054_),
    .C(_07055_),
    .Y(_07681_));
 sky130_fd_sc_hd__nand3b_2 _29306_ (.A_N(_07681_),
    .B(_07261_),
    .C(_07466_),
    .Y(_07682_));
 sky130_vsdinv _29307_ (.A(_07682_),
    .Y(_07683_));
 sky130_fd_sc_hd__nand3_2 _29308_ (.A(_07460_),
    .B(_07454_),
    .C(_07458_),
    .Y(_07684_));
 sky130_fd_sc_hd__o21ai_2 _29309_ (.A1(_07259_),
    .A2(_07461_),
    .B1(_07684_),
    .Y(_07685_));
 sky130_fd_sc_hd__a31oi_2 _29310_ (.A1(_07261_),
    .A2(_07466_),
    .A3(_07262_),
    .B1(_07685_),
    .Y(_07686_));
 sky130_fd_sc_hd__a21bo_2 _29311_ (.A1(_06878_),
    .A2(_07683_),
    .B1_N(_07686_),
    .X(_07687_));
 sky130_fd_sc_hd__xnor2_2 _29312_ (.A(_07680_),
    .B(_07687_),
    .Y(_02639_));
 sky130_fd_sc_hd__buf_1 _29313_ (.A(_06452_),
    .X(_07688_));
 sky130_fd_sc_hd__a22oi_2 _29314_ (.A1(_06881_),
    .A2(_19237_),
    .B1(_05992_),
    .B2(_07688_),
    .Y(_07689_));
 sky130_fd_sc_hd__buf_1 _29315_ (.A(_07098_),
    .X(_07690_));
 sky130_fd_sc_hd__nand2_2 _29316_ (.A(_18828_),
    .B(_07690_),
    .Y(_07691_));
 sky130_fd_sc_hd__nand2_2 _29317_ (.A(_06226_),
    .B(_06607_),
    .Y(_07692_));
 sky130_fd_sc_hd__nor2_2 _29318_ (.A(_07691_),
    .B(_07692_),
    .Y(_07693_));
 sky130_fd_sc_hd__buf_1 _29319_ (.A(_19224_),
    .X(_07694_));
 sky130_fd_sc_hd__and2_2 _29320_ (.A(_06100_),
    .B(_07694_),
    .X(_07695_));
 sky130_fd_sc_hd__o21bai_2 _29321_ (.A1(_07689_),
    .A2(_07693_),
    .B1_N(_07695_),
    .Y(_07696_));
 sky130_fd_sc_hd__buf_1 _29322_ (.A(_05872_),
    .X(_07697_));
 sky130_fd_sc_hd__buf_1 _29323_ (.A(_19230_),
    .X(_07698_));
 sky130_fd_sc_hd__buf_1 _29324_ (.A(_07698_),
    .X(_07699_));
 sky130_fd_sc_hd__nand3b_2 _29325_ (.A_N(_07691_),
    .B(_07697_),
    .C(_07699_),
    .Y(_07700_));
 sky130_fd_sc_hd__nand3b_2 _29326_ (.A_N(_07689_),
    .B(_07700_),
    .C(_07695_),
    .Y(_07701_));
 sky130_fd_sc_hd__nand2_2 _29327_ (.A(_07696_),
    .B(_07701_),
    .Y(_07702_));
 sky130_fd_sc_hd__a21oi_2 _29328_ (.A1(_07514_),
    .A2(_07516_),
    .B1(_07512_),
    .Y(_07703_));
 sky130_fd_sc_hd__nand2_2 _29329_ (.A(_07702_),
    .B(_07703_),
    .Y(_07704_));
 sky130_fd_sc_hd__nand3b_2 _29330_ (.A_N(_07703_),
    .B(_07701_),
    .C(_07696_),
    .Y(_07705_));
 sky130_fd_sc_hd__buf_1 _29331_ (.A(_07705_),
    .X(_07706_));
 sky130_fd_sc_hd__a21oi_2 _29332_ (.A1(_07559_),
    .A2(_07554_),
    .B1(_07553_),
    .Y(_07707_));
 sky130_vsdinv _29333_ (.A(_07707_),
    .Y(_07708_));
 sky130_fd_sc_hd__a21oi_2 _29334_ (.A1(_07704_),
    .A2(_07706_),
    .B1(_07708_),
    .Y(_07709_));
 sky130_fd_sc_hd__nand3_2 _29335_ (.A(_07704_),
    .B(_07708_),
    .C(_07705_),
    .Y(_07710_));
 sky130_vsdinv _29336_ (.A(_07710_),
    .Y(_07711_));
 sky130_vsdinv _29337_ (.A(_07509_),
    .Y(_07712_));
 sky130_fd_sc_hd__a21oi_2 _29338_ (.A1(_07520_),
    .A2(_07508_),
    .B1(_07712_),
    .Y(_07713_));
 sky130_fd_sc_hd__o21ai_2 _29339_ (.A1(_07709_),
    .A2(_07711_),
    .B1(_07713_),
    .Y(_07714_));
 sky130_fd_sc_hd__a21o_2 _29340_ (.A1(_07520_),
    .A2(_07508_),
    .B1(_07712_),
    .X(_07715_));
 sky130_fd_sc_hd__a21o_2 _29341_ (.A1(_07704_),
    .A2(_07706_),
    .B1(_07708_),
    .X(_07716_));
 sky130_fd_sc_hd__nand3_2 _29342_ (.A(_07715_),
    .B(_07716_),
    .C(_07710_),
    .Y(_07717_));
 sky130_fd_sc_hd__a21boi_2 _29343_ (.A1(_07563_),
    .A2(_07566_),
    .B1_N(_07564_),
    .Y(_07718_));
 sky130_vsdinv _29344_ (.A(_07718_),
    .Y(_07719_));
 sky130_fd_sc_hd__a21oi_2 _29345_ (.A1(_07714_),
    .A2(_07717_),
    .B1(_07719_),
    .Y(_07720_));
 sky130_fd_sc_hd__nand3_2 _29346_ (.A(_07714_),
    .B(_07719_),
    .C(_07717_),
    .Y(_07721_));
 sky130_vsdinv _29347_ (.A(_07721_),
    .Y(_07722_));
 sky130_fd_sc_hd__a21oi_2 _29348_ (.A1(_07572_),
    .A2(_07568_),
    .B1(_07570_),
    .Y(_07723_));
 sky130_fd_sc_hd__o21ai_2 _29349_ (.A1(_07575_),
    .A2(_07723_),
    .B1(_07574_),
    .Y(_07724_));
 sky130_fd_sc_hd__o21bai_2 _29350_ (.A1(_07720_),
    .A2(_07722_),
    .B1_N(_07724_),
    .Y(_07725_));
 sky130_fd_sc_hd__a21oi_2 _29351_ (.A1(_07716_),
    .A2(_07710_),
    .B1(_07715_),
    .Y(_07726_));
 sky130_fd_sc_hd__nor3_2 _29352_ (.A(_07709_),
    .B(_07713_),
    .C(_07711_),
    .Y(_07727_));
 sky130_fd_sc_hd__o21bai_2 _29353_ (.A1(_07726_),
    .A2(_07727_),
    .B1_N(_07719_),
    .Y(_07728_));
 sky130_fd_sc_hd__nand3_2 _29354_ (.A(_07728_),
    .B(_07721_),
    .C(_07724_),
    .Y(_07729_));
 sky130_fd_sc_hd__nand2_2 _29355_ (.A(_05496_),
    .B(_07115_),
    .Y(_07730_));
 sky130_fd_sc_hd__nand2_2 _29356_ (.A(_05637_),
    .B(_06936_),
    .Y(_07731_));
 sky130_fd_sc_hd__nor2_2 _29357_ (.A(_07730_),
    .B(_07731_),
    .Y(_07732_));
 sky130_fd_sc_hd__buf_1 _29358_ (.A(\pcpi_mul.rs1[21] ),
    .X(_07733_));
 sky130_fd_sc_hd__and2_2 _29359_ (.A(_05647_),
    .B(_07733_),
    .X(_07734_));
 sky130_fd_sc_hd__nand2_2 _29360_ (.A(_07730_),
    .B(_07731_),
    .Y(_07735_));
 sky130_fd_sc_hd__nand3b_2 _29361_ (.A_N(_07732_),
    .B(_07734_),
    .C(_07735_),
    .Y(_07736_));
 sky130_fd_sc_hd__buf_1 _29362_ (.A(_19211_),
    .X(_07737_));
 sky130_fd_sc_hd__a22oi_2 _29363_ (.A1(_05634_),
    .A2(_07116_),
    .B1(_05939_),
    .B2(_07737_),
    .Y(_07738_));
 sky130_fd_sc_hd__o21bai_2 _29364_ (.A1(_07738_),
    .A2(_07732_),
    .B1_N(_07734_),
    .Y(_07739_));
 sky130_fd_sc_hd__a21oi_2 _29365_ (.A1(_07593_),
    .A2(_07592_),
    .B1(_07590_),
    .Y(_07740_));
 sky130_fd_sc_hd__a21bo_2 _29366_ (.A1(_07736_),
    .A2(_07739_),
    .B1_N(_07740_),
    .X(_07741_));
 sky130_fd_sc_hd__nand3b_2 _29367_ (.A_N(_07740_),
    .B(_07736_),
    .C(_07739_),
    .Y(_07742_));
 sky130_fd_sc_hd__buf_1 _29368_ (.A(\pcpi_mul.rs1[19] ),
    .X(_07743_));
 sky130_fd_sc_hd__nand2_2 _29369_ (.A(_05661_),
    .B(_07743_),
    .Y(_07744_));
 sky130_fd_sc_hd__buf_1 _29370_ (.A(\pcpi_mul.rs1[20] ),
    .X(_07745_));
 sky130_fd_sc_hd__nand2_2 _29371_ (.A(_05535_),
    .B(_07745_),
    .Y(_07746_));
 sky130_fd_sc_hd__xor2_2 _29372_ (.A(_07744_),
    .B(_07746_),
    .X(_07747_));
 sky130_fd_sc_hd__buf_1 _29373_ (.A(\pcpi_mul.rs1[18] ),
    .X(_07748_));
 sky130_fd_sc_hd__and2_2 _29374_ (.A(_05458_),
    .B(_07748_),
    .X(_07749_));
 sky130_fd_sc_hd__nand2_2 _29375_ (.A(_07747_),
    .B(_07749_),
    .Y(_07750_));
 sky130_fd_sc_hd__buf_1 _29376_ (.A(_07743_),
    .X(_07751_));
 sky130_fd_sc_hd__buf_1 _29377_ (.A(_07745_),
    .X(_07752_));
 sky130_fd_sc_hd__a22oi_2 _29378_ (.A1(_05662_),
    .A2(_07751_),
    .B1(_18872_),
    .B2(_07752_),
    .Y(_07753_));
 sky130_fd_sc_hd__nor2_2 _29379_ (.A(_07744_),
    .B(_07746_),
    .Y(_07754_));
 sky130_fd_sc_hd__o21bai_2 _29380_ (.A1(_07753_),
    .A2(_07754_),
    .B1_N(_07749_),
    .Y(_07755_));
 sky130_fd_sc_hd__nand2_2 _29381_ (.A(_07750_),
    .B(_07755_),
    .Y(_07756_));
 sky130_fd_sc_hd__a21boi_2 _29382_ (.A1(_07741_),
    .A2(_07742_),
    .B1_N(_07756_),
    .Y(_07757_));
 sky130_fd_sc_hd__nand3b_2 _29383_ (.A_N(_07756_),
    .B(_07742_),
    .C(_07741_),
    .Y(_07758_));
 sky130_vsdinv _29384_ (.A(_07758_),
    .Y(_07759_));
 sky130_fd_sc_hd__a21boi_2 _29385_ (.A1(_07594_),
    .A2(_07597_),
    .B1_N(_07598_),
    .Y(_07760_));
 sky130_fd_sc_hd__o21ai_2 _29386_ (.A1(_07760_),
    .A2(_07611_),
    .B1(_07600_),
    .Y(_07761_));
 sky130_fd_sc_hd__o21bai_2 _29387_ (.A1(_07757_),
    .A2(_07759_),
    .B1_N(_07761_),
    .Y(_07762_));
 sky130_fd_sc_hd__nand3b_2 _29388_ (.A_N(_07757_),
    .B(_07758_),
    .C(_07761_),
    .Y(_07763_));
 sky130_fd_sc_hd__nand2_2 _29389_ (.A(_07762_),
    .B(_07763_),
    .Y(_07764_));
 sky130_fd_sc_hd__o21a_2 _29390_ (.A1(_07602_),
    .A2(_07603_),
    .B1(_07608_),
    .X(_07765_));
 sky130_fd_sc_hd__nand2_2 _29391_ (.A(_07764_),
    .B(_07765_),
    .Y(_07766_));
 sky130_fd_sc_hd__nand3b_2 _29392_ (.A_N(_07765_),
    .B(_07762_),
    .C(_07763_),
    .Y(_07767_));
 sky130_fd_sc_hd__nand2_2 _29393_ (.A(_07766_),
    .B(_07767_),
    .Y(_07768_));
 sky130_fd_sc_hd__a21boi_2 _29394_ (.A1(_07725_),
    .A2(_07729_),
    .B1_N(_07768_),
    .Y(_07769_));
 sky130_fd_sc_hd__buf_1 _29395_ (.A(_07768_),
    .X(_07770_));
 sky130_fd_sc_hd__a21oi_2 _29396_ (.A1(_07728_),
    .A2(_07721_),
    .B1(_07724_),
    .Y(_07771_));
 sky130_vsdinv _29397_ (.A(_07729_),
    .Y(_07772_));
 sky130_fd_sc_hd__nor3_2 _29398_ (.A(_07770_),
    .B(_07771_),
    .C(_07772_),
    .Y(_07773_));
 sky130_vsdinv _29399_ (.A(_07530_),
    .Y(_07774_));
 sky130_fd_sc_hd__o21bai_2 _29400_ (.A1(_07769_),
    .A2(_07773_),
    .B1_N(_07774_),
    .Y(_07775_));
 sky130_fd_sc_hd__buf_1 _29401_ (.A(_07775_),
    .X(_07776_));
 sky130_fd_sc_hd__o21ai_2 _29402_ (.A1(_07771_),
    .A2(_07772_),
    .B1(_07770_),
    .Y(_07777_));
 sky130_fd_sc_hd__nand3b_2 _29403_ (.A_N(_07770_),
    .B(_07729_),
    .C(_07725_),
    .Y(_07778_));
 sky130_fd_sc_hd__nand3_2 _29404_ (.A(_07777_),
    .B(_07774_),
    .C(_07778_),
    .Y(_07779_));
 sky130_fd_sc_hd__buf_1 _29405_ (.A(_07779_),
    .X(_07780_));
 sky130_fd_sc_hd__o21a_2 _29406_ (.A1(_07625_),
    .A2(_07627_),
    .B1(_07587_),
    .X(_07781_));
 sky130_vsdinv _29407_ (.A(_07781_),
    .Y(_07782_));
 sky130_fd_sc_hd__a21oi_2 _29408_ (.A1(_07776_),
    .A2(_07780_),
    .B1(_07782_),
    .Y(_07783_));
 sky130_fd_sc_hd__o211a_2 _29409_ (.A1(_07628_),
    .A2(_07629_),
    .B1(_07779_),
    .C1(_07776_),
    .X(_07784_));
 sky130_fd_sc_hd__buf_1 _29410_ (.A(\pcpi_mul.rs2[17] ),
    .X(_07785_));
 sky130_fd_sc_hd__buf_1 _29411_ (.A(_07785_),
    .X(_07786_));
 sky130_fd_sc_hd__buf_1 _29412_ (.A(_07167_),
    .X(_07787_));
 sky130_fd_sc_hd__buf_1 _29413_ (.A(_07787_),
    .X(_07788_));
 sky130_fd_sc_hd__a22oi_2 _29414_ (.A1(_07786_),
    .A2(_05533_),
    .B1(_07788_),
    .B2(_06820_),
    .Y(_07789_));
 sky130_fd_sc_hd__buf_1 _29415_ (.A(_19281_),
    .X(_07790_));
 sky130_fd_sc_hd__and4_2 _29416_ (.A(_18780_),
    .B(_18785_),
    .C(_06991_),
    .D(_07790_),
    .X(_07791_));
 sky130_fd_sc_hd__and2_2 _29417_ (.A(_07012_),
    .B(_19272_),
    .X(_07792_));
 sky130_fd_sc_hd__o21bai_2 _29418_ (.A1(_07789_),
    .A2(_07791_),
    .B1_N(_07792_),
    .Y(_07793_));
 sky130_fd_sc_hd__buf_1 _29419_ (.A(_19281_),
    .X(_07794_));
 sky130_fd_sc_hd__nand2_2 _29420_ (.A(_07472_),
    .B(_07794_),
    .Y(_07795_));
 sky130_fd_sc_hd__nand3b_2 _29421_ (.A_N(_07795_),
    .B(_07480_),
    .C(_06102_),
    .Y(_07796_));
 sky130_fd_sc_hd__nand3b_2 _29422_ (.A_N(_07789_),
    .B(_07796_),
    .C(_07792_),
    .Y(_07797_));
 sky130_fd_sc_hd__nand2_2 _29423_ (.A(_07793_),
    .B(_07797_),
    .Y(_07798_));
 sky130_fd_sc_hd__nand2_2 _29424_ (.A(_07536_),
    .B(_07538_),
    .Y(_07799_));
 sky130_fd_sc_hd__nor2_2 _29425_ (.A(_07536_),
    .B(_07538_),
    .Y(_07800_));
 sky130_fd_sc_hd__a21oi_2 _29426_ (.A1(_07799_),
    .A2(_07534_),
    .B1(_07800_),
    .Y(_07801_));
 sky130_fd_sc_hd__nand2_2 _29427_ (.A(_07798_),
    .B(_07801_),
    .Y(_07802_));
 sky130_fd_sc_hd__nand3b_2 _29428_ (.A_N(_07801_),
    .B(_07793_),
    .C(_07797_),
    .Y(_07803_));
 sky130_fd_sc_hd__nand2_2 _29429_ (.A(_07802_),
    .B(_07803_),
    .Y(_07804_));
 sky130_fd_sc_hd__o31a_2 _29430_ (.A1(_18792_),
    .A2(_19278_),
    .A3(_07471_),
    .B1(_07481_),
    .X(_07805_));
 sky130_fd_sc_hd__nand2_2 _29431_ (.A(_07804_),
    .B(_07805_),
    .Y(_07806_));
 sky130_vsdinv _29432_ (.A(_07805_),
    .Y(_07807_));
 sky130_fd_sc_hd__nand3_2 _29433_ (.A(_07802_),
    .B(_07807_),
    .C(_07803_),
    .Y(_07808_));
 sky130_fd_sc_hd__o21ai_2 _29434_ (.A1(_07487_),
    .A2(_07484_),
    .B1(_07485_),
    .Y(_07809_));
 sky130_fd_sc_hd__a21oi_2 _29435_ (.A1(_07806_),
    .A2(_07808_),
    .B1(_07809_),
    .Y(_07810_));
 sky130_fd_sc_hd__nand3_2 _29436_ (.A(_07806_),
    .B(_07808_),
    .C(_07809_),
    .Y(_07811_));
 sky130_vsdinv _29437_ (.A(_07811_),
    .Y(_07812_));
 sky130_fd_sc_hd__nand2_2 _29438_ (.A(_06811_),
    .B(_06069_),
    .Y(_07813_));
 sky130_fd_sc_hd__nand2_2 _29439_ (.A(_06812_),
    .B(_06589_),
    .Y(_07814_));
 sky130_fd_sc_hd__nand2_2 _29440_ (.A(_07813_),
    .B(_07814_),
    .Y(_07815_));
 sky130_fd_sc_hd__nor2_2 _29441_ (.A(_07813_),
    .B(_07814_),
    .Y(_07816_));
 sky130_vsdinv _29442_ (.A(_07816_),
    .Y(_07817_));
 sky130_fd_sc_hd__buf_1 _29443_ (.A(_18823_),
    .X(_07818_));
 sky130_fd_sc_hd__o2bb2ai_2 _29444_ (.A1_N(_07815_),
    .A2_N(_07817_),
    .B1(_07818_),
    .B2(_19244_),
    .Y(_07819_));
 sky130_fd_sc_hd__and2_2 _29445_ (.A(_06680_),
    .B(_06729_),
    .X(_07820_));
 sky130_fd_sc_hd__nand3b_2 _29446_ (.A_N(_07816_),
    .B(_07820_),
    .C(_07815_),
    .Y(_07821_));
 sky130_fd_sc_hd__nand2_2 _29447_ (.A(_07819_),
    .B(_07821_),
    .Y(_07822_));
 sky130_fd_sc_hd__nand2_2 _29448_ (.A(_07503_),
    .B(_06180_),
    .Y(_07823_));
 sky130_fd_sc_hd__buf_1 _29449_ (.A(_07192_),
    .X(_07824_));
 sky130_fd_sc_hd__nand2_2 _29450_ (.A(_07824_),
    .B(_06075_),
    .Y(_07825_));
 sky130_fd_sc_hd__nor2_2 _29451_ (.A(_07823_),
    .B(_07825_),
    .Y(_07826_));
 sky130_fd_sc_hd__and2_2 _29452_ (.A(_06275_),
    .B(_06343_),
    .X(_07827_));
 sky130_fd_sc_hd__nand2_2 _29453_ (.A(_07823_),
    .B(_07825_),
    .Y(_07828_));
 sky130_fd_sc_hd__nand3b_2 _29454_ (.A_N(_07826_),
    .B(_07827_),
    .C(_07828_),
    .Y(_07829_));
 sky130_fd_sc_hd__a22oi_2 _29455_ (.A1(_06535_),
    .A2(_06486_),
    .B1(_06394_),
    .B2(_05848_),
    .Y(_07830_));
 sky130_fd_sc_hd__o21bai_2 _29456_ (.A1(_07830_),
    .A2(_07826_),
    .B1_N(_07827_),
    .Y(_07831_));
 sky130_fd_sc_hd__a21oi_2 _29457_ (.A1(_07501_),
    .A2(_07500_),
    .B1(_07498_),
    .Y(_07832_));
 sky130_fd_sc_hd__a21bo_2 _29458_ (.A1(_07829_),
    .A2(_07831_),
    .B1_N(_07832_),
    .X(_07833_));
 sky130_fd_sc_hd__nand3b_2 _29459_ (.A_N(_07832_),
    .B(_07829_),
    .C(_07831_),
    .Y(_07834_));
 sky130_fd_sc_hd__nand2_2 _29460_ (.A(_07833_),
    .B(_07834_),
    .Y(_07835_));
 sky130_fd_sc_hd__xnor2_2 _29461_ (.A(_07822_),
    .B(_07835_),
    .Y(_07836_));
 sky130_fd_sc_hd__o21ai_2 _29462_ (.A1(_07810_),
    .A2(_07812_),
    .B1(_07836_),
    .Y(_07837_));
 sky130_fd_sc_hd__xor2_2 _29463_ (.A(_07822_),
    .B(_07835_),
    .X(_07838_));
 sky130_fd_sc_hd__nand3b_2 _29464_ (.A_N(_07810_),
    .B(_07838_),
    .C(_07811_),
    .Y(_07839_));
 sky130_fd_sc_hd__nand2_2 _29465_ (.A(_07525_),
    .B(_07494_),
    .Y(_07840_));
 sky130_fd_sc_hd__a21oi_2 _29466_ (.A1(_07837_),
    .A2(_07839_),
    .B1(_07840_),
    .Y(_07841_));
 sky130_fd_sc_hd__nand3_2 _29467_ (.A(_07840_),
    .B(_07837_),
    .C(_07839_),
    .Y(_07842_));
 sky130_vsdinv _29468_ (.A(_07842_),
    .Y(_07843_));
 sky130_fd_sc_hd__buf_1 _29469_ (.A(\pcpi_mul.rs2[21] ),
    .X(_07844_));
 sky130_fd_sc_hd__buf_1 _29470_ (.A(_07844_),
    .X(_07845_));
 sky130_fd_sc_hd__buf_1 _29471_ (.A(_07845_),
    .X(_07846_));
 sky130_fd_sc_hd__buf_1 _29472_ (.A(_07846_),
    .X(_07847_));
 sky130_fd_sc_hd__and2_2 _29473_ (.A(_07847_),
    .B(_05589_),
    .X(_07848_));
 sky130_fd_sc_hd__and2_2 _29474_ (.A(_07533_),
    .B(_06827_),
    .X(_07849_));
 sky130_fd_sc_hd__buf_1 _29475_ (.A(\pcpi_mul.rs2[20] ),
    .X(_07850_));
 sky130_fd_sc_hd__buf_1 _29476_ (.A(_07850_),
    .X(_07851_));
 sky130_fd_sc_hd__nand2_2 _29477_ (.A(_07851_),
    .B(_05424_),
    .Y(_07852_));
 sky130_fd_sc_hd__buf_1 _29478_ (.A(_18769_),
    .X(_07853_));
 sky130_fd_sc_hd__nand2_2 _29479_ (.A(_07853_),
    .B(_05431_),
    .Y(_07854_));
 sky130_fd_sc_hd__xnor2_2 _29480_ (.A(_07852_),
    .B(_07854_),
    .Y(_07855_));
 sky130_fd_sc_hd__xor2_2 _29481_ (.A(_07849_),
    .B(_07855_),
    .X(_07856_));
 sky130_fd_sc_hd__xnor2_2 _29482_ (.A(_07848_),
    .B(_07856_),
    .Y(_07857_));
 sky130_fd_sc_hd__o21bai_2 _29483_ (.A1(_07841_),
    .A2(_07843_),
    .B1_N(_07857_),
    .Y(_07858_));
 sky130_fd_sc_hd__a21o_2 _29484_ (.A1(_07837_),
    .A2(_07839_),
    .B1(_07840_),
    .X(_07859_));
 sky130_fd_sc_hd__nand3_2 _29485_ (.A(_07859_),
    .B(_07857_),
    .C(_07842_),
    .Y(_07860_));
 sky130_fd_sc_hd__a21oi_2 _29486_ (.A1(_07858_),
    .A2(_07860_),
    .B1(_07546_),
    .Y(_07861_));
 sky130_fd_sc_hd__a21oi_2 _29487_ (.A1(_07859_),
    .A2(_07842_),
    .B1(_07857_),
    .Y(_07862_));
 sky130_vsdinv _29488_ (.A(_07860_),
    .Y(_07863_));
 sky130_fd_sc_hd__nor3_2 _29489_ (.A(_07543_),
    .B(_07862_),
    .C(_07863_),
    .Y(_07864_));
 sky130_fd_sc_hd__nor2_2 _29490_ (.A(_07861_),
    .B(_07864_),
    .Y(_07865_));
 sky130_fd_sc_hd__o21bai_2 _29491_ (.A1(_07783_),
    .A2(_07784_),
    .B1_N(_07865_),
    .Y(_07866_));
 sky130_fd_sc_hd__nand2_2 _29492_ (.A(_07775_),
    .B(_07779_),
    .Y(_07867_));
 sky130_fd_sc_hd__nand2_2 _29493_ (.A(_07867_),
    .B(_07781_),
    .Y(_07868_));
 sky130_fd_sc_hd__nand3_2 _29494_ (.A(_07776_),
    .B(_07782_),
    .C(_07780_),
    .Y(_07869_));
 sky130_fd_sc_hd__nand3_2 _29495_ (.A(_07868_),
    .B(_07865_),
    .C(_07869_),
    .Y(_07870_));
 sky130_fd_sc_hd__nand2_2 _29496_ (.A(_07866_),
    .B(_07870_),
    .Y(_07871_));
 sky130_fd_sc_hd__a31oi_2 _29497_ (.A1(_07644_),
    .A2(_07645_),
    .A3(_07646_),
    .B1(_07547_),
    .Y(_07872_));
 sky130_fd_sc_hd__nand2_2 _29498_ (.A(_07871_),
    .B(_07872_),
    .Y(_07873_));
 sky130_vsdinv _29499_ (.A(_07547_),
    .Y(_07874_));
 sky130_fd_sc_hd__nand2_2 _29500_ (.A(_07647_),
    .B(_07874_),
    .Y(_07875_));
 sky130_fd_sc_hd__nand3_2 _29501_ (.A(_07875_),
    .B(_07866_),
    .C(_07870_),
    .Y(_07876_));
 sky130_fd_sc_hd__buf_1 _29502_ (.A(_07876_),
    .X(_07877_));
 sky130_fd_sc_hd__a21boi_2 _29503_ (.A1(_07616_),
    .A2(_07622_),
    .B1_N(_07617_),
    .Y(_07878_));
 sky130_fd_sc_hd__o21ai_2 _29504_ (.A1(_07637_),
    .A2(_07640_),
    .B1(_07636_),
    .Y(_07879_));
 sky130_fd_sc_hd__xnor2_2 _29505_ (.A(_07878_),
    .B(_07879_),
    .Y(_07880_));
 sky130_fd_sc_hd__a21oi_2 _29506_ (.A1(_07873_),
    .A2(_07877_),
    .B1(_07880_),
    .Y(_07881_));
 sky130_vsdinv _29507_ (.A(_07880_),
    .Y(_07882_));
 sky130_fd_sc_hd__a21oi_2 _29508_ (.A1(_07866_),
    .A2(_07870_),
    .B1(_07875_),
    .Y(_07883_));
 sky130_fd_sc_hd__nor3b_2 _29509_ (.A(_07882_),
    .B(_07883_),
    .C_N(_07877_),
    .Y(_07884_));
 sky130_fd_sc_hd__o21ai_2 _29510_ (.A1(_07657_),
    .A2(_07660_),
    .B1(_07654_),
    .Y(_07885_));
 sky130_fd_sc_hd__o21bai_2 _29511_ (.A1(_07881_),
    .A2(_07884_),
    .B1_N(_07885_),
    .Y(_07886_));
 sky130_fd_sc_hd__nand2_2 _29512_ (.A(_07873_),
    .B(_07876_),
    .Y(_07887_));
 sky130_fd_sc_hd__nand2_2 _29513_ (.A(_07887_),
    .B(_07882_),
    .Y(_07888_));
 sky130_fd_sc_hd__nand3_2 _29514_ (.A(_07873_),
    .B(_07880_),
    .C(_07877_),
    .Y(_07889_));
 sky130_fd_sc_hd__nand3_2 _29515_ (.A(_07888_),
    .B(_07889_),
    .C(_07885_),
    .Y(_07890_));
 sky130_fd_sc_hd__buf_1 _29516_ (.A(_07890_),
    .X(_07891_));
 sky130_fd_sc_hd__a21oi_2 _29517_ (.A1(_07435_),
    .A2(_07357_),
    .B1(_07655_),
    .Y(_07892_));
 sky130_fd_sc_hd__buf_1 _29518_ (.A(_07892_),
    .X(_07893_));
 sky130_fd_sc_hd__a21oi_2 _29519_ (.A1(_07886_),
    .A2(_07891_),
    .B1(_07893_),
    .Y(_07894_));
 sky130_vsdinv _29520_ (.A(_07892_),
    .Y(_07895_));
 sky130_fd_sc_hd__a21oi_2 _29521_ (.A1(_07888_),
    .A2(_07889_),
    .B1(_07885_),
    .Y(_07896_));
 sky130_vsdinv _29522_ (.A(_07890_),
    .Y(_07897_));
 sky130_fd_sc_hd__nor3_2 _29523_ (.A(_07895_),
    .B(_07896_),
    .C(_07897_),
    .Y(_07898_));
 sky130_fd_sc_hd__o21ai_2 _29524_ (.A1(_07670_),
    .A2(_07671_),
    .B1(_07667_),
    .Y(_07899_));
 sky130_fd_sc_hd__o21bai_2 _29525_ (.A1(_07894_),
    .A2(_07898_),
    .B1_N(_07899_),
    .Y(_07900_));
 sky130_fd_sc_hd__o21bai_2 _29526_ (.A1(_07896_),
    .A2(_07897_),
    .B1_N(_07893_),
    .Y(_07901_));
 sky130_fd_sc_hd__nand3_2 _29527_ (.A(_07886_),
    .B(_07893_),
    .C(_07891_),
    .Y(_07902_));
 sky130_fd_sc_hd__nand3_2 _29528_ (.A(_07901_),
    .B(_07899_),
    .C(_07902_),
    .Y(_07903_));
 sky130_fd_sc_hd__nand2_2 _29529_ (.A(_07900_),
    .B(_07903_),
    .Y(_07904_));
 sky130_fd_sc_hd__a21boi_2 _29530_ (.A1(_07687_),
    .A2(_07676_),
    .B1_N(_07679_),
    .Y(_07905_));
 sky130_fd_sc_hd__xor2_2 _29531_ (.A(_07904_),
    .B(_07905_),
    .X(_02640_));
 sky130_fd_sc_hd__buf_1 _29532_ (.A(_07694_),
    .X(_07906_));
 sky130_fd_sc_hd__a22oi_2 _29533_ (.A1(_06105_),
    .A2(_07699_),
    .B1(_05873_),
    .B2(_07906_),
    .Y(_07907_));
 sky130_fd_sc_hd__nand2_2 _29534_ (.A(_06224_),
    .B(_06453_),
    .Y(_07908_));
 sky130_fd_sc_hd__nand2_2 _29535_ (.A(_06890_),
    .B(_06596_),
    .Y(_07909_));
 sky130_fd_sc_hd__nor2_2 _29536_ (.A(_07908_),
    .B(_07909_),
    .Y(_07910_));
 sky130_fd_sc_hd__and2_2 _29537_ (.A(_06771_),
    .B(_07116_),
    .X(_07911_));
 sky130_fd_sc_hd__o21bai_2 _29538_ (.A1(_07907_),
    .A2(_07910_),
    .B1_N(_07911_),
    .Y(_07912_));
 sky130_fd_sc_hd__buf_1 _29539_ (.A(_07306_),
    .X(_07913_));
 sky130_fd_sc_hd__nand3b_2 _29540_ (.A_N(_07908_),
    .B(_06227_),
    .C(_07913_),
    .Y(_07914_));
 sky130_fd_sc_hd__nand3b_2 _29541_ (.A_N(_07907_),
    .B(_07914_),
    .C(_07911_),
    .Y(_07915_));
 sky130_fd_sc_hd__nand2_2 _29542_ (.A(_07912_),
    .B(_07915_),
    .Y(_07916_));
 sky130_fd_sc_hd__a21oi_2 _29543_ (.A1(_07815_),
    .A2(_07820_),
    .B1(_07816_),
    .Y(_07917_));
 sky130_fd_sc_hd__nand2_2 _29544_ (.A(_07916_),
    .B(_07917_),
    .Y(_07918_));
 sky130_fd_sc_hd__nand3b_2 _29545_ (.A_N(_07917_),
    .B(_07915_),
    .C(_07912_),
    .Y(_07919_));
 sky130_fd_sc_hd__buf_1 _29546_ (.A(_06113_),
    .X(_07920_));
 sky130_fd_sc_hd__o31a_2 _29547_ (.A1(_07920_),
    .A2(_19227_),
    .A3(_07689_),
    .B1(_07700_),
    .X(_07921_));
 sky130_vsdinv _29548_ (.A(_07921_),
    .Y(_07922_));
 sky130_fd_sc_hd__a21oi_2 _29549_ (.A1(_07918_),
    .A2(_07919_),
    .B1(_07922_),
    .Y(_07923_));
 sky130_fd_sc_hd__nand3_2 _29550_ (.A(_07918_),
    .B(_07922_),
    .C(_07919_),
    .Y(_07924_));
 sky130_vsdinv _29551_ (.A(_07924_),
    .Y(_07925_));
 sky130_fd_sc_hd__a21boi_2 _29552_ (.A1(_07829_),
    .A2(_07831_),
    .B1_N(_07832_),
    .Y(_07926_));
 sky130_fd_sc_hd__o21ai_2 _29553_ (.A1(_07822_),
    .A2(_07926_),
    .B1(_07834_),
    .Y(_07927_));
 sky130_fd_sc_hd__o21bai_2 _29554_ (.A1(_07923_),
    .A2(_07925_),
    .B1_N(_07927_),
    .Y(_07928_));
 sky130_fd_sc_hd__a21o_2 _29555_ (.A1(_07918_),
    .A2(_07919_),
    .B1(_07922_),
    .X(_07929_));
 sky130_fd_sc_hd__nand3_2 _29556_ (.A(_07929_),
    .B(_07927_),
    .C(_07924_),
    .Y(_07930_));
 sky130_fd_sc_hd__buf_1 _29557_ (.A(_07930_),
    .X(_07931_));
 sky130_fd_sc_hd__a21boi_2 _29558_ (.A1(_07704_),
    .A2(_07708_),
    .B1_N(_07706_),
    .Y(_07932_));
 sky130_vsdinv _29559_ (.A(_07932_),
    .Y(_07933_));
 sky130_fd_sc_hd__a21oi_2 _29560_ (.A1(_07928_),
    .A2(_07931_),
    .B1(_07933_),
    .Y(_07934_));
 sky130_vsdinv _29561_ (.A(_07706_),
    .Y(_07935_));
 sky130_fd_sc_hd__o211a_2 _29562_ (.A1(_07935_),
    .A2(_07711_),
    .B1(_07930_),
    .C1(_07928_),
    .X(_07936_));
 sky130_fd_sc_hd__o21ai_2 _29563_ (.A1(_07718_),
    .A2(_07726_),
    .B1(_07717_),
    .Y(_07937_));
 sky130_fd_sc_hd__o21bai_2 _29564_ (.A1(_07934_),
    .A2(_07936_),
    .B1_N(_07937_),
    .Y(_07938_));
 sky130_fd_sc_hd__a21o_2 _29565_ (.A1(_07928_),
    .A2(_07931_),
    .B1(_07933_),
    .X(_07939_));
 sky130_fd_sc_hd__nand3_2 _29566_ (.A(_07928_),
    .B(_07933_),
    .C(_07931_),
    .Y(_07940_));
 sky130_fd_sc_hd__nand3_2 _29567_ (.A(_07939_),
    .B(_07940_),
    .C(_07937_),
    .Y(_07941_));
 sky130_fd_sc_hd__buf_1 _29568_ (.A(_07748_),
    .X(_07942_));
 sky130_fd_sc_hd__a22o_2 _29569_ (.A1(_07595_),
    .A2(_07606_),
    .B1(_05504_),
    .B2(_07942_),
    .X(_07943_));
 sky130_fd_sc_hd__buf_1 _29570_ (.A(_19207_),
    .X(_07944_));
 sky130_fd_sc_hd__nand2_2 _29571_ (.A(_05939_),
    .B(_07944_),
    .Y(_07945_));
 sky130_fd_sc_hd__buf_1 _29572_ (.A(\pcpi_mul.rs1[17] ),
    .X(_07946_));
 sky130_fd_sc_hd__buf_1 _29573_ (.A(_07946_),
    .X(_07947_));
 sky130_fd_sc_hd__buf_1 _29574_ (.A(_07947_),
    .X(_07948_));
 sky130_fd_sc_hd__nand3b_2 _29575_ (.A_N(_07945_),
    .B(_05825_),
    .C(_07948_),
    .Y(_07949_));
 sky130_fd_sc_hd__o2bb2ai_2 _29576_ (.A1_N(_07943_),
    .A2_N(_07949_),
    .B1(_06347_),
    .B2(_19188_),
    .Y(_07950_));
 sky130_fd_sc_hd__buf_1 _29577_ (.A(_19184_),
    .X(_07951_));
 sky130_fd_sc_hd__buf_1 _29578_ (.A(_07951_),
    .X(_07952_));
 sky130_fd_sc_hd__and2_2 _29579_ (.A(_05236_),
    .B(_07952_),
    .X(_07953_));
 sky130_fd_sc_hd__nand3_2 _29580_ (.A(_07949_),
    .B(_07943_),
    .C(_07953_),
    .Y(_07954_));
 sky130_fd_sc_hd__a21oi_2 _29581_ (.A1(_07735_),
    .A2(_07734_),
    .B1(_07732_),
    .Y(_07955_));
 sky130_vsdinv _29582_ (.A(_07955_),
    .Y(_07956_));
 sky130_fd_sc_hd__a21o_2 _29583_ (.A1(_07950_),
    .A2(_07954_),
    .B1(_07956_),
    .X(_07957_));
 sky130_fd_sc_hd__nand3_2 _29584_ (.A(_07950_),
    .B(_07956_),
    .C(_07954_),
    .Y(_07958_));
 sky130_fd_sc_hd__buf_1 _29585_ (.A(_07958_),
    .X(_07959_));
 sky130_fd_sc_hd__buf_1 _29586_ (.A(\pcpi_mul.rs1[20] ),
    .X(_07960_));
 sky130_fd_sc_hd__buf_1 _29587_ (.A(_07960_),
    .X(_07961_));
 sky130_fd_sc_hd__nand2_2 _29588_ (.A(_18866_),
    .B(_07961_),
    .Y(_07962_));
 sky130_fd_sc_hd__buf_1 _29589_ (.A(_19190_),
    .X(_07963_));
 sky130_fd_sc_hd__nand2_2 _29590_ (.A(_05663_),
    .B(_07963_),
    .Y(_07964_));
 sky130_fd_sc_hd__xor2_2 _29591_ (.A(_07962_),
    .B(_07964_),
    .X(_07965_));
 sky130_fd_sc_hd__buf_1 _29592_ (.A(_07309_),
    .X(_07966_));
 sky130_fd_sc_hd__buf_1 _29593_ (.A(_07966_),
    .X(_07967_));
 sky130_fd_sc_hd__and2_2 _29594_ (.A(_07121_),
    .B(_07967_),
    .X(_07968_));
 sky130_fd_sc_hd__nand2_2 _29595_ (.A(_07965_),
    .B(_07968_),
    .Y(_07969_));
 sky130_fd_sc_hd__xnor2_2 _29596_ (.A(_07962_),
    .B(_07964_),
    .Y(_07970_));
 sky130_fd_sc_hd__o21ai_2 _29597_ (.A1(_18857_),
    .A2(_19205_),
    .B1(_07970_),
    .Y(_07971_));
 sky130_fd_sc_hd__nand2_2 _29598_ (.A(_07969_),
    .B(_07971_),
    .Y(_07972_));
 sky130_fd_sc_hd__buf_1 _29599_ (.A(_07972_),
    .X(_07973_));
 sky130_fd_sc_hd__a21boi_2 _29600_ (.A1(_07957_),
    .A2(_07959_),
    .B1_N(_07973_),
    .Y(_07974_));
 sky130_fd_sc_hd__a21oi_2 _29601_ (.A1(_07950_),
    .A2(_07954_),
    .B1(_07956_),
    .Y(_07975_));
 sky130_fd_sc_hd__nor3b_2 _29602_ (.A(_07973_),
    .B(_07975_),
    .C_N(_07958_),
    .Y(_07976_));
 sky130_fd_sc_hd__a21boi_2 _29603_ (.A1(_07736_),
    .A2(_07739_),
    .B1_N(_07740_),
    .Y(_07977_));
 sky130_fd_sc_hd__o21ai_2 _29604_ (.A1(_07756_),
    .A2(_07977_),
    .B1(_07742_),
    .Y(_07978_));
 sky130_fd_sc_hd__o21bai_2 _29605_ (.A1(_07974_),
    .A2(_07976_),
    .B1_N(_07978_),
    .Y(_07979_));
 sky130_vsdinv _29606_ (.A(_07972_),
    .Y(_07980_));
 sky130_fd_sc_hd__a21o_2 _29607_ (.A1(_07957_),
    .A2(_07959_),
    .B1(_07980_),
    .X(_07981_));
 sky130_fd_sc_hd__nand3b_2 _29608_ (.A_N(_07973_),
    .B(_07957_),
    .C(_07959_),
    .Y(_07982_));
 sky130_fd_sc_hd__nand3_2 _29609_ (.A(_07981_),
    .B(_07978_),
    .C(_07982_),
    .Y(_07983_));
 sky130_fd_sc_hd__a21oi_2 _29610_ (.A1(_07747_),
    .A2(_07749_),
    .B1(_07754_),
    .Y(_07984_));
 sky130_vsdinv _29611_ (.A(_07984_),
    .Y(_07985_));
 sky130_fd_sc_hd__a21oi_2 _29612_ (.A1(_07979_),
    .A2(_07983_),
    .B1(_07985_),
    .Y(_07986_));
 sky130_fd_sc_hd__nand3_2 _29613_ (.A(_07979_),
    .B(_07985_),
    .C(_07983_),
    .Y(_07987_));
 sky130_vsdinv _29614_ (.A(_07987_),
    .Y(_07988_));
 sky130_fd_sc_hd__nor2_2 _29615_ (.A(_07986_),
    .B(_07988_),
    .Y(_07989_));
 sky130_fd_sc_hd__a21oi_2 _29616_ (.A1(_07938_),
    .A2(_07941_),
    .B1(_07989_),
    .Y(_07990_));
 sky130_fd_sc_hd__or2b_2 _29617_ (.A(_07986_),
    .B_N(_07987_),
    .X(_07991_));
 sky130_fd_sc_hd__nand2_2 _29618_ (.A(_07938_),
    .B(_07941_),
    .Y(_07992_));
 sky130_fd_sc_hd__nor2_2 _29619_ (.A(_07991_),
    .B(_07992_),
    .Y(_07993_));
 sky130_fd_sc_hd__o21bai_2 _29620_ (.A1(_07990_),
    .A2(_07993_),
    .B1_N(_07843_),
    .Y(_07994_));
 sky130_fd_sc_hd__o21ai_2 _29621_ (.A1(_07770_),
    .A2(_07771_),
    .B1(_07729_),
    .Y(_07995_));
 sky130_fd_sc_hd__nand2_2 _29622_ (.A(_07992_),
    .B(_07991_),
    .Y(_07996_));
 sky130_fd_sc_hd__nand3_2 _29623_ (.A(_07989_),
    .B(_07938_),
    .C(_07941_),
    .Y(_07997_));
 sky130_fd_sc_hd__nand3_2 _29624_ (.A(_07996_),
    .B(_07843_),
    .C(_07997_),
    .Y(_07998_));
 sky130_fd_sc_hd__nand3_2 _29625_ (.A(_07994_),
    .B(_07995_),
    .C(_07998_),
    .Y(_07999_));
 sky130_fd_sc_hd__a21oi_2 _29626_ (.A1(_07996_),
    .A2(_07997_),
    .B1(_07843_),
    .Y(_08000_));
 sky130_fd_sc_hd__nor3_2 _29627_ (.A(_07842_),
    .B(_07990_),
    .C(_07993_),
    .Y(_08001_));
 sky130_fd_sc_hd__o21bai_2 _29628_ (.A1(_08000_),
    .A2(_08001_),
    .B1_N(_07995_),
    .Y(_08002_));
 sky130_fd_sc_hd__buf_1 _29629_ (.A(_05527_),
    .X(_08003_));
 sky130_fd_sc_hd__nand2_2 _29630_ (.A(_07006_),
    .B(_08003_),
    .Y(_08004_));
 sky130_fd_sc_hd__nand2_2 _29631_ (.A(_18785_),
    .B(_05851_),
    .Y(_08005_));
 sky130_fd_sc_hd__nor2_2 _29632_ (.A(_08004_),
    .B(_08005_),
    .Y(_08006_));
 sky130_fd_sc_hd__buf_1 _29633_ (.A(_19267_),
    .X(_08007_));
 sky130_fd_sc_hd__and2_2 _29634_ (.A(_07477_),
    .B(_08007_),
    .X(_08008_));
 sky130_fd_sc_hd__nand2_2 _29635_ (.A(_08004_),
    .B(_08005_),
    .Y(_08009_));
 sky130_fd_sc_hd__nand3b_2 _29636_ (.A_N(_08006_),
    .B(_08008_),
    .C(_08009_),
    .Y(_08010_));
 sky130_fd_sc_hd__buf_1 _29637_ (.A(_07165_),
    .X(_08011_));
 sky130_fd_sc_hd__buf_1 _29638_ (.A(_07167_),
    .X(_08012_));
 sky130_fd_sc_hd__buf_1 _29639_ (.A(_08012_),
    .X(_08013_));
 sky130_fd_sc_hd__a22oi_2 _29640_ (.A1(_08011_),
    .A2(_06102_),
    .B1(_08013_),
    .B2(_06052_),
    .Y(_08014_));
 sky130_fd_sc_hd__o21bai_2 _29641_ (.A1(_08014_),
    .A2(_08006_),
    .B1_N(_08008_),
    .Y(_08015_));
 sky130_fd_sc_hd__nand2_2 _29642_ (.A(_08010_),
    .B(_08015_),
    .Y(_08016_));
 sky130_fd_sc_hd__nand2_2 _29643_ (.A(_07852_),
    .B(_07854_),
    .Y(_08017_));
 sky130_fd_sc_hd__nor2_2 _29644_ (.A(_07852_),
    .B(_07854_),
    .Y(_08018_));
 sky130_fd_sc_hd__a21oi_2 _29645_ (.A1(_08017_),
    .A2(_07849_),
    .B1(_08018_),
    .Y(_08019_));
 sky130_fd_sc_hd__nand2_2 _29646_ (.A(_08016_),
    .B(_08019_),
    .Y(_08020_));
 sky130_fd_sc_hd__nand3b_2 _29647_ (.A_N(_08019_),
    .B(_08010_),
    .C(_08015_),
    .Y(_08021_));
 sky130_fd_sc_hd__o31a_2 _29648_ (.A1(_07178_),
    .A2(_19274_),
    .A3(_07789_),
    .B1(_07796_),
    .X(_08022_));
 sky130_vsdinv _29649_ (.A(_08022_),
    .Y(_08023_));
 sky130_fd_sc_hd__a21oi_2 _29650_ (.A1(_08020_),
    .A2(_08021_),
    .B1(_08023_),
    .Y(_08024_));
 sky130_fd_sc_hd__nand3_2 _29651_ (.A(_08020_),
    .B(_08023_),
    .C(_08021_),
    .Y(_08025_));
 sky130_vsdinv _29652_ (.A(_08025_),
    .Y(_08026_));
 sky130_fd_sc_hd__nand2_2 _29653_ (.A(_07808_),
    .B(_07803_),
    .Y(_08027_));
 sky130_fd_sc_hd__o21bai_2 _29654_ (.A1(_08024_),
    .A2(_08026_),
    .B1_N(_08027_),
    .Y(_08028_));
 sky130_fd_sc_hd__a21o_2 _29655_ (.A1(_08020_),
    .A2(_08021_),
    .B1(_08023_),
    .X(_08029_));
 sky130_fd_sc_hd__nand3_2 _29656_ (.A(_08027_),
    .B(_08029_),
    .C(_08025_),
    .Y(_08030_));
 sky130_fd_sc_hd__buf_1 _29657_ (.A(_08030_),
    .X(_08031_));
 sky130_fd_sc_hd__buf_1 _29658_ (.A(_06533_),
    .X(_08032_));
 sky130_fd_sc_hd__nand2_2 _29659_ (.A(_08032_),
    .B(_05841_),
    .Y(_08033_));
 sky130_fd_sc_hd__buf_1 _29660_ (.A(_18801_),
    .X(_08034_));
 sky130_fd_sc_hd__buf_1 _29661_ (.A(_19257_),
    .X(_08035_));
 sky130_fd_sc_hd__nand2_2 _29662_ (.A(_08034_),
    .B(_08035_),
    .Y(_08036_));
 sky130_fd_sc_hd__nor2_2 _29663_ (.A(_08033_),
    .B(_08036_),
    .Y(_08037_));
 sky130_fd_sc_hd__buf_1 _29664_ (.A(\pcpi_mul.rs2[12] ),
    .X(_08038_));
 sky130_fd_sc_hd__buf_1 _29665_ (.A(_08038_),
    .X(_08039_));
 sky130_fd_sc_hd__and2_2 _29666_ (.A(_08039_),
    .B(_06199_),
    .X(_08040_));
 sky130_fd_sc_hd__nand2_2 _29667_ (.A(_08033_),
    .B(_08036_),
    .Y(_08041_));
 sky130_fd_sc_hd__nand3b_2 _29668_ (.A_N(_08037_),
    .B(_08040_),
    .C(_08041_),
    .Y(_08042_));
 sky130_fd_sc_hd__buf_1 _29669_ (.A(_06537_),
    .X(_08043_));
 sky130_fd_sc_hd__a22oi_2 _29670_ (.A1(_06535_),
    .A2(_05842_),
    .B1(_08043_),
    .B2(_05951_),
    .Y(_08044_));
 sky130_fd_sc_hd__o21bai_2 _29671_ (.A1(_08044_),
    .A2(_08037_),
    .B1_N(_08040_),
    .Y(_08045_));
 sky130_fd_sc_hd__a21oi_2 _29672_ (.A1(_07828_),
    .A2(_07827_),
    .B1(_07826_),
    .Y(_08046_));
 sky130_fd_sc_hd__a21boi_2 _29673_ (.A1(_08042_),
    .A2(_08045_),
    .B1_N(_08046_),
    .Y(_08047_));
 sky130_fd_sc_hd__nand2_2 _29674_ (.A(_18814_),
    .B(_06360_),
    .Y(_08048_));
 sky130_fd_sc_hd__nand2_2 _29675_ (.A(_18819_),
    .B(_06365_),
    .Y(_08049_));
 sky130_fd_sc_hd__nand2_2 _29676_ (.A(_08048_),
    .B(_08049_),
    .Y(_08050_));
 sky130_fd_sc_hd__nor2_2 _29677_ (.A(_08048_),
    .B(_08049_),
    .Y(_08051_));
 sky130_vsdinv _29678_ (.A(_08051_),
    .Y(_08052_));
 sky130_fd_sc_hd__o2bb2ai_2 _29679_ (.A1_N(_08050_),
    .A2_N(_08052_),
    .B1(_07818_),
    .B2(_19239_),
    .Y(_08053_));
 sky130_fd_sc_hd__buf_1 _29680_ (.A(_07551_),
    .X(_08054_));
 sky130_fd_sc_hd__and2_2 _29681_ (.A(_05895_),
    .B(_08054_),
    .X(_08055_));
 sky130_fd_sc_hd__nand3b_2 _29682_ (.A_N(_08051_),
    .B(_08055_),
    .C(_08050_),
    .Y(_08056_));
 sky130_fd_sc_hd__nand2_2 _29683_ (.A(_08053_),
    .B(_08056_),
    .Y(_08057_));
 sky130_vsdinv _29684_ (.A(_08057_),
    .Y(_08058_));
 sky130_fd_sc_hd__nand3b_2 _29685_ (.A_N(_08046_),
    .B(_08042_),
    .C(_08045_),
    .Y(_08059_));
 sky130_fd_sc_hd__nand3b_2 _29686_ (.A_N(_08047_),
    .B(_08058_),
    .C(_08059_),
    .Y(_08060_));
 sky130_vsdinv _29687_ (.A(_08059_),
    .Y(_08061_));
 sky130_fd_sc_hd__o21ai_2 _29688_ (.A1(_08047_),
    .A2(_08061_),
    .B1(_08057_),
    .Y(_08062_));
 sky130_fd_sc_hd__nand2_2 _29689_ (.A(_08060_),
    .B(_08062_),
    .Y(_08063_));
 sky130_vsdinv _29690_ (.A(_08063_),
    .Y(_08064_));
 sky130_fd_sc_hd__a21oi_2 _29691_ (.A1(_08028_),
    .A2(_08031_),
    .B1(_08064_),
    .Y(_08065_));
 sky130_fd_sc_hd__a21oi_2 _29692_ (.A1(_08029_),
    .A2(_08025_),
    .B1(_08027_),
    .Y(_08066_));
 sky130_fd_sc_hd__nor3b_2 _29693_ (.A(_08063_),
    .B(_08066_),
    .C_N(_08031_),
    .Y(_08067_));
 sky130_fd_sc_hd__o21ai_2 _29694_ (.A1(_07810_),
    .A2(_07836_),
    .B1(_07811_),
    .Y(_08068_));
 sky130_fd_sc_hd__o21bai_2 _29695_ (.A1(_08065_),
    .A2(_08067_),
    .B1_N(_08068_),
    .Y(_08069_));
 sky130_fd_sc_hd__a21o_2 _29696_ (.A1(_08028_),
    .A2(_08031_),
    .B1(_08064_),
    .X(_08070_));
 sky130_fd_sc_hd__nand3_2 _29697_ (.A(_08028_),
    .B(_08064_),
    .C(_08031_),
    .Y(_08071_));
 sky130_fd_sc_hd__nand3_2 _29698_ (.A(_08070_),
    .B(_08068_),
    .C(_08071_),
    .Y(_08072_));
 sky130_fd_sc_hd__buf_1 _29699_ (.A(_08072_),
    .X(_08073_));
 sky130_fd_sc_hd__buf_1 _29700_ (.A(_07850_),
    .X(_08074_));
 sky130_fd_sc_hd__nand2_2 _29701_ (.A(_08074_),
    .B(_05412_),
    .Y(_08075_));
 sky130_fd_sc_hd__nand2_2 _29702_ (.A(_07535_),
    .B(_05551_),
    .Y(_08076_));
 sky130_fd_sc_hd__nand2_2 _29703_ (.A(_08075_),
    .B(_08076_),
    .Y(_08077_));
 sky130_fd_sc_hd__nor2_2 _29704_ (.A(_08075_),
    .B(_08076_),
    .Y(_08078_));
 sky130_vsdinv _29705_ (.A(_08078_),
    .Y(_08079_));
 sky130_fd_sc_hd__o2bb2ai_2 _29706_ (.A1_N(_08077_),
    .A2_N(_08079_),
    .B1(_18777_),
    .B2(_19283_),
    .Y(_08080_));
 sky130_fd_sc_hd__and2_2 _29707_ (.A(_07533_),
    .B(_07790_),
    .X(_08081_));
 sky130_fd_sc_hd__nand3b_2 _29708_ (.A_N(_08078_),
    .B(_08081_),
    .C(_08077_),
    .Y(_08082_));
 sky130_fd_sc_hd__nand2_2 _29709_ (.A(_18755_),
    .B(_05240_),
    .Y(_08083_));
 sky130_fd_sc_hd__buf_1 _29710_ (.A(_18758_),
    .X(_08084_));
 sky130_fd_sc_hd__buf_1 _29711_ (.A(_08084_),
    .X(_08085_));
 sky130_fd_sc_hd__buf_1 _29712_ (.A(_08085_),
    .X(_08086_));
 sky130_fd_sc_hd__nand2_2 _29713_ (.A(_08086_),
    .B(_05403_),
    .Y(_08087_));
 sky130_fd_sc_hd__xor2_2 _29714_ (.A(_08083_),
    .B(_08087_),
    .X(_08088_));
 sky130_fd_sc_hd__a21o_2 _29715_ (.A1(_08080_),
    .A2(_08082_),
    .B1(_08088_),
    .X(_08089_));
 sky130_fd_sc_hd__nand3_2 _29716_ (.A(_08080_),
    .B(_08088_),
    .C(_08082_),
    .Y(_08090_));
 sky130_fd_sc_hd__nand2_2 _29717_ (.A(_08089_),
    .B(_08090_),
    .Y(_08091_));
 sky130_fd_sc_hd__o31a_2 _29718_ (.A1(_18761_),
    .A2(_19302_),
    .A3(_07856_),
    .B1(_08091_),
    .X(_08092_));
 sky130_fd_sc_hd__nand3b_2 _29719_ (.A_N(_07856_),
    .B(_07847_),
    .C(_05242_),
    .Y(_08093_));
 sky130_fd_sc_hd__nor2_2 _29720_ (.A(_08091_),
    .B(_08093_),
    .Y(_08094_));
 sky130_fd_sc_hd__buf_1 _29721_ (.A(_08094_),
    .X(_08095_));
 sky130_fd_sc_hd__nor2_2 _29722_ (.A(_08092_),
    .B(_08095_),
    .Y(_08096_));
 sky130_fd_sc_hd__a21oi_2 _29723_ (.A1(_08069_),
    .A2(_08073_),
    .B1(_08096_),
    .Y(_08097_));
 sky130_fd_sc_hd__nand3_2 _29724_ (.A(_08069_),
    .B(_08096_),
    .C(_08072_),
    .Y(_08098_));
 sky130_vsdinv _29725_ (.A(_08098_),
    .Y(_08099_));
 sky130_fd_sc_hd__nor3_2 _29726_ (.A(_07860_),
    .B(_08097_),
    .C(_08099_),
    .Y(_08100_));
 sky130_fd_sc_hd__o2bb2ai_2 _29727_ (.A1_N(_08073_),
    .A2_N(_08069_),
    .B1(_08092_),
    .B2(_08095_),
    .Y(_08101_));
 sky130_fd_sc_hd__a21boi_2 _29728_ (.A1(_08101_),
    .A2(_08098_),
    .B1_N(_07860_),
    .Y(_08102_));
 sky130_fd_sc_hd__o2bb2ai_2 _29729_ (.A1_N(_07999_),
    .A2_N(_08002_),
    .B1(_08100_),
    .B2(_08102_),
    .Y(_08103_));
 sky130_fd_sc_hd__nor2_2 _29730_ (.A(_08102_),
    .B(_08100_),
    .Y(_08104_));
 sky130_fd_sc_hd__nand3_2 _29731_ (.A(_08002_),
    .B(_08104_),
    .C(_07999_),
    .Y(_08105_));
 sky130_fd_sc_hd__nand2_2 _29732_ (.A(_08103_),
    .B(_08105_),
    .Y(_08106_));
 sky130_fd_sc_hd__a31oi_2 _29733_ (.A1(_07868_),
    .A2(_07865_),
    .A3(_07869_),
    .B1(_07864_),
    .Y(_08107_));
 sky130_fd_sc_hd__nand2_2 _29734_ (.A(_08106_),
    .B(_08107_),
    .Y(_08108_));
 sky130_fd_sc_hd__o31ai_2 _29735_ (.A1(_07543_),
    .A2(_07863_),
    .A3(_07862_),
    .B1(_07870_),
    .Y(_08109_));
 sky130_fd_sc_hd__nand3_2 _29736_ (.A(_08109_),
    .B(_08105_),
    .C(_08103_),
    .Y(_08110_));
 sky130_fd_sc_hd__o21a_2 _29737_ (.A1(_07765_),
    .A2(_07764_),
    .B1(_07763_),
    .X(_08111_));
 sky130_fd_sc_hd__a21boi_2 _29738_ (.A1(_07776_),
    .A2(_07782_),
    .B1_N(_07780_),
    .Y(_08112_));
 sky130_fd_sc_hd__xor2_2 _29739_ (.A(_08111_),
    .B(_08112_),
    .X(_08113_));
 sky130_fd_sc_hd__a21oi_2 _29740_ (.A1(_08108_),
    .A2(_08110_),
    .B1(_08113_),
    .Y(_08114_));
 sky130_fd_sc_hd__nand3_2 _29741_ (.A(_08108_),
    .B(_08110_),
    .C(_08113_),
    .Y(_08115_));
 sky130_vsdinv _29742_ (.A(_08115_),
    .Y(_08116_));
 sky130_fd_sc_hd__o21ai_2 _29743_ (.A1(_07882_),
    .A2(_07883_),
    .B1(_07877_),
    .Y(_08117_));
 sky130_fd_sc_hd__o21bai_2 _29744_ (.A1(_08114_),
    .A2(_08116_),
    .B1_N(_08117_),
    .Y(_08118_));
 sky130_fd_sc_hd__a21o_2 _29745_ (.A1(_08108_),
    .A2(_08110_),
    .B1(_08113_),
    .X(_08119_));
 sky130_fd_sc_hd__nand3_2 _29746_ (.A(_08119_),
    .B(_08115_),
    .C(_08117_),
    .Y(_08120_));
 sky130_fd_sc_hd__buf_1 _29747_ (.A(_08120_),
    .X(_08121_));
 sky130_fd_sc_hd__a21oi_2 _29748_ (.A1(_07646_),
    .A2(_07636_),
    .B1(_07878_),
    .Y(_08122_));
 sky130_fd_sc_hd__a21o_2 _29749_ (.A1(_08118_),
    .A2(_08121_),
    .B1(_08122_),
    .X(_08123_));
 sky130_fd_sc_hd__nand3_2 _29750_ (.A(_08118_),
    .B(_08122_),
    .C(_08120_),
    .Y(_08124_));
 sky130_fd_sc_hd__o21ai_2 _29751_ (.A1(_07895_),
    .A2(_07896_),
    .B1(_07891_),
    .Y(_08125_));
 sky130_fd_sc_hd__a21oi_2 _29752_ (.A1(_08123_),
    .A2(_08124_),
    .B1(_08125_),
    .Y(_08126_));
 sky130_fd_sc_hd__a21boi_2 _29753_ (.A1(_07886_),
    .A2(_07893_),
    .B1_N(_07891_),
    .Y(_08127_));
 sky130_fd_sc_hd__a21oi_2 _29754_ (.A1(_08118_),
    .A2(_08121_),
    .B1(_08122_),
    .Y(_08128_));
 sky130_fd_sc_hd__nor3b_2 _29755_ (.A(_08127_),
    .B(_08128_),
    .C_N(_08124_),
    .Y(_08129_));
 sky130_fd_sc_hd__nor2_2 _29756_ (.A(_08126_),
    .B(_08129_),
    .Y(_08130_));
 sky130_fd_sc_hd__nor2_2 _29757_ (.A(_07680_),
    .B(_07904_),
    .Y(_08131_));
 sky130_fd_sc_hd__a21oi_2 _29758_ (.A1(_07901_),
    .A2(_07902_),
    .B1(_07899_),
    .Y(_08132_));
 sky130_fd_sc_hd__a21oi_2 _29759_ (.A1(_07679_),
    .A2(_07903_),
    .B1(_08132_),
    .Y(_08133_));
 sky130_fd_sc_hd__a21oi_2 _29760_ (.A1(_07687_),
    .A2(_08131_),
    .B1(_08133_),
    .Y(_08134_));
 sky130_fd_sc_hd__xnor2_2 _29761_ (.A(_08130_),
    .B(_08134_),
    .Y(_02641_));
 sky130_fd_sc_hd__nand2_2 _29762_ (.A(_08115_),
    .B(_08110_),
    .Y(_08135_));
 sky130_fd_sc_hd__a22oi_2 _29763_ (.A1(_07392_),
    .A2(_05666_),
    .B1(_08013_),
    .B2(_05838_),
    .Y(_08136_));
 sky130_fd_sc_hd__nand2_2 _29764_ (.A(_07472_),
    .B(_07365_),
    .Y(_08137_));
 sky130_fd_sc_hd__nand2_2 _29765_ (.A(_07788_),
    .B(_06180_),
    .Y(_08138_));
 sky130_fd_sc_hd__nor2_2 _29766_ (.A(_08137_),
    .B(_08138_),
    .Y(_08139_));
 sky130_fd_sc_hd__and2_2 _29767_ (.A(_07477_),
    .B(_05728_),
    .X(_08140_));
 sky130_fd_sc_hd__o21bai_2 _29768_ (.A1(_08136_),
    .A2(_08139_),
    .B1_N(_08140_),
    .Y(_08141_));
 sky130_fd_sc_hd__buf_1 _29769_ (.A(_07004_),
    .X(_08142_));
 sky130_fd_sc_hd__nand3b_2 _29770_ (.A_N(_08137_),
    .B(_08142_),
    .C(_05964_),
    .Y(_08143_));
 sky130_fd_sc_hd__nand2_2 _29771_ (.A(_08137_),
    .B(_08138_),
    .Y(_08144_));
 sky130_fd_sc_hd__nand3_2 _29772_ (.A(_08143_),
    .B(_08140_),
    .C(_08144_),
    .Y(_08145_));
 sky130_fd_sc_hd__nand2_2 _29773_ (.A(_08141_),
    .B(_08145_),
    .Y(_08146_));
 sky130_fd_sc_hd__a21o_2 _29774_ (.A1(_08077_),
    .A2(_08081_),
    .B1(_08078_),
    .X(_08147_));
 sky130_vsdinv _29775_ (.A(_08147_),
    .Y(_08148_));
 sky130_fd_sc_hd__nand2_2 _29776_ (.A(_08146_),
    .B(_08148_),
    .Y(_08149_));
 sky130_fd_sc_hd__nand3_2 _29777_ (.A(_08141_),
    .B(_08147_),
    .C(_08145_),
    .Y(_08150_));
 sky130_fd_sc_hd__a21oi_2 _29778_ (.A1(_08009_),
    .A2(_08008_),
    .B1(_08006_),
    .Y(_08151_));
 sky130_vsdinv _29779_ (.A(_08151_),
    .Y(_08152_));
 sky130_fd_sc_hd__a21oi_2 _29780_ (.A1(_08149_),
    .A2(_08150_),
    .B1(_08152_),
    .Y(_08153_));
 sky130_fd_sc_hd__nand3_2 _29781_ (.A(_08149_),
    .B(_08152_),
    .C(_08150_),
    .Y(_08154_));
 sky130_vsdinv _29782_ (.A(_08154_),
    .Y(_08155_));
 sky130_fd_sc_hd__a21boi_2 _29783_ (.A1(_08010_),
    .A2(_08015_),
    .B1_N(_08019_),
    .Y(_08156_));
 sky130_fd_sc_hd__o21ai_2 _29784_ (.A1(_08022_),
    .A2(_08156_),
    .B1(_08021_),
    .Y(_08157_));
 sky130_fd_sc_hd__o21bai_2 _29785_ (.A1(_08153_),
    .A2(_08155_),
    .B1_N(_08157_),
    .Y(_08158_));
 sky130_fd_sc_hd__nand2_2 _29786_ (.A(_08149_),
    .B(_08150_),
    .Y(_08159_));
 sky130_fd_sc_hd__nand2_2 _29787_ (.A(_08159_),
    .B(_08151_),
    .Y(_08160_));
 sky130_fd_sc_hd__nand3_2 _29788_ (.A(_08160_),
    .B(_08157_),
    .C(_08154_),
    .Y(_08161_));
 sky130_fd_sc_hd__nand2_2 _29789_ (.A(_08158_),
    .B(_08161_),
    .Y(_08162_));
 sky130_fd_sc_hd__nand2_2 _29790_ (.A(_06534_),
    .B(_08035_),
    .Y(_08163_));
 sky130_fd_sc_hd__nand2_2 _29791_ (.A(_08034_),
    .B(_05935_),
    .Y(_08164_));
 sky130_fd_sc_hd__nor2_2 _29792_ (.A(_08163_),
    .B(_08164_),
    .Y(_08165_));
 sky130_fd_sc_hd__and2_2 _29793_ (.A(_08039_),
    .B(_06360_),
    .X(_08166_));
 sky130_fd_sc_hd__nand2_2 _29794_ (.A(_08163_),
    .B(_08164_),
    .Y(_08167_));
 sky130_fd_sc_hd__nand3b_2 _29795_ (.A_N(_08165_),
    .B(_08166_),
    .C(_08167_),
    .Y(_08168_));
 sky130_fd_sc_hd__buf_1 _29796_ (.A(_06543_),
    .X(_08169_));
 sky130_fd_sc_hd__buf_1 _29797_ (.A(_08169_),
    .X(_08170_));
 sky130_fd_sc_hd__a22oi_2 _29798_ (.A1(_08170_),
    .A2(_05959_),
    .B1(_18803_),
    .B2(_06358_),
    .Y(_08171_));
 sky130_fd_sc_hd__o21bai_2 _29799_ (.A1(_08171_),
    .A2(_08165_),
    .B1_N(_08166_),
    .Y(_08172_));
 sky130_fd_sc_hd__nand2_2 _29800_ (.A(_08168_),
    .B(_08172_),
    .Y(_08173_));
 sky130_fd_sc_hd__a21oi_2 _29801_ (.A1(_08041_),
    .A2(_08040_),
    .B1(_08037_),
    .Y(_08174_));
 sky130_fd_sc_hd__nand2_2 _29802_ (.A(_08173_),
    .B(_08174_),
    .Y(_08175_));
 sky130_fd_sc_hd__nand3b_2 _29803_ (.A_N(_08174_),
    .B(_08168_),
    .C(_08172_),
    .Y(_08176_));
 sky130_fd_sc_hd__nand2_2 _29804_ (.A(_08175_),
    .B(_08176_),
    .Y(_08177_));
 sky130_fd_sc_hd__buf_1 _29805_ (.A(_18813_),
    .X(_08178_));
 sky130_fd_sc_hd__nand2_2 _29806_ (.A(_08178_),
    .B(_06728_),
    .Y(_08179_));
 sky130_fd_sc_hd__buf_1 _29807_ (.A(_06140_),
    .X(_08180_));
 sky130_fd_sc_hd__buf_1 _29808_ (.A(_07098_),
    .X(_08181_));
 sky130_fd_sc_hd__nand2_2 _29809_ (.A(_08180_),
    .B(_08181_),
    .Y(_08182_));
 sky130_fd_sc_hd__xnor2_2 _29810_ (.A(_08179_),
    .B(_08182_),
    .Y(_08183_));
 sky130_fd_sc_hd__o21ai_2 _29811_ (.A1(_07818_),
    .A2(_19234_),
    .B1(_08183_),
    .Y(_08184_));
 sky130_fd_sc_hd__nor2_2 _29812_ (.A(_08179_),
    .B(_08182_),
    .Y(_08185_));
 sky130_fd_sc_hd__buf_1 _29813_ (.A(_06452_),
    .X(_08186_));
 sky130_fd_sc_hd__and2_2 _29814_ (.A(_06815_),
    .B(_08186_),
    .X(_08187_));
 sky130_fd_sc_hd__nand2_2 _29815_ (.A(_08179_),
    .B(_08182_),
    .Y(_08188_));
 sky130_fd_sc_hd__nand3b_2 _29816_ (.A_N(_08185_),
    .B(_08187_),
    .C(_08188_),
    .Y(_08189_));
 sky130_fd_sc_hd__nand2_2 _29817_ (.A(_08184_),
    .B(_08189_),
    .Y(_08190_));
 sky130_fd_sc_hd__nand2_2 _29818_ (.A(_08177_),
    .B(_08190_),
    .Y(_08191_));
 sky130_fd_sc_hd__nand3b_2 _29819_ (.A_N(_08190_),
    .B(_08176_),
    .C(_08175_),
    .Y(_08192_));
 sky130_fd_sc_hd__nand2_2 _29820_ (.A(_08191_),
    .B(_08192_),
    .Y(_08193_));
 sky130_fd_sc_hd__nand2_2 _29821_ (.A(_08162_),
    .B(_08193_),
    .Y(_08194_));
 sky130_vsdinv _29822_ (.A(_08193_),
    .Y(_08195_));
 sky130_fd_sc_hd__buf_1 _29823_ (.A(_08161_),
    .X(_08196_));
 sky130_fd_sc_hd__nand3_2 _29824_ (.A(_08195_),
    .B(_08158_),
    .C(_08196_),
    .Y(_08197_));
 sky130_fd_sc_hd__a21oi_2 _29825_ (.A1(_08194_),
    .A2(_08197_),
    .B1(_08095_),
    .Y(_08198_));
 sky130_vsdinv _29826_ (.A(_08094_),
    .Y(_08199_));
 sky130_fd_sc_hd__a21oi_2 _29827_ (.A1(_08158_),
    .A2(_08196_),
    .B1(_08195_),
    .Y(_08200_));
 sky130_fd_sc_hd__a21oi_2 _29828_ (.A1(_08160_),
    .A2(_08154_),
    .B1(_08157_),
    .Y(_08201_));
 sky130_fd_sc_hd__nor3b_2 _29829_ (.A(_08193_),
    .B(_08201_),
    .C_N(_08196_),
    .Y(_08202_));
 sky130_fd_sc_hd__nor3_2 _29830_ (.A(_08199_),
    .B(_08200_),
    .C(_08202_),
    .Y(_08203_));
 sky130_fd_sc_hd__o21a_2 _29831_ (.A1(_08063_),
    .A2(_08066_),
    .B1(_08030_),
    .X(_08204_));
 sky130_vsdinv _29832_ (.A(_08204_),
    .Y(_08205_));
 sky130_fd_sc_hd__o21bai_2 _29833_ (.A1(_08198_),
    .A2(_08203_),
    .B1_N(_08205_),
    .Y(_08206_));
 sky130_fd_sc_hd__o21bai_2 _29834_ (.A1(_08200_),
    .A2(_08202_),
    .B1_N(_08094_),
    .Y(_08207_));
 sky130_fd_sc_hd__nand3_2 _29835_ (.A(_08194_),
    .B(_08095_),
    .C(_08197_),
    .Y(_08208_));
 sky130_fd_sc_hd__nand3_2 _29836_ (.A(_08207_),
    .B(_08205_),
    .C(_08208_),
    .Y(_08209_));
 sky130_fd_sc_hd__nand2_2 _29837_ (.A(_08206_),
    .B(_08209_),
    .Y(_08210_));
 sky130_vsdinv _29838_ (.A(_08090_),
    .Y(_08211_));
 sky130_fd_sc_hd__nand2_2 _29839_ (.A(_07533_),
    .B(_06820_),
    .Y(_08212_));
 sky130_fd_sc_hd__nand2_2 _29840_ (.A(_18764_),
    .B(_06826_),
    .Y(_08213_));
 sky130_fd_sc_hd__buf_1 _29841_ (.A(\pcpi_mul.rs2[19] ),
    .X(_08214_));
 sky130_fd_sc_hd__buf_1 _29842_ (.A(_08214_),
    .X(_08215_));
 sky130_fd_sc_hd__nand3b_2 _29843_ (.A_N(_08213_),
    .B(_08215_),
    .C(_05814_),
    .Y(_08216_));
 sky130_fd_sc_hd__buf_1 _29844_ (.A(_18763_),
    .X(_08217_));
 sky130_fd_sc_hd__buf_1 _29845_ (.A(_08217_),
    .X(_08218_));
 sky130_fd_sc_hd__buf_1 _29846_ (.A(_08218_),
    .X(_08219_));
 sky130_fd_sc_hd__buf_1 _29847_ (.A(_08215_),
    .X(_08220_));
 sky130_fd_sc_hd__a22o_2 _29848_ (.A1(_08219_),
    .A2(_05988_),
    .B1(_08220_),
    .B2(_05471_),
    .X(_08221_));
 sky130_fd_sc_hd__nand2_2 _29849_ (.A(_08216_),
    .B(_08221_),
    .Y(_08222_));
 sky130_fd_sc_hd__xnor2_2 _29850_ (.A(_08212_),
    .B(_08222_),
    .Y(_08223_));
 sky130_fd_sc_hd__buf_1 _29851_ (.A(_18752_),
    .X(_08224_));
 sky130_fd_sc_hd__nand2_2 _29852_ (.A(_08224_),
    .B(_05510_),
    .Y(_08225_));
 sky130_fd_sc_hd__buf_1 _29853_ (.A(_18747_),
    .X(_08226_));
 sky130_fd_sc_hd__nand2_2 _29854_ (.A(_08226_),
    .B(_19300_),
    .Y(_08227_));
 sky130_fd_sc_hd__nand2_2 _29855_ (.A(_08225_),
    .B(_08227_),
    .Y(_08228_));
 sky130_fd_sc_hd__nor2_2 _29856_ (.A(_08225_),
    .B(_08227_),
    .Y(_08229_));
 sky130_vsdinv _29857_ (.A(_08229_),
    .Y(_08230_));
 sky130_fd_sc_hd__buf_1 _29858_ (.A(_18759_),
    .X(_08231_));
 sky130_fd_sc_hd__buf_1 _29859_ (.A(_08231_),
    .X(_08232_));
 sky130_fd_sc_hd__o2bb2ai_2 _29860_ (.A1_N(_08228_),
    .A2_N(_08230_),
    .B1(_08232_),
    .B2(_19295_),
    .Y(_08233_));
 sky130_fd_sc_hd__buf_1 _29861_ (.A(\pcpi_mul.rs2[21] ),
    .X(_08234_));
 sky130_fd_sc_hd__buf_1 _29862_ (.A(_08234_),
    .X(_08235_));
 sky130_fd_sc_hd__and2_2 _29863_ (.A(_08235_),
    .B(_05984_),
    .X(_08236_));
 sky130_fd_sc_hd__nand3b_2 _29864_ (.A_N(_08229_),
    .B(_08236_),
    .C(_08228_),
    .Y(_08237_));
 sky130_fd_sc_hd__nor2_2 _29865_ (.A(_08083_),
    .B(_08087_),
    .Y(_08238_));
 sky130_fd_sc_hd__a21oi_2 _29866_ (.A1(_08233_),
    .A2(_08237_),
    .B1(_08238_),
    .Y(_08239_));
 sky130_fd_sc_hd__nand3_2 _29867_ (.A(_08233_),
    .B(_08238_),
    .C(_08237_),
    .Y(_08240_));
 sky130_vsdinv _29868_ (.A(_08240_),
    .Y(_08241_));
 sky130_fd_sc_hd__nor3_2 _29869_ (.A(_08223_),
    .B(_08239_),
    .C(_08241_),
    .Y(_08242_));
 sky130_fd_sc_hd__o21ai_2 _29870_ (.A1(_08239_),
    .A2(_08241_),
    .B1(_08223_),
    .Y(_08243_));
 sky130_fd_sc_hd__and2b_2 _29871_ (.A_N(_08242_),
    .B(_08243_),
    .X(_08244_));
 sky130_fd_sc_hd__xor2_2 _29872_ (.A(_08211_),
    .B(_08244_),
    .X(_08245_));
 sky130_vsdinv _29873_ (.A(_08245_),
    .Y(_08246_));
 sky130_fd_sc_hd__nand2_2 _29874_ (.A(_08210_),
    .B(_08246_),
    .Y(_08247_));
 sky130_fd_sc_hd__nand3_2 _29875_ (.A(_08206_),
    .B(_08245_),
    .C(_08209_),
    .Y(_08248_));
 sky130_fd_sc_hd__a21oi_2 _29876_ (.A1(_08247_),
    .A2(_08248_),
    .B1(_08099_),
    .Y(_08249_));
 sky130_fd_sc_hd__nand3_2 _29877_ (.A(_08247_),
    .B(_08099_),
    .C(_08248_),
    .Y(_08250_));
 sky130_vsdinv _29878_ (.A(_08250_),
    .Y(_08251_));
 sky130_fd_sc_hd__nor2_2 _29879_ (.A(_08249_),
    .B(_08251_),
    .Y(_08252_));
 sky130_fd_sc_hd__a22oi_2 _29880_ (.A1(_05982_),
    .A2(_06745_),
    .B1(_07697_),
    .B2(_07116_),
    .Y(_08253_));
 sky130_fd_sc_hd__buf_1 _29881_ (.A(_06733_),
    .X(_08254_));
 sky130_fd_sc_hd__buf_1 _29882_ (.A(_08254_),
    .X(_08255_));
 sky130_fd_sc_hd__buf_1 _29883_ (.A(_06744_),
    .X(_08256_));
 sky130_fd_sc_hd__and4_2 _29884_ (.A(_05772_),
    .B(_07556_),
    .C(_08255_),
    .D(_08256_),
    .X(_08257_));
 sky130_fd_sc_hd__buf_1 _29885_ (.A(_06935_),
    .X(_08258_));
 sky130_fd_sc_hd__and2_2 _29886_ (.A(_05778_),
    .B(_08258_),
    .X(_08259_));
 sky130_fd_sc_hd__o21bai_2 _29887_ (.A1(_08253_),
    .A2(_08257_),
    .B1_N(_08259_),
    .Y(_08260_));
 sky130_fd_sc_hd__buf_1 _29888_ (.A(\pcpi_mul.rs1[15] ),
    .X(_08261_));
 sky130_fd_sc_hd__buf_1 _29889_ (.A(_08261_),
    .X(_08262_));
 sky130_fd_sc_hd__nand2_2 _29890_ (.A(_07548_),
    .B(_08262_),
    .Y(_08263_));
 sky130_fd_sc_hd__nand3b_2 _29891_ (.A_N(_08263_),
    .B(_06890_),
    .C(_07329_),
    .Y(_08264_));
 sky130_fd_sc_hd__nand3b_2 _29892_ (.A_N(_08253_),
    .B(_08264_),
    .C(_08259_),
    .Y(_08265_));
 sky130_fd_sc_hd__nand2_2 _29893_ (.A(_08260_),
    .B(_08265_),
    .Y(_08266_));
 sky130_fd_sc_hd__a21oi_2 _29894_ (.A1(_08050_),
    .A2(_08055_),
    .B1(_08051_),
    .Y(_08267_));
 sky130_fd_sc_hd__nand2_2 _29895_ (.A(_08266_),
    .B(_08267_),
    .Y(_08268_));
 sky130_fd_sc_hd__nand3b_2 _29896_ (.A_N(_08267_),
    .B(_08260_),
    .C(_08265_),
    .Y(_08269_));
 sky130_fd_sc_hd__o31a_2 _29897_ (.A1(_06113_),
    .A2(_19217_),
    .A3(_07907_),
    .B1(_07914_),
    .X(_08270_));
 sky130_vsdinv _29898_ (.A(_08270_),
    .Y(_08271_));
 sky130_fd_sc_hd__a21oi_2 _29899_ (.A1(_08268_),
    .A2(_08269_),
    .B1(_08271_),
    .Y(_08272_));
 sky130_fd_sc_hd__nand3_2 _29900_ (.A(_08268_),
    .B(_08271_),
    .C(_08269_),
    .Y(_08273_));
 sky130_vsdinv _29901_ (.A(_08273_),
    .Y(_08274_));
 sky130_fd_sc_hd__o21ai_2 _29902_ (.A1(_08057_),
    .A2(_08047_),
    .B1(_08059_),
    .Y(_08275_));
 sky130_fd_sc_hd__o21bai_2 _29903_ (.A1(_08272_),
    .A2(_08274_),
    .B1_N(_08275_),
    .Y(_08276_));
 sky130_fd_sc_hd__nand2_2 _29904_ (.A(_08268_),
    .B(_08269_),
    .Y(_08277_));
 sky130_fd_sc_hd__nand2_2 _29905_ (.A(_08277_),
    .B(_08270_),
    .Y(_08278_));
 sky130_fd_sc_hd__nand3_2 _29906_ (.A(_08278_),
    .B(_08275_),
    .C(_08273_),
    .Y(_08279_));
 sky130_fd_sc_hd__a21boi_2 _29907_ (.A1(_07918_),
    .A2(_07922_),
    .B1_N(_07919_),
    .Y(_08280_));
 sky130_vsdinv _29908_ (.A(_08280_),
    .Y(_08281_));
 sky130_fd_sc_hd__a21oi_2 _29909_ (.A1(_08276_),
    .A2(_08279_),
    .B1(_08281_),
    .Y(_08282_));
 sky130_fd_sc_hd__nand3_2 _29910_ (.A(_08276_),
    .B(_08281_),
    .C(_08279_),
    .Y(_08283_));
 sky130_vsdinv _29911_ (.A(_08283_),
    .Y(_08284_));
 sky130_fd_sc_hd__a21oi_2 _29912_ (.A1(_07929_),
    .A2(_07924_),
    .B1(_07927_),
    .Y(_08285_));
 sky130_fd_sc_hd__o21ai_2 _29913_ (.A1(_07932_),
    .A2(_08285_),
    .B1(_07931_),
    .Y(_08286_));
 sky130_fd_sc_hd__o21bai_2 _29914_ (.A1(_08282_),
    .A2(_08284_),
    .B1_N(_08286_),
    .Y(_08287_));
 sky130_fd_sc_hd__a21o_2 _29915_ (.A1(_08276_),
    .A2(_08279_),
    .B1(_08281_),
    .X(_08288_));
 sky130_fd_sc_hd__nand3_2 _29916_ (.A(_08288_),
    .B(_08283_),
    .C(_08286_),
    .Y(_08289_));
 sky130_fd_sc_hd__nand2_2 _29917_ (.A(_05634_),
    .B(_07106_),
    .Y(_08290_));
 sky130_fd_sc_hd__buf_1 _29918_ (.A(_05642_),
    .X(_08291_));
 sky130_fd_sc_hd__buf_1 _29919_ (.A(_07309_),
    .X(_08292_));
 sky130_fd_sc_hd__nand2_2 _29920_ (.A(_08291_),
    .B(_08292_),
    .Y(_08293_));
 sky130_fd_sc_hd__nor2_2 _29921_ (.A(_08290_),
    .B(_08293_),
    .Y(_08294_));
 sky130_fd_sc_hd__buf_1 _29922_ (.A(_19179_),
    .X(_08295_));
 sky130_fd_sc_hd__and2_2 _29923_ (.A(_06732_),
    .B(_08295_),
    .X(_08296_));
 sky130_fd_sc_hd__nand2_2 _29924_ (.A(_08290_),
    .B(_08293_),
    .Y(_08297_));
 sky130_fd_sc_hd__nand3b_2 _29925_ (.A_N(_08294_),
    .B(_08296_),
    .C(_08297_),
    .Y(_08298_));
 sky130_fd_sc_hd__buf_1 _29926_ (.A(_07324_),
    .X(_08299_));
 sky130_fd_sc_hd__buf_1 _29927_ (.A(_08299_),
    .X(_08300_));
 sky130_fd_sc_hd__buf_1 _29928_ (.A(_08300_),
    .X(_08301_));
 sky130_fd_sc_hd__buf_1 _29929_ (.A(_19202_),
    .X(_08302_));
 sky130_fd_sc_hd__buf_1 _29930_ (.A(_08302_),
    .X(_08303_));
 sky130_fd_sc_hd__buf_1 _29931_ (.A(_08303_),
    .X(_08304_));
 sky130_fd_sc_hd__a22oi_2 _29932_ (.A1(_18845_),
    .A2(_08301_),
    .B1(_18851_),
    .B2(_08304_),
    .Y(_08305_));
 sky130_fd_sc_hd__o21bai_2 _29933_ (.A1(_08305_),
    .A2(_08294_),
    .B1_N(_08296_),
    .Y(_08306_));
 sky130_fd_sc_hd__nand2_2 _29934_ (.A(_07954_),
    .B(_07949_),
    .Y(_08307_));
 sky130_fd_sc_hd__a21o_2 _29935_ (.A1(_08298_),
    .A2(_08306_),
    .B1(_08307_),
    .X(_08308_));
 sky130_fd_sc_hd__nand3_2 _29936_ (.A(_08307_),
    .B(_08298_),
    .C(_08306_),
    .Y(_08309_));
 sky130_fd_sc_hd__buf_1 _29937_ (.A(_07733_),
    .X(_08310_));
 sky130_fd_sc_hd__nand2_2 _29938_ (.A(_05953_),
    .B(_08310_),
    .Y(_08311_));
 sky130_fd_sc_hd__nand2_2 _29939_ (.A(_05554_),
    .B(_07952_),
    .Y(_08312_));
 sky130_fd_sc_hd__xor2_2 _29940_ (.A(_08311_),
    .B(_08312_),
    .X(_08313_));
 sky130_fd_sc_hd__buf_1 _29941_ (.A(_07961_),
    .X(_08314_));
 sky130_fd_sc_hd__and2_2 _29942_ (.A(_06460_),
    .B(_08314_),
    .X(_08315_));
 sky130_fd_sc_hd__nand2_2 _29943_ (.A(_08313_),
    .B(_08315_),
    .Y(_08316_));
 sky130_fd_sc_hd__xnor2_2 _29944_ (.A(_08311_),
    .B(_08312_),
    .Y(_08317_));
 sky130_fd_sc_hd__o21ai_2 _29945_ (.A1(_06923_),
    .A2(_19198_),
    .B1(_08317_),
    .Y(_08318_));
 sky130_fd_sc_hd__nand2_2 _29946_ (.A(_08316_),
    .B(_08318_),
    .Y(_08319_));
 sky130_fd_sc_hd__a21boi_2 _29947_ (.A1(_08308_),
    .A2(_08309_),
    .B1_N(_08319_),
    .Y(_08320_));
 sky130_fd_sc_hd__nand3b_2 _29948_ (.A_N(_08319_),
    .B(_08308_),
    .C(_08309_),
    .Y(_08321_));
 sky130_vsdinv _29949_ (.A(_08321_),
    .Y(_08322_));
 sky130_fd_sc_hd__o21ai_2 _29950_ (.A1(_07973_),
    .A2(_07975_),
    .B1(_07959_),
    .Y(_08323_));
 sky130_fd_sc_hd__o21bai_2 _29951_ (.A1(_08320_),
    .A2(_08322_),
    .B1_N(_08323_),
    .Y(_08324_));
 sky130_fd_sc_hd__nand3b_2 _29952_ (.A_N(_08320_),
    .B(_08321_),
    .C(_08323_),
    .Y(_08325_));
 sky130_fd_sc_hd__o21a_2 _29953_ (.A1(_07962_),
    .A2(_07964_),
    .B1(_07969_),
    .X(_08326_));
 sky130_vsdinv _29954_ (.A(_08326_),
    .Y(_08327_));
 sky130_fd_sc_hd__a21oi_2 _29955_ (.A1(_08324_),
    .A2(_08325_),
    .B1(_08327_),
    .Y(_08328_));
 sky130_fd_sc_hd__nand3_2 _29956_ (.A(_08324_),
    .B(_08327_),
    .C(_08325_),
    .Y(_08329_));
 sky130_vsdinv _29957_ (.A(_08329_),
    .Y(_08330_));
 sky130_fd_sc_hd__nor2_2 _29958_ (.A(_08328_),
    .B(_08330_),
    .Y(_08331_));
 sky130_fd_sc_hd__a21oi_2 _29959_ (.A1(_08287_),
    .A2(_08289_),
    .B1(_08331_),
    .Y(_08332_));
 sky130_fd_sc_hd__or2b_2 _29960_ (.A(_08328_),
    .B_N(_08329_),
    .X(_08333_));
 sky130_fd_sc_hd__nand2_2 _29961_ (.A(_08287_),
    .B(_08289_),
    .Y(_08334_));
 sky130_fd_sc_hd__nor2_2 _29962_ (.A(_08333_),
    .B(_08334_),
    .Y(_08335_));
 sky130_vsdinv _29963_ (.A(_08073_),
    .Y(_08336_));
 sky130_fd_sc_hd__o21bai_2 _29964_ (.A1(_08332_),
    .A2(_08335_),
    .B1_N(_08336_),
    .Y(_08337_));
 sky130_fd_sc_hd__a21boi_2 _29965_ (.A1(_07989_),
    .A2(_07938_),
    .B1_N(_07941_),
    .Y(_08338_));
 sky130_vsdinv _29966_ (.A(_08338_),
    .Y(_08339_));
 sky130_fd_sc_hd__nand2_2 _29967_ (.A(_08334_),
    .B(_08333_),
    .Y(_08340_));
 sky130_fd_sc_hd__nand3_2 _29968_ (.A(_08331_),
    .B(_08287_),
    .C(_08289_),
    .Y(_08341_));
 sky130_fd_sc_hd__nand3_2 _29969_ (.A(_08340_),
    .B(_08336_),
    .C(_08341_),
    .Y(_08342_));
 sky130_fd_sc_hd__nand3_2 _29970_ (.A(_08337_),
    .B(_08339_),
    .C(_08342_),
    .Y(_08343_));
 sky130_fd_sc_hd__buf_1 _29971_ (.A(_08343_),
    .X(_08344_));
 sky130_fd_sc_hd__a21oi_2 _29972_ (.A1(_08340_),
    .A2(_08341_),
    .B1(_08336_),
    .Y(_08345_));
 sky130_fd_sc_hd__nor3_2 _29973_ (.A(_08073_),
    .B(_08332_),
    .C(_08335_),
    .Y(_08346_));
 sky130_fd_sc_hd__o21bai_2 _29974_ (.A1(_08345_),
    .A2(_08346_),
    .B1_N(_08339_),
    .Y(_08347_));
 sky130_fd_sc_hd__buf_1 _29975_ (.A(_08347_),
    .X(_08348_));
 sky130_fd_sc_hd__nand3_2 _29976_ (.A(_08252_),
    .B(_08344_),
    .C(_08348_),
    .Y(_08349_));
 sky130_fd_sc_hd__nand2_2 _29977_ (.A(_08347_),
    .B(_08343_),
    .Y(_08350_));
 sky130_fd_sc_hd__a21oi_2 _29978_ (.A1(_08206_),
    .A2(_08209_),
    .B1(_08245_),
    .Y(_08351_));
 sky130_fd_sc_hd__a21oi_2 _29979_ (.A1(_08207_),
    .A2(_08208_),
    .B1(_08205_),
    .Y(_08352_));
 sky130_fd_sc_hd__nor3b_2 _29980_ (.A(_08246_),
    .B(_08352_),
    .C_N(_08209_),
    .Y(_08353_));
 sky130_fd_sc_hd__o21bai_2 _29981_ (.A1(_08351_),
    .A2(_08353_),
    .B1_N(_08099_),
    .Y(_08354_));
 sky130_fd_sc_hd__nand2_2 _29982_ (.A(_08354_),
    .B(_08250_),
    .Y(_08355_));
 sky130_fd_sc_hd__nand2_2 _29983_ (.A(_08350_),
    .B(_08355_),
    .Y(_08356_));
 sky130_vsdinv _29984_ (.A(_08100_),
    .Y(_08357_));
 sky130_fd_sc_hd__nand2_2 _29985_ (.A(_08105_),
    .B(_08357_),
    .Y(_08358_));
 sky130_fd_sc_hd__nand3_2 _29986_ (.A(_08349_),
    .B(_08356_),
    .C(_08358_),
    .Y(_08359_));
 sky130_fd_sc_hd__buf_1 _29987_ (.A(_08359_),
    .X(_08360_));
 sky130_fd_sc_hd__a22oi_2 _29988_ (.A1(_08354_),
    .A2(_08250_),
    .B1(_08348_),
    .B2(_08344_),
    .Y(_08361_));
 sky130_fd_sc_hd__nor2_2 _29989_ (.A(_08355_),
    .B(_08350_),
    .Y(_08362_));
 sky130_fd_sc_hd__o21bai_2 _29990_ (.A1(_08361_),
    .A2(_08362_),
    .B1_N(_08358_),
    .Y(_08363_));
 sky130_fd_sc_hd__a21boi_2 _29991_ (.A1(_07979_),
    .A2(_07985_),
    .B1_N(_07983_),
    .Y(_08364_));
 sky130_fd_sc_hd__a21oi_2 _29992_ (.A1(_07999_),
    .A2(_07998_),
    .B1(_08364_),
    .Y(_08365_));
 sky130_fd_sc_hd__and3_2 _29993_ (.A(_07999_),
    .B(_07998_),
    .C(_08364_),
    .X(_08366_));
 sky130_fd_sc_hd__o2bb2ai_2 _29994_ (.A1_N(_08360_),
    .A2_N(_08363_),
    .B1(_08365_),
    .B2(_08366_),
    .Y(_08367_));
 sky130_fd_sc_hd__a21o_2 _29995_ (.A1(_07994_),
    .A2(_07995_),
    .B1(_08001_),
    .X(_08368_));
 sky130_fd_sc_hd__xnor2_2 _29996_ (.A(_08364_),
    .B(_08368_),
    .Y(_08369_));
 sky130_fd_sc_hd__nand3_2 _29997_ (.A(_08363_),
    .B(_08359_),
    .C(_08369_),
    .Y(_08370_));
 sky130_fd_sc_hd__nand3_2 _29998_ (.A(_08135_),
    .B(_08367_),
    .C(_08370_),
    .Y(_08371_));
 sky130_fd_sc_hd__a21oi_2 _29999_ (.A1(_08363_),
    .A2(_08360_),
    .B1(_08369_),
    .Y(_08372_));
 sky130_vsdinv _30000_ (.A(_08370_),
    .Y(_08373_));
 sky130_fd_sc_hd__o21bai_2 _30001_ (.A1(_08372_),
    .A2(_08373_),
    .B1_N(_08135_),
    .Y(_08374_));
 sky130_fd_sc_hd__o2bb2ai_2 _30002_ (.A1_N(_08371_),
    .A2_N(_08374_),
    .B1(_08112_),
    .B2(_08111_),
    .Y(_08375_));
 sky130_fd_sc_hd__a21oi_2 _30003_ (.A1(_07869_),
    .A2(_07780_),
    .B1(_08111_),
    .Y(_08376_));
 sky130_fd_sc_hd__nand3_2 _30004_ (.A(_08374_),
    .B(_08376_),
    .C(_08371_),
    .Y(_08377_));
 sky130_fd_sc_hd__nand2_2 _30005_ (.A(_08124_),
    .B(_08121_),
    .Y(_08378_));
 sky130_fd_sc_hd__a21oi_2 _30006_ (.A1(_08375_),
    .A2(_08377_),
    .B1(_08378_),
    .Y(_08379_));
 sky130_fd_sc_hd__a21boi_2 _30007_ (.A1(_08118_),
    .A2(_08122_),
    .B1_N(_08121_),
    .Y(_08380_));
 sky130_fd_sc_hd__a21oi_2 _30008_ (.A1(_08374_),
    .A2(_08371_),
    .B1(_08376_),
    .Y(_08381_));
 sky130_fd_sc_hd__nor3b_2 _30009_ (.A(_08380_),
    .B(_08381_),
    .C_N(_08377_),
    .Y(_08382_));
 sky130_fd_sc_hd__nor2_2 _30010_ (.A(_08379_),
    .B(_08382_),
    .Y(_08383_));
 sky130_fd_sc_hd__o21bai_2 _30011_ (.A1(_08126_),
    .A2(_08134_),
    .B1_N(_08129_),
    .Y(_08384_));
 sky130_fd_sc_hd__xor2_2 _30012_ (.A(_08383_),
    .B(_08384_),
    .X(_02642_));
 sky130_fd_sc_hd__a22oi_2 _30013_ (.A1(_07786_),
    .A2(_08007_),
    .B1(_07470_),
    .B2(_05841_),
    .Y(_08385_));
 sky130_fd_sc_hd__nand2_2 _30014_ (.A(_07785_),
    .B(_06979_),
    .Y(_08386_));
 sky130_fd_sc_hd__nand2_2 _30015_ (.A(_08012_),
    .B(_05846_),
    .Y(_08387_));
 sky130_fd_sc_hd__nor2_2 _30016_ (.A(_08386_),
    .B(_08387_),
    .Y(_08388_));
 sky130_fd_sc_hd__and2_2 _30017_ (.A(_18790_),
    .B(_05821_),
    .X(_08389_));
 sky130_fd_sc_hd__o21bai_2 _30018_ (.A1(_08385_),
    .A2(_08388_),
    .B1_N(_08389_),
    .Y(_08390_));
 sky130_fd_sc_hd__buf_1 _30019_ (.A(_07787_),
    .X(_08391_));
 sky130_fd_sc_hd__nand3b_2 _30020_ (.A_N(_08386_),
    .B(_08391_),
    .C(_06181_),
    .Y(_08392_));
 sky130_fd_sc_hd__nand2_2 _30021_ (.A(_08386_),
    .B(_08387_),
    .Y(_08393_));
 sky130_fd_sc_hd__nand3_2 _30022_ (.A(_08392_),
    .B(_08389_),
    .C(_08393_),
    .Y(_08394_));
 sky130_fd_sc_hd__nand2_2 _30023_ (.A(_08390_),
    .B(_08394_),
    .Y(_08395_));
 sky130_fd_sc_hd__a22oi_2 _30024_ (.A1(_08074_),
    .A2(_05540_),
    .B1(_07853_),
    .B2(_05555_),
    .Y(_08396_));
 sky130_fd_sc_hd__o21ai_2 _30025_ (.A1(_08212_),
    .A2(_08396_),
    .B1(_08216_),
    .Y(_08397_));
 sky130_vsdinv _30026_ (.A(_08397_),
    .Y(_08398_));
 sky130_fd_sc_hd__nand2_2 _30027_ (.A(_08395_),
    .B(_08398_),
    .Y(_08399_));
 sky130_fd_sc_hd__nand3_2 _30028_ (.A(_08390_),
    .B(_08397_),
    .C(_08394_),
    .Y(_08400_));
 sky130_fd_sc_hd__a21oi_2 _30029_ (.A1(_08144_),
    .A2(_08140_),
    .B1(_08139_),
    .Y(_08401_));
 sky130_vsdinv _30030_ (.A(_08401_),
    .Y(_08402_));
 sky130_fd_sc_hd__a21oi_2 _30031_ (.A1(_08399_),
    .A2(_08400_),
    .B1(_08402_),
    .Y(_08403_));
 sky130_fd_sc_hd__a21oi_2 _30032_ (.A1(_08390_),
    .A2(_08394_),
    .B1(_08397_),
    .Y(_08404_));
 sky130_vsdinv _30033_ (.A(_08400_),
    .Y(_08405_));
 sky130_fd_sc_hd__nor3_2 _30034_ (.A(_08401_),
    .B(_08404_),
    .C(_08405_),
    .Y(_08406_));
 sky130_fd_sc_hd__a21oi_2 _30035_ (.A1(_08141_),
    .A2(_08145_),
    .B1(_08147_),
    .Y(_08407_));
 sky130_fd_sc_hd__o21ai_2 _30036_ (.A1(_08151_),
    .A2(_08407_),
    .B1(_08150_),
    .Y(_08408_));
 sky130_fd_sc_hd__o21bai_2 _30037_ (.A1(_08403_),
    .A2(_08406_),
    .B1_N(_08408_),
    .Y(_08409_));
 sky130_fd_sc_hd__o21bai_2 _30038_ (.A1(_08404_),
    .A2(_08405_),
    .B1_N(_08402_),
    .Y(_08410_));
 sky130_fd_sc_hd__nand3_2 _30039_ (.A(_08399_),
    .B(_08402_),
    .C(_08400_),
    .Y(_08411_));
 sky130_fd_sc_hd__nand3_2 _30040_ (.A(_08410_),
    .B(_08411_),
    .C(_08408_),
    .Y(_08412_));
 sky130_fd_sc_hd__nand2_2 _30041_ (.A(_08409_),
    .B(_08412_),
    .Y(_08413_));
 sky130_fd_sc_hd__buf_1 _30042_ (.A(_06543_),
    .X(_08414_));
 sky130_fd_sc_hd__nand2_2 _30043_ (.A(_08414_),
    .B(_06063_),
    .Y(_08415_));
 sky130_fd_sc_hd__nand2_2 _30044_ (.A(_18802_),
    .B(_06886_),
    .Y(_08416_));
 sky130_fd_sc_hd__nor2_2 _30045_ (.A(_08415_),
    .B(_08416_),
    .Y(_08417_));
 sky130_fd_sc_hd__and2_2 _30046_ (.A(_18808_),
    .B(_06187_),
    .X(_08418_));
 sky130_fd_sc_hd__nand2_2 _30047_ (.A(_08415_),
    .B(_08416_),
    .Y(_08419_));
 sky130_fd_sc_hd__nand3b_2 _30048_ (.A_N(_08417_),
    .B(_08418_),
    .C(_08419_),
    .Y(_08420_));
 sky130_fd_sc_hd__a22oi_2 _30049_ (.A1(_08170_),
    .A2(_06444_),
    .B1(_06393_),
    .B2(_06197_),
    .Y(_08421_));
 sky130_fd_sc_hd__o21bai_2 _30050_ (.A1(_08421_),
    .A2(_08417_),
    .B1_N(_08418_),
    .Y(_08422_));
 sky130_fd_sc_hd__a21oi_2 _30051_ (.A1(_08167_),
    .A2(_08166_),
    .B1(_08165_),
    .Y(_08423_));
 sky130_fd_sc_hd__a21boi_2 _30052_ (.A1(_08420_),
    .A2(_08422_),
    .B1_N(_08423_),
    .Y(_08424_));
 sky130_fd_sc_hd__nand3b_2 _30053_ (.A_N(_08423_),
    .B(_08420_),
    .C(_08422_),
    .Y(_08425_));
 sky130_vsdinv _30054_ (.A(_08425_),
    .Y(_08426_));
 sky130_fd_sc_hd__nand2_2 _30055_ (.A(_08178_),
    .B(_06350_),
    .Y(_08427_));
 sky130_fd_sc_hd__nand2_2 _30056_ (.A(_08180_),
    .B(_07698_),
    .Y(_08428_));
 sky130_fd_sc_hd__nand2_2 _30057_ (.A(_08427_),
    .B(_08428_),
    .Y(_08429_));
 sky130_fd_sc_hd__nor2_2 _30058_ (.A(_08427_),
    .B(_08428_),
    .Y(_08430_));
 sky130_vsdinv _30059_ (.A(_08430_),
    .Y(_08431_));
 sky130_fd_sc_hd__o2bb2ai_2 _30060_ (.A1_N(_08429_),
    .A2_N(_08431_),
    .B1(_07818_),
    .B2(_19228_),
    .Y(_08432_));
 sky130_fd_sc_hd__and2_2 _30061_ (.A(_06815_),
    .B(_06595_),
    .X(_08433_));
 sky130_fd_sc_hd__nand3b_2 _30062_ (.A_N(_08430_),
    .B(_08433_),
    .C(_08429_),
    .Y(_08434_));
 sky130_fd_sc_hd__nand2_2 _30063_ (.A(_08432_),
    .B(_08434_),
    .Y(_08435_));
 sky130_fd_sc_hd__o21ai_2 _30064_ (.A1(_08424_),
    .A2(_08426_),
    .B1(_08435_),
    .Y(_08436_));
 sky130_fd_sc_hd__a21bo_2 _30065_ (.A1(_08420_),
    .A2(_08422_),
    .B1_N(_08423_),
    .X(_08437_));
 sky130_fd_sc_hd__nand3b_2 _30066_ (.A_N(_08435_),
    .B(_08425_),
    .C(_08437_),
    .Y(_08438_));
 sky130_fd_sc_hd__nand2_2 _30067_ (.A(_08436_),
    .B(_08438_),
    .Y(_08439_));
 sky130_fd_sc_hd__buf_1 _30068_ (.A(_08439_),
    .X(_08440_));
 sky130_fd_sc_hd__nand2_2 _30069_ (.A(_08413_),
    .B(_08440_),
    .Y(_08441_));
 sky130_fd_sc_hd__buf_1 _30070_ (.A(_08412_),
    .X(_08442_));
 sky130_fd_sc_hd__nand3b_2 _30071_ (.A_N(_08439_),
    .B(_08409_),
    .C(_08442_),
    .Y(_08443_));
 sky130_fd_sc_hd__nand3b_2 _30072_ (.A_N(_08242_),
    .B(_08211_),
    .C(_08243_),
    .Y(_08444_));
 sky130_fd_sc_hd__a21boi_2 _30073_ (.A1(_08441_),
    .A2(_08443_),
    .B1_N(_08444_),
    .Y(_08445_));
 sky130_fd_sc_hd__a21boi_2 _30074_ (.A1(_08409_),
    .A2(_08442_),
    .B1_N(_08440_),
    .Y(_08446_));
 sky130_fd_sc_hd__a21oi_2 _30075_ (.A1(_08410_),
    .A2(_08411_),
    .B1(_08408_),
    .Y(_08447_));
 sky130_vsdinv _30076_ (.A(_08442_),
    .Y(_08448_));
 sky130_fd_sc_hd__nor3_2 _30077_ (.A(_08440_),
    .B(_08447_),
    .C(_08448_),
    .Y(_08449_));
 sky130_fd_sc_hd__nor3_2 _30078_ (.A(_08444_),
    .B(_08446_),
    .C(_08449_),
    .Y(_08450_));
 sky130_fd_sc_hd__o21a_2 _30079_ (.A1(_08193_),
    .A2(_08201_),
    .B1(_08196_),
    .X(_08451_));
 sky130_vsdinv _30080_ (.A(_08451_),
    .Y(_08452_));
 sky130_fd_sc_hd__o21bai_2 _30081_ (.A1(_08445_),
    .A2(_08450_),
    .B1_N(_08452_),
    .Y(_08453_));
 sky130_fd_sc_hd__o21ai_2 _30082_ (.A1(_08446_),
    .A2(_08449_),
    .B1(_08444_),
    .Y(_08454_));
 sky130_fd_sc_hd__nand3b_2 _30083_ (.A_N(_08444_),
    .B(_08441_),
    .C(_08443_),
    .Y(_08455_));
 sky130_fd_sc_hd__nand3_2 _30084_ (.A(_08454_),
    .B(_08452_),
    .C(_08455_),
    .Y(_08456_));
 sky130_fd_sc_hd__buf_1 _30085_ (.A(\pcpi_mul.rs2[24] ),
    .X(_08457_));
 sky130_fd_sc_hd__buf_1 _30086_ (.A(_08457_),
    .X(_08458_));
 sky130_fd_sc_hd__buf_1 _30087_ (.A(_08458_),
    .X(_08459_));
 sky130_fd_sc_hd__buf_1 _30088_ (.A(_08459_),
    .X(_08460_));
 sky130_fd_sc_hd__and2_2 _30089_ (.A(_08460_),
    .B(_05589_),
    .X(_08461_));
 sky130_fd_sc_hd__buf_1 _30090_ (.A(\pcpi_mul.rs2[23] ),
    .X(_08462_));
 sky130_fd_sc_hd__buf_1 _30091_ (.A(_08462_),
    .X(_08463_));
 sky130_fd_sc_hd__nand2_2 _30092_ (.A(_08463_),
    .B(_05423_),
    .Y(_08464_));
 sky130_fd_sc_hd__buf_1 _30093_ (.A(\pcpi_mul.rs2[22] ),
    .X(_08465_));
 sky130_fd_sc_hd__nand2_2 _30094_ (.A(_08465_),
    .B(_05430_),
    .Y(_08466_));
 sky130_fd_sc_hd__nor2_2 _30095_ (.A(_08464_),
    .B(_08466_),
    .Y(_08467_));
 sky130_fd_sc_hd__and2_2 _30096_ (.A(_07844_),
    .B(_07171_),
    .X(_08468_));
 sky130_fd_sc_hd__nand2_2 _30097_ (.A(_08464_),
    .B(_08466_),
    .Y(_08469_));
 sky130_fd_sc_hd__nand3b_2 _30098_ (.A_N(_08467_),
    .B(_08468_),
    .C(_08469_),
    .Y(_08470_));
 sky130_fd_sc_hd__buf_1 _30099_ (.A(\pcpi_mul.rs2[23] ),
    .X(_08471_));
 sky130_fd_sc_hd__buf_1 _30100_ (.A(_08471_),
    .X(_08472_));
 sky130_fd_sc_hd__buf_1 _30101_ (.A(_08465_),
    .X(_08473_));
 sky130_fd_sc_hd__a22oi_2 _30102_ (.A1(_08472_),
    .A2(_06143_),
    .B1(_08473_),
    .B2(_05636_),
    .Y(_08474_));
 sky130_fd_sc_hd__o21bai_2 _30103_ (.A1(_08474_),
    .A2(_08467_),
    .B1_N(_08468_),
    .Y(_08475_));
 sky130_fd_sc_hd__a21o_2 _30104_ (.A1(_08228_),
    .A2(_08236_),
    .B1(_08229_),
    .X(_08476_));
 sky130_fd_sc_hd__nand3_2 _30105_ (.A(_08470_),
    .B(_08475_),
    .C(_08476_),
    .Y(_08477_));
 sky130_fd_sc_hd__nand2_2 _30106_ (.A(_08470_),
    .B(_08475_),
    .Y(_08478_));
 sky130_fd_sc_hd__nand3_2 _30107_ (.A(_08478_),
    .B(_08230_),
    .C(_08237_),
    .Y(_08479_));
 sky130_fd_sc_hd__buf_1 _30108_ (.A(_05664_),
    .X(_08480_));
 sky130_fd_sc_hd__nand2_2 _30109_ (.A(_07532_),
    .B(_08480_),
    .Y(_08481_));
 sky130_fd_sc_hd__nand2_2 _30110_ (.A(_08217_),
    .B(_05469_),
    .Y(_08482_));
 sky130_fd_sc_hd__nand2_2 _30111_ (.A(_08214_),
    .B(_19277_),
    .Y(_08483_));
 sky130_fd_sc_hd__nor2_2 _30112_ (.A(_08482_),
    .B(_08483_),
    .Y(_08484_));
 sky130_fd_sc_hd__nand2_2 _30113_ (.A(_08482_),
    .B(_08483_),
    .Y(_08485_));
 sky130_fd_sc_hd__nor3b_2 _30114_ (.A(_08481_),
    .B(_08484_),
    .C_N(_08485_),
    .Y(_08486_));
 sky130_vsdinv _30115_ (.A(_08484_),
    .Y(_08487_));
 sky130_vsdinv _30116_ (.A(_08481_),
    .Y(_08488_));
 sky130_fd_sc_hd__a21oi_2 _30117_ (.A1(_08487_),
    .A2(_08485_),
    .B1(_08488_),
    .Y(_08489_));
 sky130_fd_sc_hd__o2bb2ai_2 _30118_ (.A1_N(_08477_),
    .A2_N(_08479_),
    .B1(_08486_),
    .B2(_08489_),
    .Y(_08490_));
 sky130_fd_sc_hd__nor2_2 _30119_ (.A(_08486_),
    .B(_08489_),
    .Y(_08491_));
 sky130_fd_sc_hd__nand3_2 _30120_ (.A(_08479_),
    .B(_08491_),
    .C(_08477_),
    .Y(_08492_));
 sky130_fd_sc_hd__o21ai_2 _30121_ (.A1(_08223_),
    .A2(_08239_),
    .B1(_08240_),
    .Y(_08493_));
 sky130_fd_sc_hd__a21o_2 _30122_ (.A1(_08490_),
    .A2(_08492_),
    .B1(_08493_),
    .X(_08494_));
 sky130_fd_sc_hd__nand3_2 _30123_ (.A(_08493_),
    .B(_08490_),
    .C(_08492_),
    .Y(_08495_));
 sky130_fd_sc_hd__nand2_2 _30124_ (.A(_08494_),
    .B(_08495_),
    .Y(_08496_));
 sky130_fd_sc_hd__xor2_2 _30125_ (.A(_08461_),
    .B(_08496_),
    .X(_08497_));
 sky130_vsdinv _30126_ (.A(_08497_),
    .Y(_08498_));
 sky130_fd_sc_hd__a21oi_2 _30127_ (.A1(_08453_),
    .A2(_08456_),
    .B1(_08498_),
    .Y(_08499_));
 sky130_fd_sc_hd__a21oi_2 _30128_ (.A1(_08454_),
    .A2(_08455_),
    .B1(_08452_),
    .Y(_08500_));
 sky130_vsdinv _30129_ (.A(_08456_),
    .Y(_08501_));
 sky130_fd_sc_hd__nor3_2 _30130_ (.A(_08497_),
    .B(_08500_),
    .C(_08501_),
    .Y(_08502_));
 sky130_fd_sc_hd__o22ai_2 _30131_ (.A1(_08246_),
    .A2(_08210_),
    .B1(_08499_),
    .B2(_08502_),
    .Y(_08503_));
 sky130_fd_sc_hd__nand2_2 _30132_ (.A(_08453_),
    .B(_08456_),
    .Y(_08504_));
 sky130_fd_sc_hd__nand2_2 _30133_ (.A(_08504_),
    .B(_08497_),
    .Y(_08505_));
 sky130_fd_sc_hd__nand3_2 _30134_ (.A(_08453_),
    .B(_08498_),
    .C(_08456_),
    .Y(_08506_));
 sky130_fd_sc_hd__nand3b_2 _30135_ (.A_N(_08248_),
    .B(_08505_),
    .C(_08506_),
    .Y(_08507_));
 sky130_vsdinv _30136_ (.A(_08289_),
    .Y(_08508_));
 sky130_fd_sc_hd__a21oi_2 _30137_ (.A1(_08331_),
    .A2(_08287_),
    .B1(_08508_),
    .Y(_08509_));
 sky130_fd_sc_hd__buf_1 _30138_ (.A(_19215_),
    .X(_08510_));
 sky130_fd_sc_hd__a22oi_2 _30139_ (.A1(_06224_),
    .A2(_08510_),
    .B1(_07556_),
    .B2(_07947_),
    .Y(_08511_));
 sky130_fd_sc_hd__nand2_2 _30140_ (.A(_05771_),
    .B(_08254_),
    .Y(_08512_));
 sky130_fd_sc_hd__nand2_2 _30141_ (.A(_05872_),
    .B(_06936_),
    .Y(_08513_));
 sky130_fd_sc_hd__nor2_2 _30142_ (.A(_08512_),
    .B(_08513_),
    .Y(_08514_));
 sky130_fd_sc_hd__and2_2 _30143_ (.A(_06100_),
    .B(_07105_),
    .X(_08515_));
 sky130_fd_sc_hd__o21bai_2 _30144_ (.A1(_08511_),
    .A2(_08514_),
    .B1_N(_08515_),
    .Y(_08516_));
 sky130_fd_sc_hd__nand3b_2 _30145_ (.A_N(_08512_),
    .B(_07697_),
    .C(_07737_),
    .Y(_08517_));
 sky130_fd_sc_hd__nand2_2 _30146_ (.A(_08512_),
    .B(_08513_),
    .Y(_08518_));
 sky130_fd_sc_hd__nand3_2 _30147_ (.A(_08517_),
    .B(_08515_),
    .C(_08518_),
    .Y(_08519_));
 sky130_fd_sc_hd__nand2_2 _30148_ (.A(_08516_),
    .B(_08519_),
    .Y(_08520_));
 sky130_fd_sc_hd__a21oi_2 _30149_ (.A1(_08188_),
    .A2(_08187_),
    .B1(_08185_),
    .Y(_08521_));
 sky130_fd_sc_hd__nand2_2 _30150_ (.A(_08520_),
    .B(_08521_),
    .Y(_08522_));
 sky130_fd_sc_hd__nand3b_2 _30151_ (.A_N(_08521_),
    .B(_08519_),
    .C(_08516_),
    .Y(_08523_));
 sky130_fd_sc_hd__buf_1 _30152_ (.A(_19212_),
    .X(_08524_));
 sky130_fd_sc_hd__o31a_2 _30153_ (.A1(_06113_),
    .A2(_08524_),
    .A3(_08253_),
    .B1(_08264_),
    .X(_08525_));
 sky130_vsdinv _30154_ (.A(_08525_),
    .Y(_08526_));
 sky130_fd_sc_hd__a21oi_2 _30155_ (.A1(_08522_),
    .A2(_08523_),
    .B1(_08526_),
    .Y(_08527_));
 sky130_fd_sc_hd__nand2_2 _30156_ (.A(_08522_),
    .B(_08523_),
    .Y(_08528_));
 sky130_fd_sc_hd__nor2_2 _30157_ (.A(_08525_),
    .B(_08528_),
    .Y(_08529_));
 sky130_fd_sc_hd__a21boi_2 _30158_ (.A1(_08168_),
    .A2(_08172_),
    .B1_N(_08174_),
    .Y(_08530_));
 sky130_fd_sc_hd__o21ai_2 _30159_ (.A1(_08190_),
    .A2(_08530_),
    .B1(_08176_),
    .Y(_08531_));
 sky130_fd_sc_hd__o21bai_2 _30160_ (.A1(_08527_),
    .A2(_08529_),
    .B1_N(_08531_),
    .Y(_08532_));
 sky130_fd_sc_hd__nand2_2 _30161_ (.A(_08528_),
    .B(_08525_),
    .Y(_08533_));
 sky130_fd_sc_hd__nand3_2 _30162_ (.A(_08522_),
    .B(_08526_),
    .C(_08523_),
    .Y(_08534_));
 sky130_fd_sc_hd__nand3_2 _30163_ (.A(_08531_),
    .B(_08533_),
    .C(_08534_),
    .Y(_08535_));
 sky130_fd_sc_hd__buf_1 _30164_ (.A(_08535_),
    .X(_08536_));
 sky130_fd_sc_hd__a21boi_2 _30165_ (.A1(_08268_),
    .A2(_08271_),
    .B1_N(_08269_),
    .Y(_08537_));
 sky130_vsdinv _30166_ (.A(_08537_),
    .Y(_08538_));
 sky130_fd_sc_hd__a21oi_2 _30167_ (.A1(_08532_),
    .A2(_08536_),
    .B1(_08538_),
    .Y(_08539_));
 sky130_fd_sc_hd__a21oi_2 _30168_ (.A1(_08533_),
    .A2(_08534_),
    .B1(_08531_),
    .Y(_08540_));
 sky130_fd_sc_hd__nor3b_2 _30169_ (.A(_08537_),
    .B(_08540_),
    .C_N(_08536_),
    .Y(_08541_));
 sky130_fd_sc_hd__a21oi_2 _30170_ (.A1(_08278_),
    .A2(_08273_),
    .B1(_08275_),
    .Y(_08542_));
 sky130_fd_sc_hd__o21ai_2 _30171_ (.A1(_08280_),
    .A2(_08542_),
    .B1(_08279_),
    .Y(_08543_));
 sky130_fd_sc_hd__o21bai_2 _30172_ (.A1(_08539_),
    .A2(_08541_),
    .B1_N(_08543_),
    .Y(_08544_));
 sky130_fd_sc_hd__nand2_2 _30173_ (.A(_08532_),
    .B(_08536_),
    .Y(_08545_));
 sky130_fd_sc_hd__nand2_2 _30174_ (.A(_08545_),
    .B(_08537_),
    .Y(_08546_));
 sky130_fd_sc_hd__nand3_2 _30175_ (.A(_08532_),
    .B(_08538_),
    .C(_08536_),
    .Y(_08547_));
 sky130_fd_sc_hd__nand3_2 _30176_ (.A(_08546_),
    .B(_08543_),
    .C(_08547_),
    .Y(_08548_));
 sky130_fd_sc_hd__buf_1 _30177_ (.A(_07960_),
    .X(_08549_));
 sky130_fd_sc_hd__a22o_2 _30178_ (.A1(_05926_),
    .A2(_07966_),
    .B1(_05929_),
    .B2(_08549_),
    .X(_08550_));
 sky130_fd_sc_hd__buf_1 _30179_ (.A(_19202_),
    .X(_08551_));
 sky130_fd_sc_hd__nand2_2 _30180_ (.A(_06040_),
    .B(_08551_),
    .Y(_08552_));
 sky130_fd_sc_hd__buf_1 _30181_ (.A(_07745_),
    .X(_08553_));
 sky130_fd_sc_hd__nand3b_2 _30182_ (.A_N(_08552_),
    .B(_05638_),
    .C(_08553_),
    .Y(_08554_));
 sky130_fd_sc_hd__o2bb2ai_2 _30183_ (.A1_N(_08550_),
    .A2_N(_08554_),
    .B1(_18880_),
    .B2(_19174_),
    .Y(_08555_));
 sky130_fd_sc_hd__buf_1 _30184_ (.A(\pcpi_mul.rs1[24] ),
    .X(_08556_));
 sky130_fd_sc_hd__buf_1 _30185_ (.A(_08556_),
    .X(_08557_));
 sky130_fd_sc_hd__and2_2 _30186_ (.A(_06732_),
    .B(_08557_),
    .X(_08558_));
 sky130_fd_sc_hd__nand3_2 _30187_ (.A(_08554_),
    .B(_08550_),
    .C(_08558_),
    .Y(_08559_));
 sky130_fd_sc_hd__a21oi_2 _30188_ (.A1(_08297_),
    .A2(_08296_),
    .B1(_08294_),
    .Y(_08560_));
 sky130_vsdinv _30189_ (.A(_08560_),
    .Y(_08561_));
 sky130_fd_sc_hd__a21o_2 _30190_ (.A1(_08555_),
    .A2(_08559_),
    .B1(_08561_),
    .X(_08562_));
 sky130_fd_sc_hd__nand3_2 _30191_ (.A(_08555_),
    .B(_08561_),
    .C(_08559_),
    .Y(_08563_));
 sky130_fd_sc_hd__buf_1 _30192_ (.A(_08563_),
    .X(_08564_));
 sky130_fd_sc_hd__buf_1 _30193_ (.A(_19184_),
    .X(_08565_));
 sky130_fd_sc_hd__nand2_2 _30194_ (.A(_05549_),
    .B(_08565_),
    .Y(_08566_));
 sky130_fd_sc_hd__nand2_2 _30195_ (.A(_07323_),
    .B(_19180_),
    .Y(_08567_));
 sky130_fd_sc_hd__xor2_2 _30196_ (.A(_08566_),
    .B(_08567_),
    .X(_08568_));
 sky130_fd_sc_hd__buf_1 _30197_ (.A(\pcpi_mul.rs1[21] ),
    .X(_08569_));
 sky130_fd_sc_hd__buf_1 _30198_ (.A(_08569_),
    .X(_08570_));
 sky130_fd_sc_hd__buf_1 _30199_ (.A(_08570_),
    .X(_08571_));
 sky130_fd_sc_hd__and2_2 _30200_ (.A(_05459_),
    .B(_08571_),
    .X(_08572_));
 sky130_fd_sc_hd__nand2_2 _30201_ (.A(_08568_),
    .B(_08572_),
    .Y(_08573_));
 sky130_fd_sc_hd__xnor2_2 _30202_ (.A(_08566_),
    .B(_08567_),
    .Y(_08574_));
 sky130_fd_sc_hd__o21ai_2 _30203_ (.A1(_07332_),
    .A2(_19193_),
    .B1(_08574_),
    .Y(_08575_));
 sky130_fd_sc_hd__nand2_2 _30204_ (.A(_08573_),
    .B(_08575_),
    .Y(_08576_));
 sky130_fd_sc_hd__buf_1 _30205_ (.A(_08576_),
    .X(_08577_));
 sky130_fd_sc_hd__a21boi_2 _30206_ (.A1(_08562_),
    .A2(_08564_),
    .B1_N(_08577_),
    .Y(_08578_));
 sky130_fd_sc_hd__a21oi_2 _30207_ (.A1(_08555_),
    .A2(_08559_),
    .B1(_08561_),
    .Y(_08579_));
 sky130_fd_sc_hd__nor3b_2 _30208_ (.A(_08577_),
    .B(_08579_),
    .C_N(_08563_),
    .Y(_08580_));
 sky130_fd_sc_hd__a21oi_2 _30209_ (.A1(_08306_),
    .A2(_08298_),
    .B1(_08307_),
    .Y(_08581_));
 sky130_fd_sc_hd__o21ai_2 _30210_ (.A1(_08319_),
    .A2(_08581_),
    .B1(_08309_),
    .Y(_08582_));
 sky130_fd_sc_hd__o21bai_2 _30211_ (.A1(_08578_),
    .A2(_08580_),
    .B1_N(_08582_),
    .Y(_08583_));
 sky130_fd_sc_hd__nand2_2 _30212_ (.A(_08562_),
    .B(_08564_),
    .Y(_08584_));
 sky130_fd_sc_hd__nand2_2 _30213_ (.A(_08584_),
    .B(_08577_),
    .Y(_08585_));
 sky130_fd_sc_hd__nand3b_2 _30214_ (.A_N(_08577_),
    .B(_08562_),
    .C(_08564_),
    .Y(_08586_));
 sky130_fd_sc_hd__nand3_2 _30215_ (.A(_08585_),
    .B(_08586_),
    .C(_08582_),
    .Y(_08587_));
 sky130_fd_sc_hd__o21a_2 _30216_ (.A1(_08311_),
    .A2(_08312_),
    .B1(_08316_),
    .X(_08588_));
 sky130_vsdinv _30217_ (.A(_08588_),
    .Y(_08589_));
 sky130_fd_sc_hd__a21oi_2 _30218_ (.A1(_08583_),
    .A2(_08587_),
    .B1(_08589_),
    .Y(_08590_));
 sky130_fd_sc_hd__nand3_2 _30219_ (.A(_08583_),
    .B(_08589_),
    .C(_08587_),
    .Y(_08591_));
 sky130_vsdinv _30220_ (.A(_08591_),
    .Y(_08592_));
 sky130_fd_sc_hd__nor2_2 _30221_ (.A(_08590_),
    .B(_08592_),
    .Y(_08593_));
 sky130_fd_sc_hd__a21oi_2 _30222_ (.A1(_08544_),
    .A2(_08548_),
    .B1(_08593_),
    .Y(_08594_));
 sky130_fd_sc_hd__nand2_2 _30223_ (.A(_08583_),
    .B(_08587_),
    .Y(_08595_));
 sky130_fd_sc_hd__nand2_2 _30224_ (.A(_08595_),
    .B(_08588_),
    .Y(_08596_));
 sky130_fd_sc_hd__nand2_2 _30225_ (.A(_08596_),
    .B(_08591_),
    .Y(_08597_));
 sky130_fd_sc_hd__a21oi_2 _30226_ (.A1(_08546_),
    .A2(_08547_),
    .B1(_08543_),
    .Y(_08598_));
 sky130_vsdinv _30227_ (.A(_08548_),
    .Y(_08599_));
 sky130_fd_sc_hd__nor3_2 _30228_ (.A(_08597_),
    .B(_08598_),
    .C(_08599_),
    .Y(_08600_));
 sky130_fd_sc_hd__o21ai_2 _30229_ (.A1(_08204_),
    .A2(_08198_),
    .B1(_08208_),
    .Y(_08601_));
 sky130_fd_sc_hd__o21bai_2 _30230_ (.A1(_08594_),
    .A2(_08600_),
    .B1_N(_08601_),
    .Y(_08602_));
 sky130_fd_sc_hd__o2bb2ai_2 _30231_ (.A1_N(_08548_),
    .A2_N(_08544_),
    .B1(_08592_),
    .B2(_08590_),
    .Y(_08603_));
 sky130_fd_sc_hd__nand3_2 _30232_ (.A(_08593_),
    .B(_08544_),
    .C(_08548_),
    .Y(_08604_));
 sky130_fd_sc_hd__nand3_2 _30233_ (.A(_08603_),
    .B(_08604_),
    .C(_08601_),
    .Y(_08605_));
 sky130_fd_sc_hd__nand3b_2 _30234_ (.A_N(_08509_),
    .B(_08602_),
    .C(_08605_),
    .Y(_08606_));
 sky130_fd_sc_hd__buf_1 _30235_ (.A(_08606_),
    .X(_08607_));
 sky130_fd_sc_hd__nand2_2 _30236_ (.A(_08602_),
    .B(_08605_),
    .Y(_08608_));
 sky130_fd_sc_hd__nand2_2 _30237_ (.A(_08608_),
    .B(_08509_),
    .Y(_08609_));
 sky130_fd_sc_hd__buf_1 _30238_ (.A(_08609_),
    .X(_08610_));
 sky130_fd_sc_hd__a22oi_2 _30239_ (.A1(_08503_),
    .A2(_08507_),
    .B1(_08607_),
    .B2(_08610_),
    .Y(_08611_));
 sky130_fd_sc_hd__nand2_2 _30240_ (.A(_08503_),
    .B(_08507_),
    .Y(_08612_));
 sky130_fd_sc_hd__nand2_2 _30241_ (.A(_08610_),
    .B(_08606_),
    .Y(_08613_));
 sky130_fd_sc_hd__nor2_2 _30242_ (.A(_08612_),
    .B(_08613_),
    .Y(_08614_));
 sky130_fd_sc_hd__a31oi_2 _30243_ (.A1(_08348_),
    .A2(_08354_),
    .A3(_08344_),
    .B1(_08251_),
    .Y(_08615_));
 sky130_fd_sc_hd__o21ai_2 _30244_ (.A1(_08611_),
    .A2(_08614_),
    .B1(_08615_),
    .Y(_08616_));
 sky130_fd_sc_hd__a31o_2 _30245_ (.A1(_08348_),
    .A2(_08354_),
    .A3(_08343_),
    .B1(_08251_),
    .X(_08617_));
 sky130_fd_sc_hd__a21oi_2 _30246_ (.A1(_08505_),
    .A2(_08506_),
    .B1(_08353_),
    .Y(_08618_));
 sky130_fd_sc_hd__nor3_2 _30247_ (.A(_08248_),
    .B(_08499_),
    .C(_08502_),
    .Y(_08619_));
 sky130_fd_sc_hd__nor2_2 _30248_ (.A(_08618_),
    .B(_08619_),
    .Y(_08620_));
 sky130_fd_sc_hd__nand3_2 _30249_ (.A(_08620_),
    .B(_08607_),
    .C(_08610_),
    .Y(_08621_));
 sky130_fd_sc_hd__nand2_2 _30250_ (.A(_08613_),
    .B(_08612_),
    .Y(_08622_));
 sky130_fd_sc_hd__nand3_2 _30251_ (.A(_08617_),
    .B(_08621_),
    .C(_08622_),
    .Y(_08623_));
 sky130_fd_sc_hd__nand2_2 _30252_ (.A(_08616_),
    .B(_08623_),
    .Y(_08624_));
 sky130_fd_sc_hd__a21boi_2 _30253_ (.A1(_08324_),
    .A2(_08327_),
    .B1_N(_08325_),
    .Y(_08625_));
 sky130_fd_sc_hd__o21ai_2 _30254_ (.A1(_08338_),
    .A2(_08345_),
    .B1(_08342_),
    .Y(_08626_));
 sky130_fd_sc_hd__xnor2_2 _30255_ (.A(_08625_),
    .B(_08626_),
    .Y(_08627_));
 sky130_vsdinv _30256_ (.A(_08627_),
    .Y(_08628_));
 sky130_fd_sc_hd__nand2_2 _30257_ (.A(_08624_),
    .B(_08628_),
    .Y(_08629_));
 sky130_fd_sc_hd__nand3_2 _30258_ (.A(_08616_),
    .B(_08623_),
    .C(_08627_),
    .Y(_08630_));
 sky130_fd_sc_hd__nand2_2 _30259_ (.A(_08629_),
    .B(_08630_),
    .Y(_08631_));
 sky130_fd_sc_hd__a21boi_2 _30260_ (.A1(_08363_),
    .A2(_08369_),
    .B1_N(_08360_),
    .Y(_08632_));
 sky130_fd_sc_hd__nand2_2 _30261_ (.A(_08631_),
    .B(_08632_),
    .Y(_08633_));
 sky130_fd_sc_hd__nand2_2 _30262_ (.A(_08370_),
    .B(_08360_),
    .Y(_08634_));
 sky130_fd_sc_hd__nand3_2 _30263_ (.A(_08634_),
    .B(_08630_),
    .C(_08629_),
    .Y(_08635_));
 sky130_fd_sc_hd__buf_1 _30264_ (.A(_08365_),
    .X(_08636_));
 sky130_fd_sc_hd__a21oi_2 _30265_ (.A1(_08633_),
    .A2(_08635_),
    .B1(_08636_),
    .Y(_08637_));
 sky130_vsdinv _30266_ (.A(_08636_),
    .Y(_08638_));
 sky130_fd_sc_hd__a21oi_2 _30267_ (.A1(_08629_),
    .A2(_08630_),
    .B1(_08634_),
    .Y(_08639_));
 sky130_fd_sc_hd__nor2_2 _30268_ (.A(_08632_),
    .B(_08631_),
    .Y(_08640_));
 sky130_fd_sc_hd__nor3_2 _30269_ (.A(_08638_),
    .B(_08639_),
    .C(_08640_),
    .Y(_08641_));
 sky130_vsdinv _30270_ (.A(_08376_),
    .Y(_08642_));
 sky130_fd_sc_hd__a21oi_2 _30271_ (.A1(_08367_),
    .A2(_08370_),
    .B1(_08135_),
    .Y(_08643_));
 sky130_fd_sc_hd__o21ai_2 _30272_ (.A1(_08642_),
    .A2(_08643_),
    .B1(_08371_),
    .Y(_08644_));
 sky130_fd_sc_hd__o21bai_2 _30273_ (.A1(_08637_),
    .A2(_08641_),
    .B1_N(_08644_),
    .Y(_08645_));
 sky130_fd_sc_hd__o21bai_2 _30274_ (.A1(_08639_),
    .A2(_08640_),
    .B1_N(_08636_),
    .Y(_08646_));
 sky130_fd_sc_hd__nand3_2 _30275_ (.A(_08633_),
    .B(_08636_),
    .C(_08635_),
    .Y(_08647_));
 sky130_fd_sc_hd__nand3_2 _30276_ (.A(_08646_),
    .B(_08647_),
    .C(_08644_),
    .Y(_08648_));
 sky130_fd_sc_hd__nand2_2 _30277_ (.A(_08645_),
    .B(_08648_),
    .Y(_08649_));
 sky130_fd_sc_hd__nand3_2 _30278_ (.A(_08131_),
    .B(_08130_),
    .C(_08383_),
    .Y(_08650_));
 sky130_fd_sc_hd__nor2_2 _30279_ (.A(_08650_),
    .B(_07682_),
    .Y(_08651_));
 sky130_fd_sc_hd__nand3_2 _30280_ (.A(_08123_),
    .B(_08124_),
    .C(_08125_),
    .Y(_08652_));
 sky130_fd_sc_hd__nand3_2 _30281_ (.A(_08375_),
    .B(_08378_),
    .C(_08377_),
    .Y(_08653_));
 sky130_fd_sc_hd__o21ai_2 _30282_ (.A1(_08652_),
    .A2(_08379_),
    .B1(_08653_),
    .Y(_08654_));
 sky130_fd_sc_hd__a31oi_2 _30283_ (.A1(_08383_),
    .A2(_08130_),
    .A3(_08133_),
    .B1(_08654_),
    .Y(_08655_));
 sky130_fd_sc_hd__o21ai_2 _30284_ (.A1(_08650_),
    .A2(_07686_),
    .B1(_08655_),
    .Y(_08656_));
 sky130_fd_sc_hd__a21oi_2 _30285_ (.A1(_06877_),
    .A2(_08651_),
    .B1(_08656_),
    .Y(_08657_));
 sky130_fd_sc_hd__xor2_2 _30286_ (.A(_08649_),
    .B(_08657_),
    .X(_02643_));
 sky130_fd_sc_hd__a22oi_2 _30287_ (.A1(_07785_),
    .A2(_05840_),
    .B1(_18784_),
    .B2(_05949_),
    .Y(_08658_));
 sky130_fd_sc_hd__nand2_2 _30288_ (.A(_07164_),
    .B(_05727_),
    .Y(_08659_));
 sky130_fd_sc_hd__nand2_2 _30289_ (.A(_07168_),
    .B(_06342_),
    .Y(_08660_));
 sky130_fd_sc_hd__nor2_2 _30290_ (.A(_08659_),
    .B(_08660_),
    .Y(_08661_));
 sky130_fd_sc_hd__and2_2 _30291_ (.A(_18789_),
    .B(_06062_),
    .X(_08662_));
 sky130_fd_sc_hd__o21bai_2 _30292_ (.A1(_08658_),
    .A2(_08661_),
    .B1_N(_08662_),
    .Y(_08663_));
 sky130_fd_sc_hd__nand3b_2 _30293_ (.A_N(_08659_),
    .B(_08012_),
    .C(_06060_),
    .Y(_08664_));
 sky130_fd_sc_hd__nand3b_2 _30294_ (.A_N(_08658_),
    .B(_08664_),
    .C(_08662_),
    .Y(_08665_));
 sky130_fd_sc_hd__nand2_2 _30295_ (.A(_08663_),
    .B(_08665_),
    .Y(_08666_));
 sky130_fd_sc_hd__a21oi_2 _30296_ (.A1(_08485_),
    .A2(_08488_),
    .B1(_08484_),
    .Y(_08667_));
 sky130_fd_sc_hd__nand2_2 _30297_ (.A(_08666_),
    .B(_08667_),
    .Y(_08668_));
 sky130_fd_sc_hd__nand3b_2 _30298_ (.A_N(_08667_),
    .B(_08665_),
    .C(_08663_),
    .Y(_08669_));
 sky130_fd_sc_hd__buf_1 _30299_ (.A(_08669_),
    .X(_08670_));
 sky130_fd_sc_hd__nand2_2 _30300_ (.A(_08668_),
    .B(_08670_),
    .Y(_08671_));
 sky130_fd_sc_hd__a21oi_2 _30301_ (.A1(_08393_),
    .A2(_08389_),
    .B1(_08388_),
    .Y(_08672_));
 sky130_fd_sc_hd__nand2_2 _30302_ (.A(_08671_),
    .B(_08672_),
    .Y(_08673_));
 sky130_vsdinv _30303_ (.A(_08672_),
    .Y(_08674_));
 sky130_fd_sc_hd__nand3_2 _30304_ (.A(_08668_),
    .B(_08674_),
    .C(_08669_),
    .Y(_08675_));
 sky130_fd_sc_hd__o21ai_2 _30305_ (.A1(_08401_),
    .A2(_08404_),
    .B1(_08400_),
    .Y(_08676_));
 sky130_fd_sc_hd__a21oi_2 _30306_ (.A1(_08673_),
    .A2(_08675_),
    .B1(_08676_),
    .Y(_08677_));
 sky130_fd_sc_hd__a21oi_2 _30307_ (.A1(_08399_),
    .A2(_08402_),
    .B1(_08405_),
    .Y(_08678_));
 sky130_fd_sc_hd__a21oi_2 _30308_ (.A1(_08668_),
    .A2(_08670_),
    .B1(_08674_),
    .Y(_08679_));
 sky130_vsdinv _30309_ (.A(_08675_),
    .Y(_08680_));
 sky130_fd_sc_hd__nor3_2 _30310_ (.A(_08678_),
    .B(_08679_),
    .C(_08680_),
    .Y(_08681_));
 sky130_fd_sc_hd__nand2_2 _30311_ (.A(_07190_),
    .B(_07515_),
    .Y(_08682_));
 sky130_fd_sc_hd__nand2_2 _30312_ (.A(_07200_),
    .B(_06477_),
    .Y(_08683_));
 sky130_fd_sc_hd__nor2_2 _30313_ (.A(_08682_),
    .B(_08683_),
    .Y(_08684_));
 sky130_fd_sc_hd__and2_2 _30314_ (.A(_06274_),
    .B(_08181_),
    .X(_08685_));
 sky130_fd_sc_hd__nand2_2 _30315_ (.A(_08682_),
    .B(_08683_),
    .Y(_08686_));
 sky130_fd_sc_hd__nand3b_2 _30316_ (.A_N(_08684_),
    .B(_08685_),
    .C(_08686_),
    .Y(_08687_));
 sky130_fd_sc_hd__buf_1 _30317_ (.A(_06392_),
    .X(_08688_));
 sky130_fd_sc_hd__a22oi_2 _30318_ (.A1(_18798_),
    .A2(_06203_),
    .B1(_08688_),
    .B2(_06478_),
    .Y(_08689_));
 sky130_fd_sc_hd__o21bai_2 _30319_ (.A1(_08689_),
    .A2(_08684_),
    .B1_N(_08685_),
    .Y(_08690_));
 sky130_fd_sc_hd__a21oi_2 _30320_ (.A1(_08419_),
    .A2(_08418_),
    .B1(_08417_),
    .Y(_08691_));
 sky130_fd_sc_hd__a21bo_2 _30321_ (.A1(_08687_),
    .A2(_08690_),
    .B1_N(_08691_),
    .X(_08692_));
 sky130_fd_sc_hd__nand3b_2 _30322_ (.A_N(_08691_),
    .B(_08687_),
    .C(_08690_),
    .Y(_08693_));
 sky130_fd_sc_hd__nand2_2 _30323_ (.A(_08692_),
    .B(_08693_),
    .Y(_08694_));
 sky130_fd_sc_hd__nand2_2 _30324_ (.A(_08178_),
    .B(_19231_),
    .Y(_08695_));
 sky130_fd_sc_hd__nand2_2 _30325_ (.A(_08180_),
    .B(_06744_),
    .Y(_08696_));
 sky130_fd_sc_hd__nand2_2 _30326_ (.A(_08695_),
    .B(_08696_),
    .Y(_08697_));
 sky130_fd_sc_hd__nor2_2 _30327_ (.A(_08695_),
    .B(_08696_),
    .Y(_08698_));
 sky130_vsdinv _30328_ (.A(_08698_),
    .Y(_08699_));
 sky130_fd_sc_hd__o2bb2ai_2 _30329_ (.A1_N(_08697_),
    .A2_N(_08699_),
    .B1(_07214_),
    .B2(_19217_),
    .Y(_08700_));
 sky130_fd_sc_hd__and2_2 _30330_ (.A(_18822_),
    .B(_06734_),
    .X(_08701_));
 sky130_fd_sc_hd__nand3b_2 _30331_ (.A_N(_08698_),
    .B(_08701_),
    .C(_08697_),
    .Y(_08702_));
 sky130_fd_sc_hd__nand2_2 _30332_ (.A(_08700_),
    .B(_08702_),
    .Y(_08703_));
 sky130_fd_sc_hd__nand2_2 _30333_ (.A(_08694_),
    .B(_08703_),
    .Y(_08704_));
 sky130_fd_sc_hd__nand3b_2 _30334_ (.A_N(_08703_),
    .B(_08693_),
    .C(_08692_),
    .Y(_08705_));
 sky130_fd_sc_hd__nand2_2 _30335_ (.A(_08704_),
    .B(_08705_),
    .Y(_08706_));
 sky130_fd_sc_hd__o21ai_2 _30336_ (.A1(_08677_),
    .A2(_08681_),
    .B1(_08706_),
    .Y(_08707_));
 sky130_fd_sc_hd__o21bai_2 _30337_ (.A1(_08679_),
    .A2(_08680_),
    .B1_N(_08676_),
    .Y(_08708_));
 sky130_fd_sc_hd__nand3_2 _30338_ (.A(_08673_),
    .B(_08675_),
    .C(_08676_),
    .Y(_08709_));
 sky130_fd_sc_hd__nand3b_2 _30339_ (.A_N(_08706_),
    .B(_08708_),
    .C(_08709_),
    .Y(_08710_));
 sky130_vsdinv _30340_ (.A(_08495_),
    .Y(_08711_));
 sky130_fd_sc_hd__a21oi_2 _30341_ (.A1(_08707_),
    .A2(_08710_),
    .B1(_08711_),
    .Y(_08712_));
 sky130_fd_sc_hd__nand3_2 _30342_ (.A(_08707_),
    .B(_08711_),
    .C(_08710_),
    .Y(_08713_));
 sky130_vsdinv _30343_ (.A(_08713_),
    .Y(_08714_));
 sky130_fd_sc_hd__o21a_2 _30344_ (.A1(_08440_),
    .A2(_08447_),
    .B1(_08442_),
    .X(_08715_));
 sky130_vsdinv _30345_ (.A(_08715_),
    .Y(_08716_));
 sky130_fd_sc_hd__o21bai_2 _30346_ (.A1(_08712_),
    .A2(_08714_),
    .B1_N(_08716_),
    .Y(_08717_));
 sky130_fd_sc_hd__nand2_2 _30347_ (.A(_08707_),
    .B(_08710_),
    .Y(_08718_));
 sky130_fd_sc_hd__nand2_2 _30348_ (.A(_08718_),
    .B(_08495_),
    .Y(_08719_));
 sky130_fd_sc_hd__nand3_2 _30349_ (.A(_08719_),
    .B(_08716_),
    .C(_08713_),
    .Y(_08720_));
 sky130_fd_sc_hd__buf_1 _30350_ (.A(_08720_),
    .X(_08721_));
 sky130_fd_sc_hd__nand2_2 _30351_ (.A(_08463_),
    .B(_05635_),
    .Y(_08722_));
 sky130_fd_sc_hd__nand2_2 _30352_ (.A(_08465_),
    .B(_06826_),
    .Y(_08723_));
 sky130_fd_sc_hd__nor2_2 _30353_ (.A(_08722_),
    .B(_08723_),
    .Y(_08724_));
 sky130_fd_sc_hd__buf_1 _30354_ (.A(_05468_),
    .X(_08725_));
 sky130_fd_sc_hd__and2_2 _30355_ (.A(_18758_),
    .B(_08725_),
    .X(_08726_));
 sky130_fd_sc_hd__nand2_2 _30356_ (.A(_08722_),
    .B(_08723_),
    .Y(_08727_));
 sky130_fd_sc_hd__nand3b_2 _30357_ (.A_N(_08724_),
    .B(_08726_),
    .C(_08727_),
    .Y(_08728_));
 sky130_fd_sc_hd__buf_1 _30358_ (.A(_08462_),
    .X(_08729_));
 sky130_fd_sc_hd__buf_1 _30359_ (.A(_08729_),
    .X(_08730_));
 sky130_fd_sc_hd__buf_1 _30360_ (.A(_08465_),
    .X(_08731_));
 sky130_fd_sc_hd__a22oi_2 _30361_ (.A1(_08730_),
    .A2(_05636_),
    .B1(_08731_),
    .B2(_05639_),
    .Y(_08732_));
 sky130_fd_sc_hd__o21bai_2 _30362_ (.A1(_08732_),
    .A2(_08724_),
    .B1_N(_08726_),
    .Y(_08733_));
 sky130_fd_sc_hd__nand2_2 _30363_ (.A(_08728_),
    .B(_08733_),
    .Y(_08734_));
 sky130_fd_sc_hd__a21oi_2 _30364_ (.A1(_08469_),
    .A2(_08468_),
    .B1(_08467_),
    .Y(_08735_));
 sky130_fd_sc_hd__nand2_2 _30365_ (.A(_08734_),
    .B(_08735_),
    .Y(_08736_));
 sky130_fd_sc_hd__nand3b_2 _30366_ (.A_N(_08735_),
    .B(_08728_),
    .C(_08733_),
    .Y(_08737_));
 sky130_fd_sc_hd__nand2_2 _30367_ (.A(_08736_),
    .B(_08737_),
    .Y(_08738_));
 sky130_fd_sc_hd__nand2_2 _30368_ (.A(_08217_),
    .B(_19277_),
    .Y(_08739_));
 sky130_fd_sc_hd__nand2_2 _30369_ (.A(_08214_),
    .B(_08480_),
    .Y(_08740_));
 sky130_fd_sc_hd__nand2_2 _30370_ (.A(_08739_),
    .B(_08740_),
    .Y(_08741_));
 sky130_fd_sc_hd__nor2_2 _30371_ (.A(_08739_),
    .B(_08740_),
    .Y(_08742_));
 sky130_vsdinv _30372_ (.A(_08742_),
    .Y(_08743_));
 sky130_fd_sc_hd__o2bb2ai_2 _30373_ (.A1_N(_08741_),
    .A2_N(_08743_),
    .B1(_18776_),
    .B2(_19269_),
    .Y(_08744_));
 sky130_fd_sc_hd__and2_2 _30374_ (.A(_07532_),
    .B(_07208_),
    .X(_08745_));
 sky130_fd_sc_hd__nand3b_2 _30375_ (.A_N(_08742_),
    .B(_08745_),
    .C(_08741_),
    .Y(_08746_));
 sky130_fd_sc_hd__nand2_2 _30376_ (.A(_08744_),
    .B(_08746_),
    .Y(_08747_));
 sky130_fd_sc_hd__nand2_2 _30377_ (.A(_08738_),
    .B(_08747_),
    .Y(_08748_));
 sky130_fd_sc_hd__nand3b_2 _30378_ (.A_N(_08747_),
    .B(_08737_),
    .C(_08736_),
    .Y(_08749_));
 sky130_fd_sc_hd__nand2_2 _30379_ (.A(_08492_),
    .B(_08477_),
    .Y(_08750_));
 sky130_fd_sc_hd__a21oi_2 _30380_ (.A1(_08748_),
    .A2(_08749_),
    .B1(_08750_),
    .Y(_08751_));
 sky130_fd_sc_hd__nand3_2 _30381_ (.A(_08750_),
    .B(_08749_),
    .C(_08748_),
    .Y(_08752_));
 sky130_vsdinv _30382_ (.A(_08752_),
    .Y(_08753_));
 sky130_fd_sc_hd__buf_1 _30383_ (.A(\pcpi_mul.rs2[25] ),
    .X(_08754_));
 sky130_fd_sc_hd__buf_1 _30384_ (.A(_08754_),
    .X(_08755_));
 sky130_fd_sc_hd__buf_1 _30385_ (.A(_08755_),
    .X(_08756_));
 sky130_fd_sc_hd__nand2_2 _30386_ (.A(_08756_),
    .B(_05239_),
    .Y(_08757_));
 sky130_fd_sc_hd__buf_1 _30387_ (.A(\pcpi_mul.rs2[24] ),
    .X(_08758_));
 sky130_fd_sc_hd__buf_1 _30388_ (.A(_08758_),
    .X(_08759_));
 sky130_fd_sc_hd__nand2_2 _30389_ (.A(_08759_),
    .B(_05425_),
    .Y(_08760_));
 sky130_fd_sc_hd__xor2_2 _30390_ (.A(_08757_),
    .B(_08760_),
    .X(_08761_));
 sky130_fd_sc_hd__o21bai_2 _30391_ (.A1(_08751_),
    .A2(_08753_),
    .B1_N(_08761_),
    .Y(_08762_));
 sky130_fd_sc_hd__a21o_2 _30392_ (.A1(_08748_),
    .A2(_08749_),
    .B1(_08750_),
    .X(_08763_));
 sky130_fd_sc_hd__nand3_2 _30393_ (.A(_08763_),
    .B(_08761_),
    .C(_08752_),
    .Y(_08764_));
 sky130_fd_sc_hd__buf_1 _30394_ (.A(_08764_),
    .X(_08765_));
 sky130_fd_sc_hd__nand3_2 _30395_ (.A(_08494_),
    .B(_08461_),
    .C(_08495_),
    .Y(_08766_));
 sky130_fd_sc_hd__a21boi_2 _30396_ (.A1(_08762_),
    .A2(_08765_),
    .B1_N(_08766_),
    .Y(_08767_));
 sky130_fd_sc_hd__a21oi_2 _30397_ (.A1(_08763_),
    .A2(_08752_),
    .B1(_08761_),
    .Y(_08768_));
 sky130_vsdinv _30398_ (.A(_08764_),
    .Y(_08769_));
 sky130_fd_sc_hd__nor3_2 _30399_ (.A(_08766_),
    .B(_08768_),
    .C(_08769_),
    .Y(_08770_));
 sky130_fd_sc_hd__nor2_2 _30400_ (.A(_08767_),
    .B(_08770_),
    .Y(_08771_));
 sky130_fd_sc_hd__a21oi_2 _30401_ (.A1(_08717_),
    .A2(_08721_),
    .B1(_08771_),
    .Y(_08772_));
 sky130_fd_sc_hd__o21ai_2 _30402_ (.A1(_08768_),
    .A2(_08769_),
    .B1(_08766_),
    .Y(_08773_));
 sky130_fd_sc_hd__nand3b_2 _30403_ (.A_N(_08766_),
    .B(_08762_),
    .C(_08765_),
    .Y(_08774_));
 sky130_fd_sc_hd__nand2_2 _30404_ (.A(_08773_),
    .B(_08774_),
    .Y(_08775_));
 sky130_fd_sc_hd__a21oi_2 _30405_ (.A1(_08719_),
    .A2(_08713_),
    .B1(_08716_),
    .Y(_08776_));
 sky130_fd_sc_hd__nor3b_2 _30406_ (.A(_08775_),
    .B(_08776_),
    .C_N(_08720_),
    .Y(_08777_));
 sky130_fd_sc_hd__o22ai_2 _30407_ (.A1(_08497_),
    .A2(_08504_),
    .B1(_08772_),
    .B2(_08777_),
    .Y(_08778_));
 sky130_fd_sc_hd__buf_1 _30408_ (.A(_08778_),
    .X(_08779_));
 sky130_fd_sc_hd__o2bb2ai_2 _30409_ (.A1_N(_08721_),
    .A2_N(_08717_),
    .B1(_08770_),
    .B2(_08767_),
    .Y(_08780_));
 sky130_fd_sc_hd__nand3_2 _30410_ (.A(_08717_),
    .B(_08771_),
    .C(_08721_),
    .Y(_08781_));
 sky130_fd_sc_hd__nand3_2 _30411_ (.A(_08780_),
    .B(_08502_),
    .C(_08781_),
    .Y(_08782_));
 sky130_fd_sc_hd__a22oi_2 _30412_ (.A1(_06881_),
    .A2(_06936_),
    .B1(_07271_),
    .B2(_08299_),
    .Y(_08783_));
 sky130_fd_sc_hd__and4_2 _30413_ (.A(_07548_),
    .B(_07271_),
    .C(_07325_),
    .D(_07321_),
    .X(_08784_));
 sky130_fd_sc_hd__and2_2 _30414_ (.A(_05586_),
    .B(_08302_),
    .X(_08785_));
 sky130_fd_sc_hd__o21bai_2 _30415_ (.A1(_08783_),
    .A2(_08784_),
    .B1_N(_08785_),
    .Y(_08786_));
 sky130_fd_sc_hd__nand2_2 _30416_ (.A(_18828_),
    .B(_07946_),
    .Y(_08787_));
 sky130_fd_sc_hd__nand3b_2 _30417_ (.A_N(_08787_),
    .B(_18833_),
    .C(_07106_),
    .Y(_08788_));
 sky130_fd_sc_hd__nand3b_2 _30418_ (.A_N(_08783_),
    .B(_08788_),
    .C(_08785_),
    .Y(_08789_));
 sky130_fd_sc_hd__nand2_2 _30419_ (.A(_08786_),
    .B(_08789_),
    .Y(_08790_));
 sky130_fd_sc_hd__a21oi_2 _30420_ (.A1(_08429_),
    .A2(_08433_),
    .B1(_08430_),
    .Y(_08791_));
 sky130_fd_sc_hd__nand2_2 _30421_ (.A(_08790_),
    .B(_08791_),
    .Y(_08792_));
 sky130_fd_sc_hd__nand3b_2 _30422_ (.A_N(_08791_),
    .B(_08786_),
    .C(_08789_),
    .Y(_08793_));
 sky130_fd_sc_hd__a21oi_2 _30423_ (.A1(_08518_),
    .A2(_08515_),
    .B1(_08514_),
    .Y(_08794_));
 sky130_vsdinv _30424_ (.A(_08794_),
    .Y(_08795_));
 sky130_fd_sc_hd__a21oi_2 _30425_ (.A1(_08792_),
    .A2(_08793_),
    .B1(_08795_),
    .Y(_08796_));
 sky130_fd_sc_hd__nand3_2 _30426_ (.A(_08792_),
    .B(_08795_),
    .C(_08793_),
    .Y(_08797_));
 sky130_vsdinv _30427_ (.A(_08797_),
    .Y(_08798_));
 sky130_fd_sc_hd__o21ai_2 _30428_ (.A1(_08435_),
    .A2(_08424_),
    .B1(_08425_),
    .Y(_08799_));
 sky130_fd_sc_hd__o21bai_2 _30429_ (.A1(_08796_),
    .A2(_08798_),
    .B1_N(_08799_),
    .Y(_08800_));
 sky130_fd_sc_hd__a21o_2 _30430_ (.A1(_08792_),
    .A2(_08793_),
    .B1(_08795_),
    .X(_08801_));
 sky130_fd_sc_hd__nand3_2 _30431_ (.A(_08801_),
    .B(_08799_),
    .C(_08797_),
    .Y(_08802_));
 sky130_fd_sc_hd__nand2_2 _30432_ (.A(_08800_),
    .B(_08802_),
    .Y(_08803_));
 sky130_fd_sc_hd__a21boi_2 _30433_ (.A1(_08522_),
    .A2(_08526_),
    .B1_N(_08523_),
    .Y(_08804_));
 sky130_fd_sc_hd__nand2_2 _30434_ (.A(_08803_),
    .B(_08804_),
    .Y(_08805_));
 sky130_fd_sc_hd__nand3b_2 _30435_ (.A_N(_08804_),
    .B(_08800_),
    .C(_08802_),
    .Y(_08806_));
 sky130_fd_sc_hd__nand2_2 _30436_ (.A(_08805_),
    .B(_08806_),
    .Y(_08807_));
 sky130_fd_sc_hd__o21ai_2 _30437_ (.A1(_08537_),
    .A2(_08540_),
    .B1(_08535_),
    .Y(_08808_));
 sky130_vsdinv _30438_ (.A(_08808_),
    .Y(_08809_));
 sky130_fd_sc_hd__nand2_2 _30439_ (.A(_08807_),
    .B(_08809_),
    .Y(_08810_));
 sky130_fd_sc_hd__nand3_2 _30440_ (.A(_08805_),
    .B(_08806_),
    .C(_08808_),
    .Y(_08811_));
 sky130_fd_sc_hd__buf_1 _30441_ (.A(_19195_),
    .X(_08812_));
 sky130_fd_sc_hd__nand2_2 _30442_ (.A(_05513_),
    .B(_08812_),
    .Y(_08813_));
 sky130_fd_sc_hd__nand2_2 _30443_ (.A(_05509_),
    .B(_08570_),
    .Y(_08814_));
 sky130_fd_sc_hd__nor2_2 _30444_ (.A(_08813_),
    .B(_08814_),
    .Y(_08815_));
 sky130_fd_sc_hd__nand2_2 _30445_ (.A(_08813_),
    .B(_08814_),
    .Y(_08816_));
 sky130_vsdinv _30446_ (.A(_08816_),
    .Y(_08817_));
 sky130_fd_sc_hd__buf_1 _30447_ (.A(\pcpi_mul.rs1[25] ),
    .X(_08818_));
 sky130_fd_sc_hd__and2_2 _30448_ (.A(_18878_),
    .B(_08818_),
    .X(_08819_));
 sky130_fd_sc_hd__o21bai_2 _30449_ (.A1(_08815_),
    .A2(_08817_),
    .B1_N(_08819_),
    .Y(_08820_));
 sky130_fd_sc_hd__nand3b_2 _30450_ (.A_N(_08815_),
    .B(_08816_),
    .C(_08819_),
    .Y(_08821_));
 sky130_fd_sc_hd__nand2_2 _30451_ (.A(_08559_),
    .B(_08554_),
    .Y(_08822_));
 sky130_fd_sc_hd__a21o_2 _30452_ (.A1(_08820_),
    .A2(_08821_),
    .B1(_08822_),
    .X(_08823_));
 sky130_fd_sc_hd__nand3_2 _30453_ (.A(_08822_),
    .B(_08820_),
    .C(_08821_),
    .Y(_08824_));
 sky130_fd_sc_hd__buf_1 _30454_ (.A(\pcpi_mul.rs1[22] ),
    .X(_08825_));
 sky130_fd_sc_hd__buf_1 _30455_ (.A(_08825_),
    .X(_08826_));
 sky130_fd_sc_hd__buf_1 _30456_ (.A(_08826_),
    .X(_08827_));
 sky130_fd_sc_hd__and2_2 _30457_ (.A(_06460_),
    .B(_08827_),
    .X(_08828_));
 sky130_fd_sc_hd__buf_1 _30458_ (.A(\pcpi_mul.rs1[23] ),
    .X(_08829_));
 sky130_fd_sc_hd__buf_1 _30459_ (.A(_08829_),
    .X(_08830_));
 sky130_fd_sc_hd__nand2_2 _30460_ (.A(_05835_),
    .B(_08830_),
    .Y(_08831_));
 sky130_fd_sc_hd__buf_1 _30461_ (.A(_19171_),
    .X(_08832_));
 sky130_fd_sc_hd__buf_1 _30462_ (.A(_08832_),
    .X(_08833_));
 sky130_fd_sc_hd__nand2_2 _30463_ (.A(_18872_),
    .B(_08833_),
    .Y(_08834_));
 sky130_fd_sc_hd__xnor2_2 _30464_ (.A(_08831_),
    .B(_08834_),
    .Y(_08835_));
 sky130_fd_sc_hd__xnor2_2 _30465_ (.A(_08828_),
    .B(_08835_),
    .Y(_08836_));
 sky130_fd_sc_hd__a21oi_2 _30466_ (.A1(_08823_),
    .A2(_08824_),
    .B1(_08836_),
    .Y(_08837_));
 sky130_fd_sc_hd__nand3_2 _30467_ (.A(_08836_),
    .B(_08823_),
    .C(_08824_),
    .Y(_08838_));
 sky130_vsdinv _30468_ (.A(_08838_),
    .Y(_08839_));
 sky130_fd_sc_hd__o21ai_2 _30469_ (.A1(_08576_),
    .A2(_08579_),
    .B1(_08564_),
    .Y(_08840_));
 sky130_fd_sc_hd__o21bai_2 _30470_ (.A1(_08837_),
    .A2(_08839_),
    .B1_N(_08840_),
    .Y(_08841_));
 sky130_fd_sc_hd__nand3b_2 _30471_ (.A_N(_08837_),
    .B(_08838_),
    .C(_08840_),
    .Y(_08842_));
 sky130_fd_sc_hd__nor2_2 _30472_ (.A(_08566_),
    .B(_08567_),
    .Y(_08843_));
 sky130_fd_sc_hd__a21oi_2 _30473_ (.A1(_08568_),
    .A2(_08572_),
    .B1(_08843_),
    .Y(_08844_));
 sky130_vsdinv _30474_ (.A(_08844_),
    .Y(_08845_));
 sky130_fd_sc_hd__a21oi_2 _30475_ (.A1(_08841_),
    .A2(_08842_),
    .B1(_08845_),
    .Y(_08846_));
 sky130_fd_sc_hd__nand3_2 _30476_ (.A(_08841_),
    .B(_08845_),
    .C(_08842_),
    .Y(_08847_));
 sky130_vsdinv _30477_ (.A(_08847_),
    .Y(_08848_));
 sky130_fd_sc_hd__nor2_2 _30478_ (.A(_08846_),
    .B(_08848_),
    .Y(_08849_));
 sky130_fd_sc_hd__a21oi_2 _30479_ (.A1(_08810_),
    .A2(_08811_),
    .B1(_08849_),
    .Y(_08850_));
 sky130_fd_sc_hd__or2b_2 _30480_ (.A(_08846_),
    .B_N(_08847_),
    .X(_08851_));
 sky130_fd_sc_hd__nand2_2 _30481_ (.A(_08810_),
    .B(_08811_),
    .Y(_08852_));
 sky130_fd_sc_hd__nor2_2 _30482_ (.A(_08851_),
    .B(_08852_),
    .Y(_08853_));
 sky130_fd_sc_hd__o21ai_2 _30483_ (.A1(_08451_),
    .A2(_08445_),
    .B1(_08455_),
    .Y(_08854_));
 sky130_fd_sc_hd__o21bai_2 _30484_ (.A1(_08850_),
    .A2(_08853_),
    .B1_N(_08854_),
    .Y(_08855_));
 sky130_fd_sc_hd__nand3_2 _30485_ (.A(_08849_),
    .B(_08810_),
    .C(_08811_),
    .Y(_08856_));
 sky130_fd_sc_hd__nand3b_2 _30486_ (.A_N(_08850_),
    .B(_08854_),
    .C(_08856_),
    .Y(_08857_));
 sky130_fd_sc_hd__nand2_2 _30487_ (.A(_08855_),
    .B(_08857_),
    .Y(_08858_));
 sky130_fd_sc_hd__a21oi_2 _30488_ (.A1(_08593_),
    .A2(_08544_),
    .B1(_08599_),
    .Y(_08859_));
 sky130_fd_sc_hd__nand2_2 _30489_ (.A(_08858_),
    .B(_08859_),
    .Y(_08860_));
 sky130_fd_sc_hd__buf_1 _30490_ (.A(_08860_),
    .X(_08861_));
 sky130_fd_sc_hd__nand3b_2 _30491_ (.A_N(_08859_),
    .B(_08855_),
    .C(_08857_),
    .Y(_08862_));
 sky130_fd_sc_hd__buf_1 _30492_ (.A(_08862_),
    .X(_08863_));
 sky130_fd_sc_hd__a22oi_2 _30493_ (.A1(_08779_),
    .A2(_08782_),
    .B1(_08861_),
    .B2(_08863_),
    .Y(_08864_));
 sky130_fd_sc_hd__nand2_2 _30494_ (.A(_08779_),
    .B(_08782_),
    .Y(_08865_));
 sky130_fd_sc_hd__nand2_2 _30495_ (.A(_08860_),
    .B(_08862_),
    .Y(_08866_));
 sky130_fd_sc_hd__nor2_2 _30496_ (.A(_08865_),
    .B(_08866_),
    .Y(_08867_));
 sky130_fd_sc_hd__a31oi_2 _30497_ (.A1(_08610_),
    .A2(_08503_),
    .A3(_08607_),
    .B1(_08619_),
    .Y(_08868_));
 sky130_fd_sc_hd__o21ai_2 _30498_ (.A1(_08864_),
    .A2(_08867_),
    .B1(_08868_),
    .Y(_08869_));
 sky130_fd_sc_hd__and2_2 _30499_ (.A(_08778_),
    .B(_08782_),
    .X(_08870_));
 sky130_fd_sc_hd__nand3_2 _30500_ (.A(_08870_),
    .B(_08863_),
    .C(_08861_),
    .Y(_08871_));
 sky130_fd_sc_hd__a31o_2 _30501_ (.A1(_08609_),
    .A2(_08503_),
    .A3(_08606_),
    .B1(_08619_),
    .X(_08872_));
 sky130_fd_sc_hd__nand2_2 _30502_ (.A(_08866_),
    .B(_08865_),
    .Y(_08873_));
 sky130_fd_sc_hd__nand3_2 _30503_ (.A(_08871_),
    .B(_08872_),
    .C(_08873_),
    .Y(_08874_));
 sky130_fd_sc_hd__nand2_2 _30504_ (.A(_08869_),
    .B(_08874_),
    .Y(_08875_));
 sky130_fd_sc_hd__a21boi_2 _30505_ (.A1(_08583_),
    .A2(_08589_),
    .B1_N(_08587_),
    .Y(_08876_));
 sky130_fd_sc_hd__a21oi_2 _30506_ (.A1(_08607_),
    .A2(_08605_),
    .B1(_08876_),
    .Y(_08877_));
 sky130_fd_sc_hd__and3_2 _30507_ (.A(_08606_),
    .B(_08605_),
    .C(_08876_),
    .X(_08878_));
 sky130_fd_sc_hd__nor2_2 _30508_ (.A(_08877_),
    .B(_08878_),
    .Y(_08879_));
 sky130_vsdinv _30509_ (.A(_08879_),
    .Y(_08880_));
 sky130_fd_sc_hd__nand2_2 _30510_ (.A(_08875_),
    .B(_08880_),
    .Y(_08881_));
 sky130_fd_sc_hd__nand3_2 _30511_ (.A(_08869_),
    .B(_08874_),
    .C(_08879_),
    .Y(_08882_));
 sky130_fd_sc_hd__nand2_2 _30512_ (.A(_08881_),
    .B(_08882_),
    .Y(_08883_));
 sky130_fd_sc_hd__a21boi_2 _30513_ (.A1(_08616_),
    .A2(_08627_),
    .B1_N(_08623_),
    .Y(_08884_));
 sky130_fd_sc_hd__nand2_2 _30514_ (.A(_08883_),
    .B(_08884_),
    .Y(_08885_));
 sky130_fd_sc_hd__nand2_2 _30515_ (.A(_08630_),
    .B(_08623_),
    .Y(_08886_));
 sky130_fd_sc_hd__nand3_2 _30516_ (.A(_08886_),
    .B(_08881_),
    .C(_08882_),
    .Y(_08887_));
 sky130_fd_sc_hd__a21oi_2 _30517_ (.A1(_08344_),
    .A2(_08342_),
    .B1(_08625_),
    .Y(_08888_));
 sky130_fd_sc_hd__a21oi_2 _30518_ (.A1(_08885_),
    .A2(_08887_),
    .B1(_08888_),
    .Y(_08889_));
 sky130_vsdinv _30519_ (.A(_08888_),
    .Y(_08890_));
 sky130_fd_sc_hd__a21oi_2 _30520_ (.A1(_08881_),
    .A2(_08882_),
    .B1(_08886_),
    .Y(_08891_));
 sky130_fd_sc_hd__nor3b_2 _30521_ (.A(_08890_),
    .B(_08891_),
    .C_N(_08887_),
    .Y(_08892_));
 sky130_fd_sc_hd__o21ai_2 _30522_ (.A1(_08638_),
    .A2(_08639_),
    .B1(_08635_),
    .Y(_08893_));
 sky130_fd_sc_hd__o21bai_2 _30523_ (.A1(_08889_),
    .A2(_08892_),
    .B1_N(_08893_),
    .Y(_08894_));
 sky130_fd_sc_hd__nor2_2 _30524_ (.A(_08884_),
    .B(_08883_),
    .Y(_08895_));
 sky130_fd_sc_hd__o21bai_2 _30525_ (.A1(_08891_),
    .A2(_08895_),
    .B1_N(_08888_),
    .Y(_08896_));
 sky130_fd_sc_hd__nand3_2 _30526_ (.A(_08885_),
    .B(_08888_),
    .C(_08887_),
    .Y(_08897_));
 sky130_fd_sc_hd__nand3_2 _30527_ (.A(_08896_),
    .B(_08893_),
    .C(_08897_),
    .Y(_08898_));
 sky130_fd_sc_hd__nand2_2 _30528_ (.A(_08894_),
    .B(_08898_),
    .Y(_08899_));
 sky130_fd_sc_hd__o21ai_2 _30529_ (.A1(_08649_),
    .A2(_08657_),
    .B1(_08648_),
    .Y(_08900_));
 sky130_fd_sc_hd__xnor2_2 _30530_ (.A(_08899_),
    .B(_08900_),
    .Y(_02644_));
 sky130_fd_sc_hd__a22oi_2 _30531_ (.A1(_07786_),
    .A2(_05958_),
    .B1(_07788_),
    .B2(_06063_),
    .Y(_08901_));
 sky130_fd_sc_hd__nand2_2 _30532_ (.A(_18779_),
    .B(_05949_),
    .Y(_08902_));
 sky130_fd_sc_hd__nand2_2 _30533_ (.A(_07168_),
    .B(_06068_),
    .Y(_08903_));
 sky130_fd_sc_hd__nor2_2 _30534_ (.A(_08902_),
    .B(_08903_),
    .Y(_08904_));
 sky130_fd_sc_hd__buf_1 _30535_ (.A(_06201_),
    .X(_08905_));
 sky130_fd_sc_hd__and2_2 _30536_ (.A(_06665_),
    .B(_08905_),
    .X(_08906_));
 sky130_fd_sc_hd__o21bai_2 _30537_ (.A1(_08901_),
    .A2(_08904_),
    .B1_N(_08906_),
    .Y(_08907_));
 sky130_fd_sc_hd__buf_1 _30538_ (.A(_07787_),
    .X(_08908_));
 sky130_fd_sc_hd__nand3b_2 _30539_ (.A_N(_08902_),
    .B(_08908_),
    .C(_06883_),
    .Y(_08909_));
 sky130_fd_sc_hd__nand2_2 _30540_ (.A(_08902_),
    .B(_08903_),
    .Y(_08910_));
 sky130_fd_sc_hd__nand3_2 _30541_ (.A(_08909_),
    .B(_08906_),
    .C(_08910_),
    .Y(_08911_));
 sky130_fd_sc_hd__nand2_2 _30542_ (.A(_08907_),
    .B(_08911_),
    .Y(_08912_));
 sky130_fd_sc_hd__a21o_2 _30543_ (.A1(_08741_),
    .A2(_08745_),
    .B1(_08742_),
    .X(_08913_));
 sky130_vsdinv _30544_ (.A(_08913_),
    .Y(_08914_));
 sky130_fd_sc_hd__nand2_2 _30545_ (.A(_08912_),
    .B(_08914_),
    .Y(_08915_));
 sky130_fd_sc_hd__nand3_2 _30546_ (.A(_08907_),
    .B(_08913_),
    .C(_08911_),
    .Y(_08916_));
 sky130_fd_sc_hd__nand2_2 _30547_ (.A(_08915_),
    .B(_08916_),
    .Y(_08917_));
 sky130_fd_sc_hd__buf_1 _30548_ (.A(_18791_),
    .X(_08918_));
 sky130_fd_sc_hd__o31ai_2 _30549_ (.A1(_08918_),
    .A2(_19253_),
    .A3(_08658_),
    .B1(_08664_),
    .Y(_08919_));
 sky130_vsdinv _30550_ (.A(_08919_),
    .Y(_08920_));
 sky130_fd_sc_hd__nand2_2 _30551_ (.A(_08917_),
    .B(_08920_),
    .Y(_08921_));
 sky130_fd_sc_hd__nand3_2 _30552_ (.A(_08915_),
    .B(_08919_),
    .C(_08916_),
    .Y(_08922_));
 sky130_fd_sc_hd__nand2_2 _30553_ (.A(_08921_),
    .B(_08922_),
    .Y(_08923_));
 sky130_fd_sc_hd__a21boi_2 _30554_ (.A1(_08668_),
    .A2(_08674_),
    .B1_N(_08670_),
    .Y(_08924_));
 sky130_fd_sc_hd__nand2_2 _30555_ (.A(_08923_),
    .B(_08924_),
    .Y(_08925_));
 sky130_fd_sc_hd__nand2_2 _30556_ (.A(_08675_),
    .B(_08670_),
    .Y(_08926_));
 sky130_fd_sc_hd__nand3_2 _30557_ (.A(_08926_),
    .B(_08922_),
    .C(_08921_),
    .Y(_08927_));
 sky130_fd_sc_hd__buf_1 _30558_ (.A(_08927_),
    .X(_08928_));
 sky130_fd_sc_hd__nand2_2 _30559_ (.A(_08925_),
    .B(_08928_),
    .Y(_08929_));
 sky130_fd_sc_hd__nand2_2 _30560_ (.A(_18797_),
    .B(_06477_),
    .Y(_08930_));
 sky130_fd_sc_hd__nand2_2 _30561_ (.A(_06536_),
    .B(_07551_),
    .Y(_08931_));
 sky130_fd_sc_hd__nor2_2 _30562_ (.A(_08930_),
    .B(_08931_),
    .Y(_08932_));
 sky130_fd_sc_hd__and2_2 _30563_ (.A(_08038_),
    .B(_19231_),
    .X(_08933_));
 sky130_fd_sc_hd__nand2_2 _30564_ (.A(_08930_),
    .B(_08931_),
    .Y(_08934_));
 sky130_fd_sc_hd__nand3b_2 _30565_ (.A_N(_08932_),
    .B(_08933_),
    .C(_08934_),
    .Y(_08935_));
 sky130_fd_sc_hd__a22oi_2 _30566_ (.A1(_08032_),
    .A2(_06187_),
    .B1(_08034_),
    .B2(_07557_),
    .Y(_08936_));
 sky130_fd_sc_hd__o21bai_2 _30567_ (.A1(_08936_),
    .A2(_08932_),
    .B1_N(_08933_),
    .Y(_08937_));
 sky130_fd_sc_hd__a21oi_2 _30568_ (.A1(_08686_),
    .A2(_08685_),
    .B1(_08684_),
    .Y(_08938_));
 sky130_fd_sc_hd__a21boi_2 _30569_ (.A1(_08935_),
    .A2(_08937_),
    .B1_N(_08938_),
    .Y(_08939_));
 sky130_fd_sc_hd__nand3b_2 _30570_ (.A_N(_08938_),
    .B(_08935_),
    .C(_08937_),
    .Y(_08940_));
 sky130_vsdinv _30571_ (.A(_08940_),
    .Y(_08941_));
 sky130_fd_sc_hd__nand2_2 _30572_ (.A(_18813_),
    .B(_08261_),
    .Y(_08942_));
 sky130_fd_sc_hd__nand2_2 _30573_ (.A(_18818_),
    .B(_19215_),
    .Y(_08943_));
 sky130_fd_sc_hd__nand2_2 _30574_ (.A(_08942_),
    .B(_08943_),
    .Y(_08944_));
 sky130_fd_sc_hd__nor2_2 _30575_ (.A(_08942_),
    .B(_08943_),
    .Y(_08945_));
 sky130_vsdinv _30576_ (.A(_08945_),
    .Y(_08946_));
 sky130_fd_sc_hd__o2bb2ai_2 _30577_ (.A1_N(_08944_),
    .A2_N(_08946_),
    .B1(_07214_),
    .B2(_08524_),
    .Y(_08947_));
 sky130_fd_sc_hd__and2_2 _30578_ (.A(_06136_),
    .B(_07946_),
    .X(_08948_));
 sky130_fd_sc_hd__nand3b_2 _30579_ (.A_N(_08945_),
    .B(_08948_),
    .C(_08944_),
    .Y(_08949_));
 sky130_fd_sc_hd__nand2_2 _30580_ (.A(_08947_),
    .B(_08949_),
    .Y(_08950_));
 sky130_fd_sc_hd__o21ai_2 _30581_ (.A1(_08939_),
    .A2(_08941_),
    .B1(_08950_),
    .Y(_08951_));
 sky130_fd_sc_hd__nand2_2 _30582_ (.A(_08935_),
    .B(_08937_),
    .Y(_08952_));
 sky130_fd_sc_hd__nand2_2 _30583_ (.A(_08952_),
    .B(_08938_),
    .Y(_08953_));
 sky130_fd_sc_hd__nand3b_2 _30584_ (.A_N(_08950_),
    .B(_08940_),
    .C(_08953_),
    .Y(_08954_));
 sky130_fd_sc_hd__nand2_2 _30585_ (.A(_08951_),
    .B(_08954_),
    .Y(_08955_));
 sky130_fd_sc_hd__buf_1 _30586_ (.A(_08955_),
    .X(_08956_));
 sky130_fd_sc_hd__nand2_2 _30587_ (.A(_08929_),
    .B(_08956_),
    .Y(_08957_));
 sky130_fd_sc_hd__nand3b_2 _30588_ (.A_N(_08956_),
    .B(_08925_),
    .C(_08928_),
    .Y(_08958_));
 sky130_fd_sc_hd__a21oi_2 _30589_ (.A1(_08957_),
    .A2(_08958_),
    .B1(_08753_),
    .Y(_08959_));
 sky130_fd_sc_hd__a21boi_2 _30590_ (.A1(_08925_),
    .A2(_08928_),
    .B1_N(_08956_),
    .Y(_08960_));
 sky130_fd_sc_hd__a21oi_2 _30591_ (.A1(_08921_),
    .A2(_08922_),
    .B1(_08926_),
    .Y(_08961_));
 sky130_fd_sc_hd__nor3b_2 _30592_ (.A(_08956_),
    .B(_08961_),
    .C_N(_08928_),
    .Y(_08962_));
 sky130_fd_sc_hd__nor3_2 _30593_ (.A(_08752_),
    .B(_08960_),
    .C(_08962_),
    .Y(_08963_));
 sky130_fd_sc_hd__o21a_2 _30594_ (.A1(_08706_),
    .A2(_08677_),
    .B1(_08709_),
    .X(_08964_));
 sky130_vsdinv _30595_ (.A(_08964_),
    .Y(_08965_));
 sky130_fd_sc_hd__o21bai_2 _30596_ (.A1(_08959_),
    .A2(_08963_),
    .B1_N(_08965_),
    .Y(_08966_));
 sky130_fd_sc_hd__o21bai_2 _30597_ (.A1(_08960_),
    .A2(_08962_),
    .B1_N(_08753_),
    .Y(_08967_));
 sky130_fd_sc_hd__nand3_2 _30598_ (.A(_08957_),
    .B(_08753_),
    .C(_08958_),
    .Y(_08968_));
 sky130_fd_sc_hd__nand3_2 _30599_ (.A(_08967_),
    .B(_08965_),
    .C(_08968_),
    .Y(_08969_));
 sky130_fd_sc_hd__nand2_2 _30600_ (.A(_08471_),
    .B(_05986_),
    .Y(_08970_));
 sky130_fd_sc_hd__buf_1 _30601_ (.A(\pcpi_mul.rs2[22] ),
    .X(_08971_));
 sky130_fd_sc_hd__nand2_2 _30602_ (.A(_08971_),
    .B(_05532_),
    .Y(_08972_));
 sky130_fd_sc_hd__nor2_2 _30603_ (.A(_08970_),
    .B(_08972_),
    .Y(_08973_));
 sky130_fd_sc_hd__and2_2 _30604_ (.A(_08234_),
    .B(_19277_),
    .X(_08974_));
 sky130_fd_sc_hd__nand2_2 _30605_ (.A(_08970_),
    .B(_08972_),
    .Y(_08975_));
 sky130_fd_sc_hd__nand3b_2 _30606_ (.A_N(_08973_),
    .B(_08974_),
    .C(_08975_),
    .Y(_08976_));
 sky130_fd_sc_hd__a22oi_2 _30607_ (.A1(_08226_),
    .A2(_05644_),
    .B1(_18753_),
    .B2(_05533_),
    .Y(_08977_));
 sky130_fd_sc_hd__o21bai_2 _30608_ (.A1(_08977_),
    .A2(_08973_),
    .B1_N(_08974_),
    .Y(_08978_));
 sky130_fd_sc_hd__nand2_2 _30609_ (.A(_08976_),
    .B(_08978_),
    .Y(_08979_));
 sky130_fd_sc_hd__a21oi_2 _30610_ (.A1(_08727_),
    .A2(_08726_),
    .B1(_08724_),
    .Y(_08980_));
 sky130_fd_sc_hd__nand2_2 _30611_ (.A(_08979_),
    .B(_08980_),
    .Y(_08981_));
 sky130_fd_sc_hd__nand3b_2 _30612_ (.A_N(_08980_),
    .B(_08976_),
    .C(_08978_),
    .Y(_08982_));
 sky130_fd_sc_hd__nand2_2 _30613_ (.A(_08981_),
    .B(_08982_),
    .Y(_08983_));
 sky130_fd_sc_hd__nand2_2 _30614_ (.A(_18764_),
    .B(_05930_),
    .Y(_08984_));
 sky130_fd_sc_hd__buf_1 _30615_ (.A(\pcpi_mul.rs2[19] ),
    .X(_08985_));
 sky130_fd_sc_hd__nand2_2 _30616_ (.A(_08985_),
    .B(_07208_),
    .Y(_08986_));
 sky130_fd_sc_hd__nor2_2 _30617_ (.A(_08984_),
    .B(_08986_),
    .Y(_08987_));
 sky130_fd_sc_hd__nand2_2 _30618_ (.A(_08984_),
    .B(_08986_),
    .Y(_08988_));
 sky130_vsdinv _30619_ (.A(_08988_),
    .Y(_08989_));
 sky130_fd_sc_hd__buf_1 _30620_ (.A(\pcpi_mul.rs2[18] ),
    .X(_08990_));
 sky130_fd_sc_hd__and2_2 _30621_ (.A(_08990_),
    .B(_05846_),
    .X(_08991_));
 sky130_fd_sc_hd__o21bai_2 _30622_ (.A1(_08987_),
    .A2(_08989_),
    .B1_N(_08991_),
    .Y(_08992_));
 sky130_fd_sc_hd__nand3b_2 _30623_ (.A_N(_08987_),
    .B(_08991_),
    .C(_08988_),
    .Y(_08993_));
 sky130_fd_sc_hd__nand2_2 _30624_ (.A(_08992_),
    .B(_08993_),
    .Y(_08994_));
 sky130_fd_sc_hd__nand2_2 _30625_ (.A(_08983_),
    .B(_08994_),
    .Y(_08995_));
 sky130_fd_sc_hd__nand3b_2 _30626_ (.A_N(_08994_),
    .B(_08981_),
    .C(_08982_),
    .Y(_08996_));
 sky130_fd_sc_hd__a21boi_2 _30627_ (.A1(_08728_),
    .A2(_08733_),
    .B1_N(_08735_),
    .Y(_08997_));
 sky130_fd_sc_hd__o21ai_2 _30628_ (.A1(_08747_),
    .A2(_08997_),
    .B1(_08737_),
    .Y(_08998_));
 sky130_fd_sc_hd__a21o_2 _30629_ (.A1(_08995_),
    .A2(_08996_),
    .B1(_08998_),
    .X(_08999_));
 sky130_fd_sc_hd__nand3_2 _30630_ (.A(_08995_),
    .B(_08998_),
    .C(_08996_),
    .Y(_09000_));
 sky130_fd_sc_hd__buf_1 _30631_ (.A(_09000_),
    .X(_09001_));
 sky130_fd_sc_hd__nor2_2 _30632_ (.A(_08757_),
    .B(_08760_),
    .Y(_09002_));
 sky130_vsdinv _30633_ (.A(_09002_),
    .Y(_09003_));
 sky130_fd_sc_hd__nand2_2 _30634_ (.A(_08755_),
    .B(_19297_),
    .Y(_09004_));
 sky130_fd_sc_hd__buf_1 _30635_ (.A(\pcpi_mul.rs2[26] ),
    .X(_09005_));
 sky130_fd_sc_hd__buf_1 _30636_ (.A(_09005_),
    .X(_09006_));
 sky130_fd_sc_hd__nand2_2 _30637_ (.A(_09006_),
    .B(_05238_),
    .Y(_09007_));
 sky130_fd_sc_hd__nand2_2 _30638_ (.A(_09004_),
    .B(_09007_),
    .Y(_09008_));
 sky130_fd_sc_hd__nor2_2 _30639_ (.A(_09004_),
    .B(_09007_),
    .Y(_09009_));
 sky130_vsdinv _30640_ (.A(_09009_),
    .Y(_09010_));
 sky130_fd_sc_hd__buf_1 _30641_ (.A(_18740_),
    .X(_09011_));
 sky130_fd_sc_hd__o2bb2ai_2 _30642_ (.A1_N(_09008_),
    .A2_N(_09010_),
    .B1(_09011_),
    .B2(_19294_),
    .Y(_09012_));
 sky130_fd_sc_hd__and2_2 _30643_ (.A(_08758_),
    .B(_05984_),
    .X(_09013_));
 sky130_fd_sc_hd__nand3b_2 _30644_ (.A_N(_09009_),
    .B(_09013_),
    .C(_09008_),
    .Y(_09014_));
 sky130_fd_sc_hd__nand2_2 _30645_ (.A(_09012_),
    .B(_09014_),
    .Y(_09015_));
 sky130_fd_sc_hd__xor2_2 _30646_ (.A(_09003_),
    .B(_09015_),
    .X(_09016_));
 sky130_fd_sc_hd__a21o_2 _30647_ (.A1(_08999_),
    .A2(_09001_),
    .B1(_09016_),
    .X(_09017_));
 sky130_fd_sc_hd__nand3_2 _30648_ (.A(_08999_),
    .B(_09016_),
    .C(_09000_),
    .Y(_09018_));
 sky130_fd_sc_hd__a21oi_2 _30649_ (.A1(_09017_),
    .A2(_09018_),
    .B1(_08769_),
    .Y(_09019_));
 sky130_fd_sc_hd__a21oi_2 _30650_ (.A1(_08999_),
    .A2(_09001_),
    .B1(_09016_),
    .Y(_09020_));
 sky130_vsdinv _30651_ (.A(_09018_),
    .Y(_09021_));
 sky130_fd_sc_hd__nor3_2 _30652_ (.A(_08764_),
    .B(_09020_),
    .C(_09021_),
    .Y(_09022_));
 sky130_fd_sc_hd__nor2_2 _30653_ (.A(_09019_),
    .B(_09022_),
    .Y(_09023_));
 sky130_fd_sc_hd__a21oi_2 _30654_ (.A1(_08966_),
    .A2(_08969_),
    .B1(_09023_),
    .Y(_09024_));
 sky130_fd_sc_hd__buf_1 _30655_ (.A(_09021_),
    .X(_09025_));
 sky130_fd_sc_hd__o21ai_2 _30656_ (.A1(_09020_),
    .A2(_09025_),
    .B1(_08765_),
    .Y(_09026_));
 sky130_fd_sc_hd__nand3b_2 _30657_ (.A_N(_08765_),
    .B(_09017_),
    .C(_09018_),
    .Y(_09027_));
 sky130_fd_sc_hd__nand2_2 _30658_ (.A(_09026_),
    .B(_09027_),
    .Y(_09028_));
 sky130_fd_sc_hd__a21oi_2 _30659_ (.A1(_08967_),
    .A2(_08968_),
    .B1(_08965_),
    .Y(_09029_));
 sky130_vsdinv _30660_ (.A(_08969_),
    .Y(_09030_));
 sky130_fd_sc_hd__nor3_2 _30661_ (.A(_09028_),
    .B(_09029_),
    .C(_09030_),
    .Y(_09031_));
 sky130_fd_sc_hd__a31oi_2 _30662_ (.A1(_08717_),
    .A2(_08721_),
    .A3(_08773_),
    .B1(_08770_),
    .Y(_09032_));
 sky130_fd_sc_hd__o21ai_2 _30663_ (.A1(_09024_),
    .A2(_09031_),
    .B1(_09032_),
    .Y(_09033_));
 sky130_fd_sc_hd__nand2_2 _30664_ (.A(_08781_),
    .B(_08774_),
    .Y(_09034_));
 sky130_fd_sc_hd__nand3_2 _30665_ (.A(_08966_),
    .B(_09023_),
    .C(_08969_),
    .Y(_09035_));
 sky130_fd_sc_hd__o21bai_2 _30666_ (.A1(_09029_),
    .A2(_09030_),
    .B1_N(_09023_),
    .Y(_09036_));
 sky130_fd_sc_hd__nand3_2 _30667_ (.A(_09034_),
    .B(_09035_),
    .C(_09036_),
    .Y(_09037_));
 sky130_fd_sc_hd__nand2_2 _30668_ (.A(_07058_),
    .B(_07324_),
    .Y(_09038_));
 sky130_fd_sc_hd__nand2_2 _30669_ (.A(_06095_),
    .B(_07309_),
    .Y(_09039_));
 sky130_fd_sc_hd__nor2_2 _30670_ (.A(_09038_),
    .B(_09039_),
    .Y(_09040_));
 sky130_fd_sc_hd__and2_2 _30671_ (.A(_18838_),
    .B(_07960_),
    .X(_09041_));
 sky130_fd_sc_hd__nand2_2 _30672_ (.A(_09038_),
    .B(_09039_),
    .Y(_09042_));
 sky130_fd_sc_hd__nand3b_2 _30673_ (.A_N(_09040_),
    .B(_09041_),
    .C(_09042_),
    .Y(_09043_));
 sky130_fd_sc_hd__a22oi_2 _30674_ (.A1(_07059_),
    .A2(_08299_),
    .B1(_06096_),
    .B2(_08551_),
    .Y(_09044_));
 sky130_fd_sc_hd__o21bai_2 _30675_ (.A1(_09044_),
    .A2(_09040_),
    .B1_N(_09041_),
    .Y(_09045_));
 sky130_fd_sc_hd__nand2_2 _30676_ (.A(_09043_),
    .B(_09045_),
    .Y(_09046_));
 sky130_fd_sc_hd__a21oi_2 _30677_ (.A1(_08697_),
    .A2(_08701_),
    .B1(_08698_),
    .Y(_09047_));
 sky130_fd_sc_hd__nand2_2 _30678_ (.A(_09046_),
    .B(_09047_),
    .Y(_09048_));
 sky130_fd_sc_hd__nand3b_2 _30679_ (.A_N(_09047_),
    .B(_09043_),
    .C(_09045_),
    .Y(_09049_));
 sky130_fd_sc_hd__o31a_2 _30680_ (.A1(_18839_),
    .A2(_19204_),
    .A3(_08783_),
    .B1(_08788_),
    .X(_09050_));
 sky130_vsdinv _30681_ (.A(_09050_),
    .Y(_09051_));
 sky130_fd_sc_hd__a21oi_2 _30682_ (.A1(_09048_),
    .A2(_09049_),
    .B1(_09051_),
    .Y(_09052_));
 sky130_fd_sc_hd__nand3_2 _30683_ (.A(_09048_),
    .B(_09051_),
    .C(_09049_),
    .Y(_09053_));
 sky130_vsdinv _30684_ (.A(_09053_),
    .Y(_09054_));
 sky130_fd_sc_hd__a21boi_2 _30685_ (.A1(_08687_),
    .A2(_08690_),
    .B1_N(_08691_),
    .Y(_09055_));
 sky130_fd_sc_hd__o21ai_2 _30686_ (.A1(_08703_),
    .A2(_09055_),
    .B1(_08693_),
    .Y(_09056_));
 sky130_fd_sc_hd__o21bai_2 _30687_ (.A1(_09052_),
    .A2(_09054_),
    .B1_N(_09056_),
    .Y(_09057_));
 sky130_fd_sc_hd__a21o_2 _30688_ (.A1(_09048_),
    .A2(_09049_),
    .B1(_09051_),
    .X(_09058_));
 sky130_fd_sc_hd__nand3_2 _30689_ (.A(_09058_),
    .B(_09056_),
    .C(_09053_),
    .Y(_09059_));
 sky130_fd_sc_hd__a21boi_2 _30690_ (.A1(_08792_),
    .A2(_08795_),
    .B1_N(_08793_),
    .Y(_09060_));
 sky130_fd_sc_hd__buf_1 _30691_ (.A(_09060_),
    .X(_09061_));
 sky130_fd_sc_hd__a21boi_2 _30692_ (.A1(_09057_),
    .A2(_09059_),
    .B1_N(_09061_),
    .Y(_09062_));
 sky130_fd_sc_hd__nand2_2 _30693_ (.A(_09057_),
    .B(_09059_),
    .Y(_09063_));
 sky130_fd_sc_hd__nor2_2 _30694_ (.A(_09061_),
    .B(_09063_),
    .Y(_09064_));
 sky130_fd_sc_hd__a21oi_2 _30695_ (.A1(_08801_),
    .A2(_08797_),
    .B1(_08799_),
    .Y(_09065_));
 sky130_fd_sc_hd__o21ai_2 _30696_ (.A1(_08804_),
    .A2(_09065_),
    .B1(_08802_),
    .Y(_09066_));
 sky130_fd_sc_hd__o21bai_2 _30697_ (.A1(_09062_),
    .A2(_09064_),
    .B1_N(_09066_),
    .Y(_09067_));
 sky130_fd_sc_hd__nand2_2 _30698_ (.A(_09063_),
    .B(_09061_),
    .Y(_09068_));
 sky130_fd_sc_hd__nand3b_2 _30699_ (.A_N(_09061_),
    .B(_09057_),
    .C(_09059_),
    .Y(_09069_));
 sky130_fd_sc_hd__nand3_2 _30700_ (.A(_09068_),
    .B(_09066_),
    .C(_09069_),
    .Y(_09070_));
 sky130_fd_sc_hd__nand2_2 _30701_ (.A(_05491_),
    .B(_07733_),
    .Y(_09071_));
 sky130_fd_sc_hd__buf_1 _30702_ (.A(_19184_),
    .X(_09072_));
 sky130_fd_sc_hd__nand2_2 _30703_ (.A(_18849_),
    .B(_09072_),
    .Y(_09073_));
 sky130_fd_sc_hd__nor2_2 _30704_ (.A(_09071_),
    .B(_09073_),
    .Y(_09074_));
 sky130_fd_sc_hd__and2_2 _30705_ (.A(_05647_),
    .B(_19161_),
    .X(_09075_));
 sky130_fd_sc_hd__nand2_2 _30706_ (.A(_09071_),
    .B(_09073_),
    .Y(_09076_));
 sky130_fd_sc_hd__nand3b_2 _30707_ (.A_N(_09074_),
    .B(_09075_),
    .C(_09076_),
    .Y(_09077_));
 sky130_fd_sc_hd__buf_1 _30708_ (.A(_19190_),
    .X(_09078_));
 sky130_fd_sc_hd__buf_1 _30709_ (.A(_09072_),
    .X(_09079_));
 sky130_fd_sc_hd__a22oi_2 _30710_ (.A1(_06051_),
    .A2(_09078_),
    .B1(_05463_),
    .B2(_09079_),
    .Y(_09080_));
 sky130_fd_sc_hd__o21bai_2 _30711_ (.A1(_09080_),
    .A2(_09074_),
    .B1_N(_09075_),
    .Y(_09081_));
 sky130_fd_sc_hd__a21oi_2 _30712_ (.A1(_08816_),
    .A2(_08819_),
    .B1(_08815_),
    .Y(_09082_));
 sky130_fd_sc_hd__a21bo_2 _30713_ (.A1(_09077_),
    .A2(_09081_),
    .B1_N(_09082_),
    .X(_09083_));
 sky130_fd_sc_hd__nand3b_2 _30714_ (.A_N(_09082_),
    .B(_09077_),
    .C(_09081_),
    .Y(_09084_));
 sky130_fd_sc_hd__nand2_2 _30715_ (.A(_05661_),
    .B(_08832_),
    .Y(_09085_));
 sky130_fd_sc_hd__buf_1 _30716_ (.A(\pcpi_mul.rs1[25] ),
    .X(_09086_));
 sky130_fd_sc_hd__nand2_2 _30717_ (.A(_05535_),
    .B(_09086_),
    .Y(_09087_));
 sky130_fd_sc_hd__xor2_2 _30718_ (.A(_09085_),
    .B(_09087_),
    .X(_09088_));
 sky130_fd_sc_hd__buf_1 _30719_ (.A(_08829_),
    .X(_09089_));
 sky130_fd_sc_hd__and2_2 _30720_ (.A(_05744_),
    .B(_09089_),
    .X(_09090_));
 sky130_fd_sc_hd__nand2_2 _30721_ (.A(_09088_),
    .B(_09090_),
    .Y(_09091_));
 sky130_fd_sc_hd__buf_1 _30722_ (.A(_19181_),
    .X(_09092_));
 sky130_fd_sc_hd__xnor2_2 _30723_ (.A(_09085_),
    .B(_09087_),
    .Y(_09093_));
 sky130_fd_sc_hd__o21ai_2 _30724_ (.A1(_07332_),
    .A2(_09092_),
    .B1(_09093_),
    .Y(_09094_));
 sky130_fd_sc_hd__nand2_2 _30725_ (.A(_09091_),
    .B(_09094_),
    .Y(_09095_));
 sky130_fd_sc_hd__a21boi_2 _30726_ (.A1(_09083_),
    .A2(_09084_),
    .B1_N(_09095_),
    .Y(_09096_));
 sky130_fd_sc_hd__nand3b_2 _30727_ (.A_N(_09095_),
    .B(_09084_),
    .C(_09083_),
    .Y(_09097_));
 sky130_vsdinv _30728_ (.A(_09097_),
    .Y(_09098_));
 sky130_fd_sc_hd__a21oi_2 _30729_ (.A1(_08820_),
    .A2(_08821_),
    .B1(_08822_),
    .Y(_09099_));
 sky130_fd_sc_hd__xor2_2 _30730_ (.A(_08828_),
    .B(_08835_),
    .X(_09100_));
 sky130_fd_sc_hd__o21ai_2 _30731_ (.A1(_09099_),
    .A2(_09100_),
    .B1(_08824_),
    .Y(_09101_));
 sky130_fd_sc_hd__o21bai_2 _30732_ (.A1(_09096_),
    .A2(_09098_),
    .B1_N(_09101_),
    .Y(_09102_));
 sky130_fd_sc_hd__nand3b_2 _30733_ (.A_N(_09096_),
    .B(_09097_),
    .C(_09101_),
    .Y(_09103_));
 sky130_fd_sc_hd__buf_1 _30734_ (.A(_19185_),
    .X(_09104_));
 sky130_fd_sc_hd__buf_1 _30735_ (.A(_09104_),
    .X(_09105_));
 sky130_fd_sc_hd__nand3b_2 _30736_ (.A_N(_08835_),
    .B(_05439_),
    .C(_09105_),
    .Y(_09106_));
 sky130_fd_sc_hd__o21a_2 _30737_ (.A1(_08831_),
    .A2(_08834_),
    .B1(_09106_),
    .X(_09107_));
 sky130_vsdinv _30738_ (.A(_09107_),
    .Y(_09108_));
 sky130_fd_sc_hd__a21oi_2 _30739_ (.A1(_09102_),
    .A2(_09103_),
    .B1(_09108_),
    .Y(_09109_));
 sky130_fd_sc_hd__nand3_2 _30740_ (.A(_09102_),
    .B(_09108_),
    .C(_09103_),
    .Y(_09110_));
 sky130_vsdinv _30741_ (.A(_09110_),
    .Y(_09111_));
 sky130_fd_sc_hd__nor2_2 _30742_ (.A(_09109_),
    .B(_09111_),
    .Y(_09112_));
 sky130_fd_sc_hd__a21oi_2 _30743_ (.A1(_09067_),
    .A2(_09070_),
    .B1(_09112_),
    .Y(_09113_));
 sky130_fd_sc_hd__nand2_2 _30744_ (.A(_09102_),
    .B(_09103_),
    .Y(_09114_));
 sky130_fd_sc_hd__nand2_2 _30745_ (.A(_09114_),
    .B(_09107_),
    .Y(_09115_));
 sky130_fd_sc_hd__nand2_2 _30746_ (.A(_09115_),
    .B(_09110_),
    .Y(_09116_));
 sky130_fd_sc_hd__a21oi_2 _30747_ (.A1(_09068_),
    .A2(_09069_),
    .B1(_09066_),
    .Y(_09117_));
 sky130_vsdinv _30748_ (.A(_09070_),
    .Y(_09118_));
 sky130_fd_sc_hd__nor3_2 _30749_ (.A(_09116_),
    .B(_09117_),
    .C(_09118_),
    .Y(_09119_));
 sky130_fd_sc_hd__o21ai_2 _30750_ (.A1(_08715_),
    .A2(_08712_),
    .B1(_08713_),
    .Y(_09120_));
 sky130_fd_sc_hd__o21bai_2 _30751_ (.A1(_09113_),
    .A2(_09119_),
    .B1_N(_09120_),
    .Y(_09121_));
 sky130_fd_sc_hd__o22ai_2 _30752_ (.A1(_09111_),
    .A2(_09109_),
    .B1(_09117_),
    .B2(_09118_),
    .Y(_09122_));
 sky130_fd_sc_hd__nand3_2 _30753_ (.A(_09112_),
    .B(_09067_),
    .C(_09070_),
    .Y(_09123_));
 sky130_fd_sc_hd__nand3_2 _30754_ (.A(_09122_),
    .B(_09123_),
    .C(_09120_),
    .Y(_09124_));
 sky130_fd_sc_hd__nand2_2 _30755_ (.A(_09121_),
    .B(_09124_),
    .Y(_09125_));
 sky130_fd_sc_hd__a21boi_2 _30756_ (.A1(_08849_),
    .A2(_08810_),
    .B1_N(_08811_),
    .Y(_09126_));
 sky130_fd_sc_hd__nand2_2 _30757_ (.A(_09125_),
    .B(_09126_),
    .Y(_09127_));
 sky130_fd_sc_hd__buf_1 _30758_ (.A(_09124_),
    .X(_09128_));
 sky130_fd_sc_hd__nand3b_2 _30759_ (.A_N(_09126_),
    .B(_09121_),
    .C(_09128_),
    .Y(_09129_));
 sky130_fd_sc_hd__buf_1 _30760_ (.A(_09129_),
    .X(_09130_));
 sky130_fd_sc_hd__a22oi_2 _30761_ (.A1(_09033_),
    .A2(_09037_),
    .B1(_09127_),
    .B2(_09130_),
    .Y(_09131_));
 sky130_fd_sc_hd__nand2_2 _30762_ (.A(_09033_),
    .B(_09037_),
    .Y(_09132_));
 sky130_fd_sc_hd__nand2_2 _30763_ (.A(_09127_),
    .B(_09130_),
    .Y(_09133_));
 sky130_fd_sc_hd__nor2_2 _30764_ (.A(_09132_),
    .B(_09133_),
    .Y(_09134_));
 sky130_vsdinv _30765_ (.A(_08782_),
    .Y(_09135_));
 sky130_fd_sc_hd__a31oi_2 _30766_ (.A1(_08861_),
    .A2(_08779_),
    .A3(_08863_),
    .B1(_09135_),
    .Y(_09136_));
 sky130_fd_sc_hd__o21ai_2 _30767_ (.A1(_09131_),
    .A2(_09134_),
    .B1(_09136_),
    .Y(_09137_));
 sky130_fd_sc_hd__a31o_2 _30768_ (.A1(_08861_),
    .A2(_08779_),
    .A3(_08862_),
    .B1(_09135_),
    .X(_09138_));
 sky130_fd_sc_hd__a21boi_2 _30769_ (.A1(_09121_),
    .A2(_09128_),
    .B1_N(_09126_),
    .Y(_09139_));
 sky130_fd_sc_hd__nor2_2 _30770_ (.A(_09126_),
    .B(_09125_),
    .Y(_09140_));
 sky130_fd_sc_hd__nor2_2 _30771_ (.A(_09139_),
    .B(_09140_),
    .Y(_09141_));
 sky130_fd_sc_hd__a21oi_2 _30772_ (.A1(_09036_),
    .A2(_09035_),
    .B1(_09034_),
    .Y(_09142_));
 sky130_fd_sc_hd__nor3_2 _30773_ (.A(_09024_),
    .B(_09031_),
    .C(_09032_),
    .Y(_09143_));
 sky130_fd_sc_hd__nor2_2 _30774_ (.A(_09142_),
    .B(_09143_),
    .Y(_09144_));
 sky130_fd_sc_hd__nand2_2 _30775_ (.A(_09141_),
    .B(_09144_),
    .Y(_09145_));
 sky130_fd_sc_hd__nand2_2 _30776_ (.A(_09133_),
    .B(_09132_),
    .Y(_09146_));
 sky130_fd_sc_hd__nand3_2 _30777_ (.A(_09138_),
    .B(_09145_),
    .C(_09146_),
    .Y(_09147_));
 sky130_fd_sc_hd__nand2_2 _30778_ (.A(_09137_),
    .B(_09147_),
    .Y(_09148_));
 sky130_fd_sc_hd__a21boi_2 _30779_ (.A1(_08841_),
    .A2(_08845_),
    .B1_N(_08842_),
    .Y(_09149_));
 sky130_fd_sc_hd__nand2_2 _30780_ (.A(_08862_),
    .B(_08857_),
    .Y(_09150_));
 sky130_fd_sc_hd__xor2_2 _30781_ (.A(_09149_),
    .B(_09150_),
    .X(_09151_));
 sky130_fd_sc_hd__nand2_2 _30782_ (.A(_09148_),
    .B(_09151_),
    .Y(_09152_));
 sky130_fd_sc_hd__nand3b_2 _30783_ (.A_N(_09151_),
    .B(_09137_),
    .C(_09147_),
    .Y(_09153_));
 sky130_fd_sc_hd__nand2_2 _30784_ (.A(_08882_),
    .B(_08874_),
    .Y(_09154_));
 sky130_fd_sc_hd__a21oi_2 _30785_ (.A1(_09152_),
    .A2(_09153_),
    .B1(_09154_),
    .Y(_09155_));
 sky130_fd_sc_hd__a21boi_2 _30786_ (.A1(_08869_),
    .A2(_08879_),
    .B1_N(_08874_),
    .Y(_09156_));
 sky130_fd_sc_hd__nand2_2 _30787_ (.A(_09152_),
    .B(_09153_),
    .Y(_09157_));
 sky130_fd_sc_hd__nor2_2 _30788_ (.A(_09156_),
    .B(_09157_),
    .Y(_09158_));
 sky130_fd_sc_hd__buf_1 _30789_ (.A(_08877_),
    .X(_09159_));
 sky130_fd_sc_hd__o21bai_2 _30790_ (.A1(_09155_),
    .A2(_09158_),
    .B1_N(_09159_),
    .Y(_09160_));
 sky130_fd_sc_hd__nand2_2 _30791_ (.A(_09157_),
    .B(_09156_),
    .Y(_09161_));
 sky130_fd_sc_hd__nand3_2 _30792_ (.A(_09154_),
    .B(_09153_),
    .C(_09152_),
    .Y(_09162_));
 sky130_fd_sc_hd__nand3_2 _30793_ (.A(_09161_),
    .B(_09159_),
    .C(_09162_),
    .Y(_09163_));
 sky130_fd_sc_hd__o21ai_2 _30794_ (.A1(_08890_),
    .A2(_08891_),
    .B1(_08887_),
    .Y(_09164_));
 sky130_fd_sc_hd__a21oi_2 _30795_ (.A1(_09160_),
    .A2(_09163_),
    .B1(_09164_),
    .Y(_09165_));
 sky130_fd_sc_hd__nand3_2 _30796_ (.A(_09160_),
    .B(_09163_),
    .C(_09164_),
    .Y(_09166_));
 sky130_vsdinv _30797_ (.A(_09166_),
    .Y(_09167_));
 sky130_fd_sc_hd__nor2_2 _30798_ (.A(_09165_),
    .B(_09167_),
    .Y(_09168_));
 sky130_fd_sc_hd__a21oi_2 _30799_ (.A1(_08896_),
    .A2(_08897_),
    .B1(_08893_),
    .Y(_09169_));
 sky130_fd_sc_hd__a21oi_2 _30800_ (.A1(_08648_),
    .A2(_08898_),
    .B1(_09169_),
    .Y(_09170_));
 sky130_vsdinv _30801_ (.A(_09170_),
    .Y(_09171_));
 sky130_fd_sc_hd__o31ai_2 _30802_ (.A1(_08649_),
    .A2(_08899_),
    .A3(_08657_),
    .B1(_09171_),
    .Y(_09172_));
 sky130_fd_sc_hd__xor2_2 _30803_ (.A(_09168_),
    .B(_09172_),
    .X(_02645_));
 sky130_fd_sc_hd__a22oi_2 _30804_ (.A1(_07059_),
    .A2(_19203_),
    .B1(_07271_),
    .B2(_19196_),
    .Y(_09173_));
 sky130_fd_sc_hd__nand2_2 _30805_ (.A(_06880_),
    .B(_19202_),
    .Y(_09174_));
 sky130_fd_sc_hd__nand2_2 _30806_ (.A(_05767_),
    .B(_07960_),
    .Y(_09175_));
 sky130_fd_sc_hd__nor2_2 _30807_ (.A(_09174_),
    .B(_09175_),
    .Y(_09176_));
 sky130_fd_sc_hd__and2_2 _30808_ (.A(_05585_),
    .B(_08569_),
    .X(_09177_));
 sky130_fd_sc_hd__o21bai_2 _30809_ (.A1(_09173_),
    .A2(_09176_),
    .B1_N(_09177_),
    .Y(_09178_));
 sky130_fd_sc_hd__nand3b_2 _30810_ (.A_N(_09174_),
    .B(_06096_),
    .C(_07591_),
    .Y(_09179_));
 sky130_fd_sc_hd__nand2_2 _30811_ (.A(_09174_),
    .B(_09175_),
    .Y(_09180_));
 sky130_fd_sc_hd__nand3_2 _30812_ (.A(_09179_),
    .B(_09177_),
    .C(_09180_),
    .Y(_09181_));
 sky130_fd_sc_hd__nand2_2 _30813_ (.A(_09178_),
    .B(_09181_),
    .Y(_09182_));
 sky130_fd_sc_hd__a21o_2 _30814_ (.A1(_08944_),
    .A2(_08948_),
    .B1(_08945_),
    .X(_09183_));
 sky130_vsdinv _30815_ (.A(_09183_),
    .Y(_09184_));
 sky130_fd_sc_hd__nand2_2 _30816_ (.A(_09182_),
    .B(_09184_),
    .Y(_09185_));
 sky130_fd_sc_hd__nand3_2 _30817_ (.A(_09178_),
    .B(_09183_),
    .C(_09181_),
    .Y(_09186_));
 sky130_fd_sc_hd__a21oi_2 _30818_ (.A1(_09042_),
    .A2(_09041_),
    .B1(_09040_),
    .Y(_09187_));
 sky130_vsdinv _30819_ (.A(_09187_),
    .Y(_09188_));
 sky130_fd_sc_hd__a21oi_2 _30820_ (.A1(_09185_),
    .A2(_09186_),
    .B1(_09188_),
    .Y(_09189_));
 sky130_fd_sc_hd__nand3_2 _30821_ (.A(_09185_),
    .B(_09188_),
    .C(_09186_),
    .Y(_09190_));
 sky130_vsdinv _30822_ (.A(_09190_),
    .Y(_09191_));
 sky130_fd_sc_hd__o21a_2 _30823_ (.A1(_08950_),
    .A2(_08939_),
    .B1(_08940_),
    .X(_09192_));
 sky130_fd_sc_hd__o21ai_2 _30824_ (.A1(_09189_),
    .A2(_09191_),
    .B1(_09192_),
    .Y(_09193_));
 sky130_fd_sc_hd__a21o_2 _30825_ (.A1(_09185_),
    .A2(_09186_),
    .B1(_09188_),
    .X(_09194_));
 sky130_fd_sc_hd__o21ai_2 _30826_ (.A1(_08950_),
    .A2(_08939_),
    .B1(_08940_),
    .Y(_09195_));
 sky130_fd_sc_hd__nand3_2 _30827_ (.A(_09194_),
    .B(_09195_),
    .C(_09190_),
    .Y(_09196_));
 sky130_fd_sc_hd__a21boi_2 _30828_ (.A1(_09048_),
    .A2(_09051_),
    .B1_N(_09049_),
    .Y(_09197_));
 sky130_vsdinv _30829_ (.A(_09197_),
    .Y(_09198_));
 sky130_fd_sc_hd__a21oi_2 _30830_ (.A1(_09193_),
    .A2(_09196_),
    .B1(_09198_),
    .Y(_09199_));
 sky130_fd_sc_hd__nand3_2 _30831_ (.A(_09193_),
    .B(_09198_),
    .C(_09196_),
    .Y(_09200_));
 sky130_vsdinv _30832_ (.A(_09200_),
    .Y(_09201_));
 sky130_fd_sc_hd__a21oi_2 _30833_ (.A1(_09058_),
    .A2(_09053_),
    .B1(_09056_),
    .Y(_09202_));
 sky130_fd_sc_hd__o21ai_2 _30834_ (.A1(_09060_),
    .A2(_09202_),
    .B1(_09059_),
    .Y(_09203_));
 sky130_fd_sc_hd__o21bai_2 _30835_ (.A1(_09199_),
    .A2(_09201_),
    .B1_N(_09203_),
    .Y(_09204_));
 sky130_fd_sc_hd__nand2_2 _30836_ (.A(_09193_),
    .B(_09196_),
    .Y(_09205_));
 sky130_fd_sc_hd__nand2_2 _30837_ (.A(_09205_),
    .B(_09197_),
    .Y(_09206_));
 sky130_fd_sc_hd__nand3_2 _30838_ (.A(_09206_),
    .B(_09203_),
    .C(_09200_),
    .Y(_09207_));
 sky130_fd_sc_hd__buf_1 _30839_ (.A(_09207_),
    .X(_09208_));
 sky130_fd_sc_hd__nand2_2 _30840_ (.A(_18843_),
    .B(_08825_),
    .Y(_09209_));
 sky130_fd_sc_hd__nand2_2 _30841_ (.A(_05637_),
    .B(_08829_),
    .Y(_09210_));
 sky130_fd_sc_hd__nor2_2 _30842_ (.A(_09209_),
    .B(_09210_),
    .Y(_09211_));
 sky130_fd_sc_hd__buf_1 _30843_ (.A(\pcpi_mul.rs1[27] ),
    .X(_09212_));
 sky130_fd_sc_hd__and2_2 _30844_ (.A(_05647_),
    .B(_09212_),
    .X(_09213_));
 sky130_fd_sc_hd__nand2_2 _30845_ (.A(_09209_),
    .B(_09210_),
    .Y(_09214_));
 sky130_fd_sc_hd__nand3b_2 _30846_ (.A_N(_09211_),
    .B(_09213_),
    .C(_09214_),
    .Y(_09215_));
 sky130_fd_sc_hd__buf_1 _30847_ (.A(_08825_),
    .X(_09216_));
 sky130_fd_sc_hd__a22oi_2 _30848_ (.A1(_05813_),
    .A2(_09216_),
    .B1(_05929_),
    .B2(_08295_),
    .Y(_09217_));
 sky130_fd_sc_hd__o21bai_2 _30849_ (.A1(_09217_),
    .A2(_09211_),
    .B1_N(_09213_),
    .Y(_09218_));
 sky130_fd_sc_hd__a21oi_2 _30850_ (.A1(_09076_),
    .A2(_09075_),
    .B1(_09074_),
    .Y(_09219_));
 sky130_fd_sc_hd__a21bo_2 _30851_ (.A1(_09215_),
    .A2(_09218_),
    .B1_N(_09219_),
    .X(_09220_));
 sky130_fd_sc_hd__nand3b_2 _30852_ (.A_N(_09219_),
    .B(_09215_),
    .C(_09218_),
    .Y(_09221_));
 sky130_fd_sc_hd__nand2_2 _30853_ (.A(_09220_),
    .B(_09221_),
    .Y(_09222_));
 sky130_fd_sc_hd__nand2_2 _30854_ (.A(_18865_),
    .B(_19166_),
    .Y(_09223_));
 sky130_fd_sc_hd__buf_1 _30855_ (.A(\pcpi_mul.rs1[26] ),
    .X(_09224_));
 sky130_fd_sc_hd__nand2_2 _30856_ (.A(_18871_),
    .B(_09224_),
    .Y(_09225_));
 sky130_fd_sc_hd__xor2_2 _30857_ (.A(_09223_),
    .B(_09225_),
    .X(_09226_));
 sky130_fd_sc_hd__and2_2 _30858_ (.A(_05437_),
    .B(_08557_),
    .X(_09227_));
 sky130_fd_sc_hd__nand2_2 _30859_ (.A(_09226_),
    .B(_09227_),
    .Y(_09228_));
 sky130_fd_sc_hd__xnor2_2 _30860_ (.A(_09223_),
    .B(_09225_),
    .Y(_09229_));
 sky130_fd_sc_hd__o21ai_2 _30861_ (.A1(_18856_),
    .A2(_19173_),
    .B1(_09229_),
    .Y(_09230_));
 sky130_fd_sc_hd__nand2_2 _30862_ (.A(_09228_),
    .B(_09230_),
    .Y(_09231_));
 sky130_fd_sc_hd__nand2_2 _30863_ (.A(_09222_),
    .B(_09231_),
    .Y(_09232_));
 sky130_fd_sc_hd__nand3b_2 _30864_ (.A_N(_09231_),
    .B(_09221_),
    .C(_09220_),
    .Y(_09233_));
 sky130_fd_sc_hd__nand2_2 _30865_ (.A(_09232_),
    .B(_09233_),
    .Y(_09234_));
 sky130_fd_sc_hd__a21boi_2 _30866_ (.A1(_09077_),
    .A2(_09081_),
    .B1_N(_09082_),
    .Y(_09235_));
 sky130_fd_sc_hd__o21ai_2 _30867_ (.A1(_09235_),
    .A2(_09095_),
    .B1(_09084_),
    .Y(_09236_));
 sky130_vsdinv _30868_ (.A(_09236_),
    .Y(_09237_));
 sky130_fd_sc_hd__nand2_2 _30869_ (.A(_09234_),
    .B(_09237_),
    .Y(_09238_));
 sky130_fd_sc_hd__nand3_2 _30870_ (.A(_09232_),
    .B(_09236_),
    .C(_09233_),
    .Y(_09239_));
 sky130_fd_sc_hd__nand2_2 _30871_ (.A(_09238_),
    .B(_09239_),
    .Y(_09240_));
 sky130_fd_sc_hd__nor2_2 _30872_ (.A(_09085_),
    .B(_09087_),
    .Y(_09241_));
 sky130_fd_sc_hd__a21oi_2 _30873_ (.A1(_09088_),
    .A2(_09090_),
    .B1(_09241_),
    .Y(_09242_));
 sky130_fd_sc_hd__nand2_2 _30874_ (.A(_09240_),
    .B(_09242_),
    .Y(_09243_));
 sky130_vsdinv _30875_ (.A(_09242_),
    .Y(_09244_));
 sky130_fd_sc_hd__nand3_2 _30876_ (.A(_09238_),
    .B(_09244_),
    .C(_09239_),
    .Y(_09245_));
 sky130_fd_sc_hd__and2_2 _30877_ (.A(_09243_),
    .B(_09245_),
    .X(_09246_));
 sky130_fd_sc_hd__a21oi_2 _30878_ (.A1(_09204_),
    .A2(_09208_),
    .B1(_09246_),
    .Y(_09247_));
 sky130_fd_sc_hd__nand2_2 _30879_ (.A(_09243_),
    .B(_09245_),
    .Y(_09248_));
 sky130_fd_sc_hd__a21oi_2 _30880_ (.A1(_09206_),
    .A2(_09200_),
    .B1(_09203_),
    .Y(_09249_));
 sky130_fd_sc_hd__nor3b_2 _30881_ (.A(_09248_),
    .B(_09249_),
    .C_N(_09208_),
    .Y(_09250_));
 sky130_fd_sc_hd__o21ai_2 _30882_ (.A1(_08964_),
    .A2(_08959_),
    .B1(_08968_),
    .Y(_09251_));
 sky130_fd_sc_hd__o21bai_2 _30883_ (.A1(_09247_),
    .A2(_09250_),
    .B1_N(_09251_),
    .Y(_09252_));
 sky130_fd_sc_hd__a21o_2 _30884_ (.A1(_09204_),
    .A2(_09207_),
    .B1(_09246_),
    .X(_09253_));
 sky130_fd_sc_hd__nand3_2 _30885_ (.A(_09246_),
    .B(_09204_),
    .C(_09208_),
    .Y(_09254_));
 sky130_fd_sc_hd__nand3_2 _30886_ (.A(_09253_),
    .B(_09251_),
    .C(_09254_),
    .Y(_09255_));
 sky130_fd_sc_hd__buf_1 _30887_ (.A(_09255_),
    .X(_09256_));
 sky130_fd_sc_hd__nand2_2 _30888_ (.A(_09252_),
    .B(_09256_),
    .Y(_09257_));
 sky130_fd_sc_hd__a21oi_2 _30889_ (.A1(_09112_),
    .A2(_09067_),
    .B1(_09118_),
    .Y(_09258_));
 sky130_fd_sc_hd__nand2_2 _30890_ (.A(_09257_),
    .B(_09258_),
    .Y(_09259_));
 sky130_vsdinv _30891_ (.A(_09258_),
    .Y(_09260_));
 sky130_fd_sc_hd__nand3_2 _30892_ (.A(_09252_),
    .B(_09260_),
    .C(_09255_),
    .Y(_09261_));
 sky130_fd_sc_hd__buf_1 _30893_ (.A(_09261_),
    .X(_09262_));
 sky130_fd_sc_hd__buf_1 _30894_ (.A(_18752_),
    .X(_09263_));
 sky130_fd_sc_hd__a22oi_2 _30895_ (.A1(_08226_),
    .A2(_05722_),
    .B1(_09263_),
    .B2(_08003_),
    .Y(_09264_));
 sky130_fd_sc_hd__nand2_2 _30896_ (.A(_18747_),
    .B(_19281_),
    .Y(_09265_));
 sky130_fd_sc_hd__buf_1 _30897_ (.A(\pcpi_mul.rs2[22] ),
    .X(_09266_));
 sky130_fd_sc_hd__nand2_2 _30898_ (.A(_09266_),
    .B(_08003_),
    .Y(_09267_));
 sky130_fd_sc_hd__nor2_2 _30899_ (.A(_09265_),
    .B(_09267_),
    .Y(_09268_));
 sky130_fd_sc_hd__nand2_2 _30900_ (.A(_18758_),
    .B(_05665_),
    .Y(_09269_));
 sky130_vsdinv _30901_ (.A(_09269_),
    .Y(_09270_));
 sky130_fd_sc_hd__o21bai_2 _30902_ (.A1(_09264_),
    .A2(_09268_),
    .B1_N(_09270_),
    .Y(_09271_));
 sky130_fd_sc_hd__buf_1 _30903_ (.A(_08971_),
    .X(_09272_));
 sky130_fd_sc_hd__nand3b_2 _30904_ (.A_N(_09265_),
    .B(_09272_),
    .C(_05518_),
    .Y(_09273_));
 sky130_fd_sc_hd__nand2_2 _30905_ (.A(_09265_),
    .B(_09267_),
    .Y(_09274_));
 sky130_fd_sc_hd__nand3_2 _30906_ (.A(_09273_),
    .B(_09270_),
    .C(_09274_),
    .Y(_09275_));
 sky130_fd_sc_hd__nand2_2 _30907_ (.A(_09271_),
    .B(_09275_),
    .Y(_09276_));
 sky130_fd_sc_hd__a21oi_2 _30908_ (.A1(_08975_),
    .A2(_08974_),
    .B1(_08973_),
    .Y(_09277_));
 sky130_fd_sc_hd__nand2_2 _30909_ (.A(_09276_),
    .B(_09277_),
    .Y(_09278_));
 sky130_fd_sc_hd__nand3b_2 _30910_ (.A_N(_09277_),
    .B(_09275_),
    .C(_09271_),
    .Y(_09279_));
 sky130_fd_sc_hd__nand2_2 _30911_ (.A(_09278_),
    .B(_09279_),
    .Y(_09280_));
 sky130_fd_sc_hd__nand2_2 _30912_ (.A(_07850_),
    .B(_06979_),
    .Y(_09281_));
 sky130_fd_sc_hd__nand2_2 _30913_ (.A(_08985_),
    .B(_19261_),
    .Y(_09282_));
 sky130_fd_sc_hd__nand2_2 _30914_ (.A(_09281_),
    .B(_09282_),
    .Y(_09283_));
 sky130_fd_sc_hd__nand3b_2 _30915_ (.A_N(_09281_),
    .B(_08215_),
    .C(_06181_),
    .Y(_09284_));
 sky130_fd_sc_hd__o2bb2ai_2 _30916_ (.A1_N(_09283_),
    .A2_N(_09284_),
    .B1(_18776_),
    .B2(_19259_),
    .Y(_09285_));
 sky130_fd_sc_hd__and2_2 _30917_ (.A(_08990_),
    .B(_06342_),
    .X(_09286_));
 sky130_fd_sc_hd__nand3_2 _30918_ (.A(_09284_),
    .B(_09286_),
    .C(_09283_),
    .Y(_09287_));
 sky130_fd_sc_hd__nand2_2 _30919_ (.A(_09285_),
    .B(_09287_),
    .Y(_09288_));
 sky130_fd_sc_hd__buf_1 _30920_ (.A(_09288_),
    .X(_09289_));
 sky130_fd_sc_hd__nand2_2 _30921_ (.A(_09280_),
    .B(_09289_),
    .Y(_09290_));
 sky130_fd_sc_hd__nand3b_2 _30922_ (.A_N(_09288_),
    .B(_09279_),
    .C(_09278_),
    .Y(_09291_));
 sky130_fd_sc_hd__nand3_2 _30923_ (.A(_09012_),
    .B(_09002_),
    .C(_09014_),
    .Y(_09292_));
 sky130_vsdinv _30924_ (.A(_09292_),
    .Y(_09293_));
 sky130_fd_sc_hd__a21oi_2 _30925_ (.A1(_09290_),
    .A2(_09291_),
    .B1(_09293_),
    .Y(_09294_));
 sky130_fd_sc_hd__a21boi_2 _30926_ (.A1(_09278_),
    .A2(_09279_),
    .B1_N(_09289_),
    .Y(_09295_));
 sky130_fd_sc_hd__nor2_2 _30927_ (.A(_09289_),
    .B(_09280_),
    .Y(_09296_));
 sky130_fd_sc_hd__nor3_2 _30928_ (.A(_09292_),
    .B(_09295_),
    .C(_09296_),
    .Y(_09297_));
 sky130_fd_sc_hd__o21a_2 _30929_ (.A1(_08979_),
    .A2(_08980_),
    .B1(_08996_),
    .X(_09298_));
 sky130_fd_sc_hd__o21ai_2 _30930_ (.A1(_09294_),
    .A2(_09297_),
    .B1(_09298_),
    .Y(_09299_));
 sky130_fd_sc_hd__o21bai_2 _30931_ (.A1(_09295_),
    .A2(_09296_),
    .B1_N(_09293_),
    .Y(_09300_));
 sky130_fd_sc_hd__nand3_2 _30932_ (.A(_09290_),
    .B(_09291_),
    .C(_09293_),
    .Y(_09301_));
 sky130_fd_sc_hd__nand3b_2 _30933_ (.A_N(_09298_),
    .B(_09300_),
    .C(_09301_),
    .Y(_09302_));
 sky130_fd_sc_hd__buf_1 _30934_ (.A(_09005_),
    .X(_09303_));
 sky130_fd_sc_hd__nand2_2 _30935_ (.A(_09303_),
    .B(_05401_),
    .Y(_09304_));
 sky130_fd_sc_hd__buf_1 _30936_ (.A(\pcpi_mul.rs2[25] ),
    .X(_09305_));
 sky130_fd_sc_hd__nand2_2 _30937_ (.A(_09305_),
    .B(_19293_),
    .Y(_09306_));
 sky130_fd_sc_hd__nor2_2 _30938_ (.A(_09304_),
    .B(_09306_),
    .Y(_09307_));
 sky130_fd_sc_hd__buf_1 _30939_ (.A(\pcpi_mul.rs2[24] ),
    .X(_09308_));
 sky130_fd_sc_hd__and2_2 _30940_ (.A(_09308_),
    .B(_05444_),
    .X(_09309_));
 sky130_fd_sc_hd__nand2_2 _30941_ (.A(_09304_),
    .B(_09306_),
    .Y(_09310_));
 sky130_fd_sc_hd__nand3b_2 _30942_ (.A_N(_09307_),
    .B(_09309_),
    .C(_09310_),
    .Y(_09311_));
 sky130_fd_sc_hd__buf_1 _30943_ (.A(_09303_),
    .X(_09312_));
 sky130_fd_sc_hd__buf_1 _30944_ (.A(_08755_),
    .X(_09313_));
 sky130_fd_sc_hd__a22oi_2 _30945_ (.A1(_09312_),
    .A2(_05493_),
    .B1(_09313_),
    .B2(_05874_),
    .Y(_09314_));
 sky130_fd_sc_hd__o21bai_2 _30946_ (.A1(_09314_),
    .A2(_09307_),
    .B1_N(_09309_),
    .Y(_09315_));
 sky130_fd_sc_hd__a21oi_2 _30947_ (.A1(_09008_),
    .A2(_09013_),
    .B1(_09009_),
    .Y(_09316_));
 sky130_fd_sc_hd__a21bo_2 _30948_ (.A1(_09311_),
    .A2(_09315_),
    .B1_N(_09316_),
    .X(_09317_));
 sky130_fd_sc_hd__nand3b_2 _30949_ (.A_N(_09316_),
    .B(_09311_),
    .C(_09315_),
    .Y(_09318_));
 sky130_fd_sc_hd__buf_1 _30950_ (.A(_18722_),
    .X(_09319_));
 sky130_fd_sc_hd__buf_1 _30951_ (.A(_09319_),
    .X(_09320_));
 sky130_fd_sc_hd__buf_1 _30952_ (.A(_09320_),
    .X(_09321_));
 sky130_fd_sc_hd__and2_2 _30953_ (.A(_09321_),
    .B(_05466_),
    .X(_09322_));
 sky130_fd_sc_hd__a21oi_2 _30954_ (.A1(_09317_),
    .A2(_09318_),
    .B1(_09322_),
    .Y(_09323_));
 sky130_fd_sc_hd__nand3_2 _30955_ (.A(_09317_),
    .B(_09322_),
    .C(_09318_),
    .Y(_09324_));
 sky130_vsdinv _30956_ (.A(_09324_),
    .Y(_09325_));
 sky130_fd_sc_hd__nor2_2 _30957_ (.A(_09323_),
    .B(_09325_),
    .Y(_09326_));
 sky130_fd_sc_hd__a21oi_2 _30958_ (.A1(_09299_),
    .A2(_09302_),
    .B1(_09326_),
    .Y(_09327_));
 sky130_fd_sc_hd__nand3_2 _30959_ (.A(_09299_),
    .B(_09326_),
    .C(_09302_),
    .Y(_09328_));
 sky130_vsdinv _30960_ (.A(_09328_),
    .Y(_09329_));
 sky130_fd_sc_hd__o21bai_2 _30961_ (.A1(_09327_),
    .A2(_09329_),
    .B1_N(_09025_),
    .Y(_09330_));
 sky130_fd_sc_hd__o2bb2ai_2 _30962_ (.A1_N(_09302_),
    .A2_N(_09299_),
    .B1(_09325_),
    .B2(_09323_),
    .Y(_09331_));
 sky130_fd_sc_hd__buf_1 _30963_ (.A(_09328_),
    .X(_09332_));
 sky130_fd_sc_hd__nand3_2 _30964_ (.A(_09331_),
    .B(_09025_),
    .C(_09332_),
    .Y(_09333_));
 sky130_fd_sc_hd__nand2_2 _30965_ (.A(_07468_),
    .B(_05934_),
    .Y(_09334_));
 sky130_fd_sc_hd__nand2_2 _30966_ (.A(_07394_),
    .B(_06202_),
    .Y(_09335_));
 sky130_fd_sc_hd__nor2_2 _30967_ (.A(_09334_),
    .B(_09335_),
    .Y(_09336_));
 sky130_fd_sc_hd__and2_2 _30968_ (.A(_18790_),
    .B(_06477_),
    .X(_09337_));
 sky130_fd_sc_hd__nand2_2 _30969_ (.A(_09334_),
    .B(_09335_),
    .Y(_09338_));
 sky130_fd_sc_hd__nand3b_2 _30970_ (.A_N(_09336_),
    .B(_09337_),
    .C(_09338_),
    .Y(_09339_));
 sky130_fd_sc_hd__buf_1 _30971_ (.A(_05934_),
    .X(_09340_));
 sky130_fd_sc_hd__buf_1 _30972_ (.A(_19248_),
    .X(_09341_));
 sky130_fd_sc_hd__a22oi_2 _30973_ (.A1(_07469_),
    .A2(_09340_),
    .B1(_08908_),
    .B2(_09341_),
    .Y(_09342_));
 sky130_fd_sc_hd__o21bai_2 _30974_ (.A1(_09342_),
    .A2(_09336_),
    .B1_N(_09337_),
    .Y(_09343_));
 sky130_fd_sc_hd__nand2_2 _30975_ (.A(_09339_),
    .B(_09343_),
    .Y(_09344_));
 sky130_fd_sc_hd__a21oi_2 _30976_ (.A1(_08988_),
    .A2(_08991_),
    .B1(_08987_),
    .Y(_09345_));
 sky130_fd_sc_hd__nand2_2 _30977_ (.A(_09344_),
    .B(_09345_),
    .Y(_09346_));
 sky130_fd_sc_hd__nand3b_2 _30978_ (.A_N(_09345_),
    .B(_09339_),
    .C(_09343_),
    .Y(_09347_));
 sky130_fd_sc_hd__a21oi_2 _30979_ (.A1(_08910_),
    .A2(_08906_),
    .B1(_08904_),
    .Y(_09348_));
 sky130_vsdinv _30980_ (.A(_09348_),
    .Y(_09349_));
 sky130_fd_sc_hd__a21oi_2 _30981_ (.A1(_09346_),
    .A2(_09347_),
    .B1(_09349_),
    .Y(_09350_));
 sky130_fd_sc_hd__nand3_2 _30982_ (.A(_09346_),
    .B(_09349_),
    .C(_09347_),
    .Y(_09351_));
 sky130_vsdinv _30983_ (.A(_09351_),
    .Y(_09352_));
 sky130_fd_sc_hd__a21boi_2 _30984_ (.A1(_08915_),
    .A2(_08919_),
    .B1_N(_08916_),
    .Y(_09353_));
 sky130_fd_sc_hd__o21ai_2 _30985_ (.A1(_09350_),
    .A2(_09352_),
    .B1(_09353_),
    .Y(_09354_));
 sky130_fd_sc_hd__nand2_2 _30986_ (.A(_08922_),
    .B(_08916_),
    .Y(_09355_));
 sky130_fd_sc_hd__nand3b_2 _30987_ (.A_N(_09350_),
    .B(_09351_),
    .C(_09355_),
    .Y(_09356_));
 sky130_fd_sc_hd__nand2_2 _30988_ (.A(_09354_),
    .B(_09356_),
    .Y(_09357_));
 sky130_fd_sc_hd__nand2_2 _30989_ (.A(_06147_),
    .B(_19216_),
    .Y(_09358_));
 sky130_fd_sc_hd__nand2_2 _30990_ (.A(_06141_),
    .B(_08258_),
    .Y(_09359_));
 sky130_fd_sc_hd__nand2_2 _30991_ (.A(_09358_),
    .B(_09359_),
    .Y(_09360_));
 sky130_fd_sc_hd__nor2_2 _30992_ (.A(_09358_),
    .B(_09359_),
    .Y(_09361_));
 sky130_vsdinv _30993_ (.A(_09361_),
    .Y(_09362_));
 sky130_fd_sc_hd__o2bb2ai_2 _30994_ (.A1_N(_09360_),
    .A2_N(_09362_),
    .B1(_18824_),
    .B2(_19208_),
    .Y(_09363_));
 sky130_fd_sc_hd__buf_1 _30995_ (.A(_07324_),
    .X(_09364_));
 sky130_fd_sc_hd__and2_2 _30996_ (.A(_06137_),
    .B(_09364_),
    .X(_09365_));
 sky130_fd_sc_hd__nand3b_2 _30997_ (.A_N(_09361_),
    .B(_09365_),
    .C(_09360_),
    .Y(_09366_));
 sky130_fd_sc_hd__nand2_2 _30998_ (.A(_09363_),
    .B(_09366_),
    .Y(_09367_));
 sky130_fd_sc_hd__nand2_2 _30999_ (.A(_07495_),
    .B(_06466_),
    .Y(_09368_));
 sky130_fd_sc_hd__nand2_2 _31000_ (.A(_06540_),
    .B(_07304_),
    .Y(_09369_));
 sky130_fd_sc_hd__nor2_2 _31001_ (.A(_09368_),
    .B(_09369_),
    .Y(_09370_));
 sky130_fd_sc_hd__and2_2 _31002_ (.A(_18808_),
    .B(_06595_),
    .X(_09371_));
 sky130_fd_sc_hd__nand2_2 _31003_ (.A(_09368_),
    .B(_09369_),
    .Y(_09372_));
 sky130_fd_sc_hd__nand3b_2 _31004_ (.A_N(_09370_),
    .B(_09371_),
    .C(_09372_),
    .Y(_09373_));
 sky130_fd_sc_hd__a22oi_2 _31005_ (.A1(_08170_),
    .A2(_06351_),
    .B1(_18803_),
    .B2(_06454_),
    .Y(_09374_));
 sky130_fd_sc_hd__o21bai_2 _31006_ (.A1(_09374_),
    .A2(_09370_),
    .B1_N(_09371_),
    .Y(_09375_));
 sky130_fd_sc_hd__a21oi_2 _31007_ (.A1(_08934_),
    .A2(_08933_),
    .B1(_08932_),
    .Y(_09376_));
 sky130_fd_sc_hd__a21bo_2 _31008_ (.A1(_09373_),
    .A2(_09375_),
    .B1_N(_09376_),
    .X(_09377_));
 sky130_fd_sc_hd__nand3b_2 _31009_ (.A_N(_09376_),
    .B(_09373_),
    .C(_09375_),
    .Y(_09378_));
 sky130_fd_sc_hd__nand2_2 _31010_ (.A(_09377_),
    .B(_09378_),
    .Y(_09379_));
 sky130_fd_sc_hd__xnor2_2 _31011_ (.A(_09367_),
    .B(_09379_),
    .Y(_09380_));
 sky130_fd_sc_hd__nand2_2 _31012_ (.A(_09357_),
    .B(_09380_),
    .Y(_09381_));
 sky130_fd_sc_hd__xor2_2 _31013_ (.A(_09367_),
    .B(_09379_),
    .X(_09382_));
 sky130_fd_sc_hd__nand3_2 _31014_ (.A(_09382_),
    .B(_09354_),
    .C(_09356_),
    .Y(_09383_));
 sky130_vsdinv _31015_ (.A(_09001_),
    .Y(_09384_));
 sky130_fd_sc_hd__a21oi_2 _31016_ (.A1(_09381_),
    .A2(_09383_),
    .B1(_09384_),
    .Y(_09385_));
 sky130_fd_sc_hd__a21oi_2 _31017_ (.A1(_09354_),
    .A2(_09356_),
    .B1(_09382_),
    .Y(_09386_));
 sky130_fd_sc_hd__nor2_2 _31018_ (.A(_09380_),
    .B(_09357_),
    .Y(_09387_));
 sky130_fd_sc_hd__nor3_2 _31019_ (.A(_09001_),
    .B(_09386_),
    .C(_09387_),
    .Y(_09388_));
 sky130_fd_sc_hd__o21a_2 _31020_ (.A1(_08955_),
    .A2(_08961_),
    .B1(_08927_),
    .X(_09389_));
 sky130_vsdinv _31021_ (.A(_09389_),
    .Y(_09390_));
 sky130_fd_sc_hd__o21bai_2 _31022_ (.A1(_09385_),
    .A2(_09388_),
    .B1_N(_09390_),
    .Y(_09391_));
 sky130_fd_sc_hd__buf_1 _31023_ (.A(_09391_),
    .X(_09392_));
 sky130_fd_sc_hd__o21bai_2 _31024_ (.A1(_09386_),
    .A2(_09387_),
    .B1_N(_09384_),
    .Y(_09393_));
 sky130_fd_sc_hd__nand3_2 _31025_ (.A(_09381_),
    .B(_09384_),
    .C(_09383_),
    .Y(_09394_));
 sky130_fd_sc_hd__nand3_2 _31026_ (.A(_09393_),
    .B(_09390_),
    .C(_09394_),
    .Y(_09395_));
 sky130_fd_sc_hd__buf_1 _31027_ (.A(_09395_),
    .X(_09396_));
 sky130_fd_sc_hd__a22oi_2 _31028_ (.A1(_09330_),
    .A2(_09333_),
    .B1(_09392_),
    .B2(_09396_),
    .Y(_09397_));
 sky130_fd_sc_hd__nand2_2 _31029_ (.A(_09330_),
    .B(_09333_),
    .Y(_09398_));
 sky130_fd_sc_hd__nand2_2 _31030_ (.A(_09391_),
    .B(_09395_),
    .Y(_09399_));
 sky130_fd_sc_hd__nor2_2 _31031_ (.A(_09398_),
    .B(_09399_),
    .Y(_09400_));
 sky130_fd_sc_hd__nand2_2 _31032_ (.A(_09035_),
    .B(_09027_),
    .Y(_09401_));
 sky130_fd_sc_hd__o21bai_2 _31033_ (.A1(_09397_),
    .A2(_09400_),
    .B1_N(_09401_),
    .Y(_09402_));
 sky130_fd_sc_hd__a21oi_2 _31034_ (.A1(_09331_),
    .A2(_09332_),
    .B1(_09025_),
    .Y(_09403_));
 sky130_vsdinv _31035_ (.A(_09333_),
    .Y(_09404_));
 sky130_fd_sc_hd__nor2_2 _31036_ (.A(_09403_),
    .B(_09404_),
    .Y(_09405_));
 sky130_fd_sc_hd__nand3_2 _31037_ (.A(_09405_),
    .B(_09396_),
    .C(_09392_),
    .Y(_09406_));
 sky130_fd_sc_hd__nand2_2 _31038_ (.A(_09399_),
    .B(_09398_),
    .Y(_09407_));
 sky130_fd_sc_hd__nand3_2 _31039_ (.A(_09406_),
    .B(_09407_),
    .C(_09401_),
    .Y(_09408_));
 sky130_fd_sc_hd__buf_1 _31040_ (.A(_09408_),
    .X(_09409_));
 sky130_fd_sc_hd__a22oi_2 _31041_ (.A1(_09259_),
    .A2(_09262_),
    .B1(_09402_),
    .B2(_09409_),
    .Y(_09410_));
 sky130_fd_sc_hd__nand2_2 _31042_ (.A(_09259_),
    .B(_09262_),
    .Y(_09411_));
 sky130_fd_sc_hd__nand2_2 _31043_ (.A(_09402_),
    .B(_09408_),
    .Y(_09412_));
 sky130_fd_sc_hd__nor2_2 _31044_ (.A(_09411_),
    .B(_09412_),
    .Y(_09413_));
 sky130_fd_sc_hd__a31oi_2 _31045_ (.A1(_09127_),
    .A2(_09033_),
    .A3(_09130_),
    .B1(_09143_),
    .Y(_09414_));
 sky130_fd_sc_hd__o21ai_2 _31046_ (.A1(_09410_),
    .A2(_09413_),
    .B1(_09414_),
    .Y(_09415_));
 sky130_fd_sc_hd__a31o_2 _31047_ (.A1(_09127_),
    .A2(_09033_),
    .A3(_09129_),
    .B1(_09143_),
    .X(_09416_));
 sky130_fd_sc_hd__a21oi_2 _31048_ (.A1(_09252_),
    .A2(_09256_),
    .B1(_09260_),
    .Y(_09417_));
 sky130_vsdinv _31049_ (.A(_09261_),
    .Y(_09418_));
 sky130_fd_sc_hd__nor2_2 _31050_ (.A(_09417_),
    .B(_09418_),
    .Y(_09419_));
 sky130_fd_sc_hd__nand3_2 _31051_ (.A(_09419_),
    .B(_09409_),
    .C(_09402_),
    .Y(_09420_));
 sky130_fd_sc_hd__nand2_2 _31052_ (.A(_09412_),
    .B(_09411_),
    .Y(_09421_));
 sky130_fd_sc_hd__nand3_2 _31053_ (.A(_09416_),
    .B(_09420_),
    .C(_09421_),
    .Y(_09422_));
 sky130_fd_sc_hd__buf_1 _31054_ (.A(_09422_),
    .X(_09423_));
 sky130_fd_sc_hd__a21boi_2 _31055_ (.A1(_09102_),
    .A2(_09108_),
    .B1_N(_09103_),
    .Y(_09424_));
 sky130_fd_sc_hd__a21oi_2 _31056_ (.A1(_09130_),
    .A2(_09128_),
    .B1(_09424_),
    .Y(_09425_));
 sky130_fd_sc_hd__and3_2 _31057_ (.A(_09129_),
    .B(_09128_),
    .C(_09424_),
    .X(_09426_));
 sky130_fd_sc_hd__nor2_2 _31058_ (.A(_09425_),
    .B(_09426_),
    .Y(_09427_));
 sky130_fd_sc_hd__a21oi_2 _31059_ (.A1(_09415_),
    .A2(_09423_),
    .B1(_09427_),
    .Y(_09428_));
 sky130_fd_sc_hd__nand3_2 _31060_ (.A(_09415_),
    .B(_09427_),
    .C(_09422_),
    .Y(_09429_));
 sky130_vsdinv _31061_ (.A(_09429_),
    .Y(_09430_));
 sky130_fd_sc_hd__a21oi_2 _31062_ (.A1(_09145_),
    .A2(_09146_),
    .B1(_09138_),
    .Y(_09431_));
 sky130_fd_sc_hd__o21ai_2 _31063_ (.A1(_09151_),
    .A2(_09431_),
    .B1(_09147_),
    .Y(_09432_));
 sky130_fd_sc_hd__o21bai_2 _31064_ (.A1(_09428_),
    .A2(_09430_),
    .B1_N(_09432_),
    .Y(_09433_));
 sky130_fd_sc_hd__o2bb2ai_2 _31065_ (.A1_N(_09423_),
    .A2_N(_09415_),
    .B1(_09425_),
    .B2(_09426_),
    .Y(_09434_));
 sky130_fd_sc_hd__nand3_2 _31066_ (.A(_09434_),
    .B(_09432_),
    .C(_09429_),
    .Y(_09435_));
 sky130_fd_sc_hd__buf_1 _31067_ (.A(_09435_),
    .X(_09436_));
 sky130_fd_sc_hd__a21oi_2 _31068_ (.A1(_08863_),
    .A2(_08857_),
    .B1(_09149_),
    .Y(_09437_));
 sky130_fd_sc_hd__buf_1 _31069_ (.A(_09437_),
    .X(_09438_));
 sky130_fd_sc_hd__a21oi_2 _31070_ (.A1(_09433_),
    .A2(_09436_),
    .B1(_09438_),
    .Y(_09439_));
 sky130_fd_sc_hd__nand3_2 _31071_ (.A(_09433_),
    .B(_09438_),
    .C(_09435_),
    .Y(_09440_));
 sky130_vsdinv _31072_ (.A(_09440_),
    .Y(_09441_));
 sky130_vsdinv _31073_ (.A(_09159_),
    .Y(_09442_));
 sky130_fd_sc_hd__o21ai_2 _31074_ (.A1(_09442_),
    .A2(_09155_),
    .B1(_09162_),
    .Y(_09443_));
 sky130_fd_sc_hd__o21bai_2 _31075_ (.A1(_09439_),
    .A2(_09441_),
    .B1_N(_09443_),
    .Y(_09444_));
 sky130_fd_sc_hd__a21oi_2 _31076_ (.A1(_09434_),
    .A2(_09429_),
    .B1(_09432_),
    .Y(_09445_));
 sky130_vsdinv _31077_ (.A(_09436_),
    .Y(_09446_));
 sky130_fd_sc_hd__o21bai_2 _31078_ (.A1(_09445_),
    .A2(_09446_),
    .B1_N(_09438_),
    .Y(_09447_));
 sky130_fd_sc_hd__nand3_2 _31079_ (.A(_09447_),
    .B(_09440_),
    .C(_09443_),
    .Y(_09448_));
 sky130_fd_sc_hd__nand2_2 _31080_ (.A(_09444_),
    .B(_09448_),
    .Y(_09449_));
 sky130_fd_sc_hd__a21oi_2 _31081_ (.A1(_09161_),
    .A2(_09162_),
    .B1(_09159_),
    .Y(_09450_));
 sky130_fd_sc_hd__nor3_2 _31082_ (.A(_09442_),
    .B(_09155_),
    .C(_09158_),
    .Y(_09451_));
 sky130_fd_sc_hd__o21bai_2 _31083_ (.A1(_09450_),
    .A2(_09451_),
    .B1_N(_09164_),
    .Y(_09452_));
 sky130_fd_sc_hd__a21oi_2 _31084_ (.A1(_09172_),
    .A2(_09452_),
    .B1(_09167_),
    .Y(_09453_));
 sky130_fd_sc_hd__xor2_2 _31085_ (.A(_09449_),
    .B(_09453_),
    .X(_02646_));
 sky130_fd_sc_hd__a22oi_2 _31086_ (.A1(_06105_),
    .A2(_07961_),
    .B1(_06230_),
    .B2(_07963_),
    .Y(_09454_));
 sky130_fd_sc_hd__nand2_2 _31087_ (.A(_05869_),
    .B(_07745_),
    .Y(_09455_));
 sky130_fd_sc_hd__buf_1 _31088_ (.A(_08569_),
    .X(_09456_));
 sky130_fd_sc_hd__nand2_2 _31089_ (.A(_06889_),
    .B(_09456_),
    .Y(_09457_));
 sky130_fd_sc_hd__nor2_2 _31090_ (.A(_09455_),
    .B(_09457_),
    .Y(_09458_));
 sky130_fd_sc_hd__and2_2 _31091_ (.A(_05586_),
    .B(_07951_),
    .X(_09459_));
 sky130_fd_sc_hd__o21bai_2 _31092_ (.A1(_09454_),
    .A2(_09458_),
    .B1_N(_09459_),
    .Y(_09460_));
 sky130_fd_sc_hd__nand3b_2 _31093_ (.A_N(_09455_),
    .B(_06237_),
    .C(_08310_),
    .Y(_09461_));
 sky130_fd_sc_hd__nand2_2 _31094_ (.A(_09455_),
    .B(_09457_),
    .Y(_09462_));
 sky130_fd_sc_hd__nand3_2 _31095_ (.A(_09461_),
    .B(_09459_),
    .C(_09462_),
    .Y(_09463_));
 sky130_fd_sc_hd__nand2_2 _31096_ (.A(_09460_),
    .B(_09463_),
    .Y(_09464_));
 sky130_fd_sc_hd__a21oi_2 _31097_ (.A1(_09360_),
    .A2(_09365_),
    .B1(_09361_),
    .Y(_09465_));
 sky130_fd_sc_hd__nand2_2 _31098_ (.A(_09464_),
    .B(_09465_),
    .Y(_09466_));
 sky130_fd_sc_hd__nand3b_2 _31099_ (.A_N(_09465_),
    .B(_09463_),
    .C(_09460_),
    .Y(_09467_));
 sky130_fd_sc_hd__a21oi_2 _31100_ (.A1(_09180_),
    .A2(_09177_),
    .B1(_09176_),
    .Y(_09468_));
 sky130_vsdinv _31101_ (.A(_09468_),
    .Y(_09469_));
 sky130_fd_sc_hd__a21oi_2 _31102_ (.A1(_09466_),
    .A2(_09467_),
    .B1(_09469_),
    .Y(_09470_));
 sky130_fd_sc_hd__nand3_2 _31103_ (.A(_09466_),
    .B(_09469_),
    .C(_09467_),
    .Y(_09471_));
 sky130_vsdinv _31104_ (.A(_09471_),
    .Y(_09472_));
 sky130_fd_sc_hd__a21boi_2 _31105_ (.A1(_09373_),
    .A2(_09375_),
    .B1_N(_09376_),
    .Y(_09473_));
 sky130_fd_sc_hd__o21a_2 _31106_ (.A1(_09367_),
    .A2(_09473_),
    .B1(_09378_),
    .X(_09474_));
 sky130_fd_sc_hd__o21ai_2 _31107_ (.A1(_09470_),
    .A2(_09472_),
    .B1(_09474_),
    .Y(_09475_));
 sky130_fd_sc_hd__a21o_2 _31108_ (.A1(_09466_),
    .A2(_09467_),
    .B1(_09469_),
    .X(_09476_));
 sky130_fd_sc_hd__o21ai_2 _31109_ (.A1(_09367_),
    .A2(_09473_),
    .B1(_09378_),
    .Y(_09477_));
 sky130_fd_sc_hd__nand3_2 _31110_ (.A(_09476_),
    .B(_09477_),
    .C(_09471_),
    .Y(_09478_));
 sky130_vsdinv _31111_ (.A(_09186_),
    .Y(_09479_));
 sky130_fd_sc_hd__a21oi_2 _31112_ (.A1(_09185_),
    .A2(_09188_),
    .B1(_09479_),
    .Y(_09480_));
 sky130_vsdinv _31113_ (.A(_09480_),
    .Y(_09481_));
 sky130_fd_sc_hd__a21oi_2 _31114_ (.A1(_09475_),
    .A2(_09478_),
    .B1(_09481_),
    .Y(_09482_));
 sky130_fd_sc_hd__nand3_2 _31115_ (.A(_09475_),
    .B(_09481_),
    .C(_09478_),
    .Y(_09483_));
 sky130_vsdinv _31116_ (.A(_09483_),
    .Y(_09484_));
 sky130_fd_sc_hd__a21oi_2 _31117_ (.A1(_09194_),
    .A2(_09190_),
    .B1(_09195_),
    .Y(_09485_));
 sky130_fd_sc_hd__o21ai_2 _31118_ (.A1(_09197_),
    .A2(_09485_),
    .B1(_09196_),
    .Y(_09486_));
 sky130_fd_sc_hd__o21bai_2 _31119_ (.A1(_09482_),
    .A2(_09484_),
    .B1_N(_09486_),
    .Y(_09487_));
 sky130_fd_sc_hd__nand2_2 _31120_ (.A(_09475_),
    .B(_09478_),
    .Y(_09488_));
 sky130_fd_sc_hd__nand2_2 _31121_ (.A(_09488_),
    .B(_09480_),
    .Y(_09489_));
 sky130_fd_sc_hd__nand3_2 _31122_ (.A(_09489_),
    .B(_09486_),
    .C(_09483_),
    .Y(_09490_));
 sky130_fd_sc_hd__buf_1 _31123_ (.A(_09490_),
    .X(_09491_));
 sky130_fd_sc_hd__buf_1 _31124_ (.A(_19179_),
    .X(_09492_));
 sky130_fd_sc_hd__buf_1 _31125_ (.A(_19171_),
    .X(_09493_));
 sky130_fd_sc_hd__a22o_2 _31126_ (.A1(_05813_),
    .A2(_09492_),
    .B1(_05816_),
    .B2(_09493_),
    .X(_09494_));
 sky130_fd_sc_hd__buf_1 _31127_ (.A(\pcpi_mul.rs1[23] ),
    .X(_09495_));
 sky130_fd_sc_hd__nand2_2 _31128_ (.A(_05724_),
    .B(_09495_),
    .Y(_09496_));
 sky130_fd_sc_hd__buf_1 _31129_ (.A(_08556_),
    .X(_09497_));
 sky130_fd_sc_hd__nand3b_2 _31130_ (.A_N(_09496_),
    .B(_05638_),
    .C(_09497_),
    .Y(_09498_));
 sky130_fd_sc_hd__o2bb2ai_2 _31131_ (.A1_N(_09494_),
    .A2_N(_09498_),
    .B1(_06346_),
    .B2(_19150_),
    .Y(_09499_));
 sky130_fd_sc_hd__buf_1 _31132_ (.A(\pcpi_mul.rs1[28] ),
    .X(_09500_));
 sky130_fd_sc_hd__and2_2 _31133_ (.A(_05820_),
    .B(_09500_),
    .X(_09501_));
 sky130_fd_sc_hd__nand3_2 _31134_ (.A(_09498_),
    .B(_09494_),
    .C(_09501_),
    .Y(_09502_));
 sky130_fd_sc_hd__a21oi_2 _31135_ (.A1(_09214_),
    .A2(_09213_),
    .B1(_09211_),
    .Y(_09503_));
 sky130_vsdinv _31136_ (.A(_09503_),
    .Y(_09504_));
 sky130_fd_sc_hd__a21o_2 _31137_ (.A1(_09499_),
    .A2(_09502_),
    .B1(_09504_),
    .X(_09505_));
 sky130_fd_sc_hd__nand3_2 _31138_ (.A(_09499_),
    .B(_09504_),
    .C(_09502_),
    .Y(_09506_));
 sky130_fd_sc_hd__buf_1 _31139_ (.A(_09506_),
    .X(_09507_));
 sky130_fd_sc_hd__nand2_2 _31140_ (.A(_18865_),
    .B(_09224_),
    .Y(_09508_));
 sky130_fd_sc_hd__nand2_2 _31141_ (.A(_05427_),
    .B(_09212_),
    .Y(_09509_));
 sky130_fd_sc_hd__xor2_2 _31142_ (.A(_09508_),
    .B(_09509_),
    .X(_09510_));
 sky130_fd_sc_hd__buf_1 _31143_ (.A(\pcpi_mul.rs1[25] ),
    .X(_09511_));
 sky130_fd_sc_hd__and2_2 _31144_ (.A(_05437_),
    .B(_09511_),
    .X(_09512_));
 sky130_fd_sc_hd__nand2_2 _31145_ (.A(_09510_),
    .B(_09512_),
    .Y(_09513_));
 sky130_fd_sc_hd__xnor2_2 _31146_ (.A(_09508_),
    .B(_09509_),
    .Y(_09514_));
 sky130_fd_sc_hd__o21ai_2 _31147_ (.A1(_18855_),
    .A2(_19168_),
    .B1(_09514_),
    .Y(_09515_));
 sky130_fd_sc_hd__nand2_2 _31148_ (.A(_09513_),
    .B(_09515_),
    .Y(_09516_));
 sky130_fd_sc_hd__buf_1 _31149_ (.A(_09516_),
    .X(_09517_));
 sky130_fd_sc_hd__a21boi_2 _31150_ (.A1(_09505_),
    .A2(_09507_),
    .B1_N(_09517_),
    .Y(_09518_));
 sky130_fd_sc_hd__a21oi_2 _31151_ (.A1(_09499_),
    .A2(_09502_),
    .B1(_09504_),
    .Y(_09519_));
 sky130_fd_sc_hd__nor3b_2 _31152_ (.A(_09517_),
    .B(_09519_),
    .C_N(_09506_),
    .Y(_09520_));
 sky130_fd_sc_hd__a21boi_2 _31153_ (.A1(_09215_),
    .A2(_09218_),
    .B1_N(_09219_),
    .Y(_09521_));
 sky130_fd_sc_hd__o21ai_2 _31154_ (.A1(_09521_),
    .A2(_09231_),
    .B1(_09221_),
    .Y(_09522_));
 sky130_fd_sc_hd__o21bai_2 _31155_ (.A1(_09518_),
    .A2(_09520_),
    .B1_N(_09522_),
    .Y(_09523_));
 sky130_vsdinv _31156_ (.A(_09516_),
    .Y(_09524_));
 sky130_fd_sc_hd__a21o_2 _31157_ (.A1(_09505_),
    .A2(_09507_),
    .B1(_09524_),
    .X(_09525_));
 sky130_fd_sc_hd__nand3b_2 _31158_ (.A_N(_09517_),
    .B(_09505_),
    .C(_09507_),
    .Y(_09526_));
 sky130_fd_sc_hd__nand3_2 _31159_ (.A(_09525_),
    .B(_09526_),
    .C(_09522_),
    .Y(_09527_));
 sky130_fd_sc_hd__nand2_2 _31160_ (.A(_09523_),
    .B(_09527_),
    .Y(_09528_));
 sky130_fd_sc_hd__o21a_2 _31161_ (.A1(_09223_),
    .A2(_09225_),
    .B1(_09228_),
    .X(_09529_));
 sky130_fd_sc_hd__nand2_2 _31162_ (.A(_09528_),
    .B(_09529_),
    .Y(_09530_));
 sky130_fd_sc_hd__nand3b_2 _31163_ (.A_N(_09529_),
    .B(_09523_),
    .C(_09527_),
    .Y(_09531_));
 sky130_fd_sc_hd__nand2_2 _31164_ (.A(_09530_),
    .B(_09531_),
    .Y(_09532_));
 sky130_fd_sc_hd__buf_1 _31165_ (.A(_09532_),
    .X(_09533_));
 sky130_fd_sc_hd__a21boi_2 _31166_ (.A1(_09487_),
    .A2(_09491_),
    .B1_N(_09533_),
    .Y(_09534_));
 sky130_fd_sc_hd__a21oi_2 _31167_ (.A1(_09489_),
    .A2(_09483_),
    .B1(_09486_),
    .Y(_09535_));
 sky130_fd_sc_hd__nor3b_2 _31168_ (.A(_09533_),
    .B(_09535_),
    .C_N(_09491_),
    .Y(_09536_));
 sky130_fd_sc_hd__o21ai_2 _31169_ (.A1(_09389_),
    .A2(_09385_),
    .B1(_09394_),
    .Y(_09537_));
 sky130_fd_sc_hd__o21bai_2 _31170_ (.A1(_09534_),
    .A2(_09536_),
    .B1_N(_09537_),
    .Y(_09538_));
 sky130_fd_sc_hd__a21bo_2 _31171_ (.A1(_09490_),
    .A2(_09487_),
    .B1_N(_09533_),
    .X(_09539_));
 sky130_fd_sc_hd__nand3b_2 _31172_ (.A_N(_09532_),
    .B(_09491_),
    .C(_09487_),
    .Y(_09540_));
 sky130_fd_sc_hd__nand3_2 _31173_ (.A(_09539_),
    .B(_09537_),
    .C(_09540_),
    .Y(_09541_));
 sky130_fd_sc_hd__nand2_2 _31174_ (.A(_09538_),
    .B(_09541_),
    .Y(_09542_));
 sky130_fd_sc_hd__o21a_2 _31175_ (.A1(_09248_),
    .A2(_09249_),
    .B1(_09208_),
    .X(_09543_));
 sky130_fd_sc_hd__nand2_2 _31176_ (.A(_09542_),
    .B(_09543_),
    .Y(_09544_));
 sky130_fd_sc_hd__buf_1 _31177_ (.A(_09541_),
    .X(_09545_));
 sky130_fd_sc_hd__nand3b_2 _31178_ (.A_N(_09543_),
    .B(_09538_),
    .C(_09545_),
    .Y(_09546_));
 sky130_fd_sc_hd__buf_1 _31179_ (.A(_09546_),
    .X(_09547_));
 sky130_fd_sc_hd__buf_1 _31180_ (.A(_18752_),
    .X(_09548_));
 sky130_fd_sc_hd__a22oi_2 _31181_ (.A1(_08226_),
    .A2(_05536_),
    .B1(_09548_),
    .B2(_05851_),
    .Y(_09549_));
 sky130_fd_sc_hd__nand2_2 _31182_ (.A(_08471_),
    .B(_05517_),
    .Y(_09550_));
 sky130_fd_sc_hd__nand2_2 _31183_ (.A(_09266_),
    .B(_05500_),
    .Y(_09551_));
 sky130_fd_sc_hd__nor2_2 _31184_ (.A(_09550_),
    .B(_09551_),
    .Y(_09552_));
 sky130_fd_sc_hd__nand2_2 _31185_ (.A(_07844_),
    .B(_05837_),
    .Y(_09553_));
 sky130_vsdinv _31186_ (.A(_09553_),
    .Y(_09554_));
 sky130_fd_sc_hd__o21bai_2 _31187_ (.A1(_09549_),
    .A2(_09552_),
    .B1_N(_09554_),
    .Y(_09555_));
 sky130_fd_sc_hd__nand3b_2 _31188_ (.A_N(_09550_),
    .B(_09272_),
    .C(_06041_),
    .Y(_09556_));
 sky130_fd_sc_hd__nand2_2 _31189_ (.A(_09550_),
    .B(_09551_),
    .Y(_09557_));
 sky130_fd_sc_hd__nand3_2 _31190_ (.A(_09556_),
    .B(_09554_),
    .C(_09557_),
    .Y(_09558_));
 sky130_fd_sc_hd__nand2_2 _31191_ (.A(_09555_),
    .B(_09558_),
    .Y(_09559_));
 sky130_fd_sc_hd__o21ai_2 _31192_ (.A1(_09269_),
    .A2(_09264_),
    .B1(_09273_),
    .Y(_09560_));
 sky130_vsdinv _31193_ (.A(_09560_),
    .Y(_09561_));
 sky130_fd_sc_hd__nand2_2 _31194_ (.A(_09559_),
    .B(_09561_),
    .Y(_09562_));
 sky130_fd_sc_hd__nand3_2 _31195_ (.A(_09555_),
    .B(_09558_),
    .C(_09560_),
    .Y(_09563_));
 sky130_fd_sc_hd__buf_1 _31196_ (.A(_09563_),
    .X(_09564_));
 sky130_fd_sc_hd__nand2_2 _31197_ (.A(_18763_),
    .B(_05727_),
    .Y(_09565_));
 sky130_fd_sc_hd__nand2_2 _31198_ (.A(_18769_),
    .B(_05957_),
    .Y(_09566_));
 sky130_fd_sc_hd__nor2_2 _31199_ (.A(_09565_),
    .B(_09566_),
    .Y(_09567_));
 sky130_fd_sc_hd__nand2_2 _31200_ (.A(_09565_),
    .B(_09566_),
    .Y(_09568_));
 sky130_vsdinv _31201_ (.A(_09568_),
    .Y(_09569_));
 sky130_fd_sc_hd__and2_2 _31202_ (.A(\pcpi_mul.rs2[18] ),
    .B(_06067_),
    .X(_09570_));
 sky130_fd_sc_hd__o21bai_2 _31203_ (.A1(_09567_),
    .A2(_09569_),
    .B1_N(_09570_),
    .Y(_09571_));
 sky130_fd_sc_hd__nand3b_2 _31204_ (.A_N(_09567_),
    .B(_09570_),
    .C(_09568_),
    .Y(_09572_));
 sky130_fd_sc_hd__nand2_2 _31205_ (.A(_09571_),
    .B(_09572_),
    .Y(_09573_));
 sky130_fd_sc_hd__buf_1 _31206_ (.A(_09573_),
    .X(_09574_));
 sky130_fd_sc_hd__a21boi_2 _31207_ (.A1(_09562_),
    .A2(_09564_),
    .B1_N(_09574_),
    .Y(_09575_));
 sky130_fd_sc_hd__a21oi_2 _31208_ (.A1(_09555_),
    .A2(_09558_),
    .B1(_09560_),
    .Y(_09576_));
 sky130_fd_sc_hd__nor3b_2 _31209_ (.A(_09574_),
    .B(_09576_),
    .C_N(_09564_),
    .Y(_09577_));
 sky130_vsdinv _31210_ (.A(_09318_),
    .Y(_09578_));
 sky130_fd_sc_hd__o21bai_2 _31211_ (.A1(_09575_),
    .A2(_09577_),
    .B1_N(_09578_),
    .Y(_09579_));
 sky130_fd_sc_hd__a21bo_2 _31212_ (.A1(_09562_),
    .A2(_09563_),
    .B1_N(_09574_),
    .X(_09580_));
 sky130_fd_sc_hd__nand3b_2 _31213_ (.A_N(_09573_),
    .B(_09562_),
    .C(_09564_),
    .Y(_09581_));
 sky130_fd_sc_hd__nand3_2 _31214_ (.A(_09580_),
    .B(_09578_),
    .C(_09581_),
    .Y(_09582_));
 sky130_fd_sc_hd__nand2_2 _31215_ (.A(_09579_),
    .B(_09582_),
    .Y(_09583_));
 sky130_fd_sc_hd__o21a_2 _31216_ (.A1(_09289_),
    .A2(_09280_),
    .B1(_09279_),
    .X(_09584_));
 sky130_fd_sc_hd__nand2_2 _31217_ (.A(_09583_),
    .B(_09584_),
    .Y(_09585_));
 sky130_fd_sc_hd__nand3b_2 _31218_ (.A_N(_09584_),
    .B(_09579_),
    .C(_09582_),
    .Y(_09586_));
 sky130_fd_sc_hd__buf_1 _31219_ (.A(\pcpi_mul.rs2[26] ),
    .X(_09587_));
 sky130_fd_sc_hd__nand2_2 _31220_ (.A(_09587_),
    .B(_05430_),
    .Y(_09588_));
 sky130_fd_sc_hd__buf_1 _31221_ (.A(\pcpi_mul.rs2[25] ),
    .X(_09589_));
 sky130_fd_sc_hd__nand2_2 _31222_ (.A(_09589_),
    .B(_05986_),
    .Y(_09590_));
 sky130_fd_sc_hd__nor2_2 _31223_ (.A(_09588_),
    .B(_09590_),
    .Y(_09591_));
 sky130_fd_sc_hd__nand2_2 _31224_ (.A(_09588_),
    .B(_09590_),
    .Y(_09592_));
 sky130_vsdinv _31225_ (.A(_09592_),
    .Y(_09593_));
 sky130_fd_sc_hd__and2_2 _31226_ (.A(_09308_),
    .B(_05674_),
    .X(_09594_));
 sky130_fd_sc_hd__o21bai_2 _31227_ (.A1(_09591_),
    .A2(_09593_),
    .B1_N(_09594_),
    .Y(_09595_));
 sky130_fd_sc_hd__nand3b_2 _31228_ (.A_N(_09591_),
    .B(_09594_),
    .C(_09592_),
    .Y(_09596_));
 sky130_fd_sc_hd__a21oi_2 _31229_ (.A1(_09310_),
    .A2(_09309_),
    .B1(_09307_),
    .Y(_09597_));
 sky130_vsdinv _31230_ (.A(_09597_),
    .Y(_09598_));
 sky130_fd_sc_hd__a21o_2 _31231_ (.A1(_09595_),
    .A2(_09596_),
    .B1(_09598_),
    .X(_09599_));
 sky130_fd_sc_hd__nand3_2 _31232_ (.A(_09598_),
    .B(_09595_),
    .C(_09596_),
    .Y(_09600_));
 sky130_fd_sc_hd__buf_1 _31233_ (.A(_09600_),
    .X(_09601_));
 sky130_fd_sc_hd__nand2_2 _31234_ (.A(_09599_),
    .B(_09601_),
    .Y(_09602_));
 sky130_fd_sc_hd__buf_1 _31235_ (.A(_18716_),
    .X(_09603_));
 sky130_fd_sc_hd__nand2_2 _31236_ (.A(_09603_),
    .B(_19301_),
    .Y(_09604_));
 sky130_fd_sc_hd__buf_1 _31237_ (.A(\pcpi_mul.rs2[27] ),
    .X(_09605_));
 sky130_fd_sc_hd__buf_1 _31238_ (.A(_09605_),
    .X(_09606_));
 sky130_fd_sc_hd__nand2_2 _31239_ (.A(_09606_),
    .B(_06143_),
    .Y(_09607_));
 sky130_fd_sc_hd__xor2_2 _31240_ (.A(_09604_),
    .B(_09607_),
    .X(_09608_));
 sky130_vsdinv _31241_ (.A(_09608_),
    .Y(_09609_));
 sky130_fd_sc_hd__nand2_2 _31242_ (.A(_09602_),
    .B(_09609_),
    .Y(_09610_));
 sky130_fd_sc_hd__nand3_2 _31243_ (.A(_09599_),
    .B(_09608_),
    .C(_09600_),
    .Y(_09611_));
 sky130_fd_sc_hd__a21oi_2 _31244_ (.A1(_09610_),
    .A2(_09611_),
    .B1(_09325_),
    .Y(_09612_));
 sky130_fd_sc_hd__a21oi_2 _31245_ (.A1(_09599_),
    .A2(_09601_),
    .B1(_09608_),
    .Y(_09613_));
 sky130_vsdinv _31246_ (.A(_09611_),
    .Y(_09614_));
 sky130_fd_sc_hd__nor3_2 _31247_ (.A(_09324_),
    .B(_09613_),
    .C(_09614_),
    .Y(_09615_));
 sky130_fd_sc_hd__nor2_2 _31248_ (.A(_09612_),
    .B(_09615_),
    .Y(_09616_));
 sky130_fd_sc_hd__a21oi_2 _31249_ (.A1(_09585_),
    .A2(_09586_),
    .B1(_09616_),
    .Y(_09617_));
 sky130_fd_sc_hd__o21ai_2 _31250_ (.A1(_09613_),
    .A2(_09614_),
    .B1(_09324_),
    .Y(_09618_));
 sky130_fd_sc_hd__nand3_2 _31251_ (.A(_09325_),
    .B(_09610_),
    .C(_09611_),
    .Y(_09619_));
 sky130_fd_sc_hd__nand2_2 _31252_ (.A(_09618_),
    .B(_09619_),
    .Y(_09620_));
 sky130_fd_sc_hd__a21boi_2 _31253_ (.A1(_09579_),
    .A2(_09582_),
    .B1_N(_09584_),
    .Y(_09621_));
 sky130_fd_sc_hd__nor3b_2 _31254_ (.A(_09620_),
    .B(_09621_),
    .C_N(_09586_),
    .Y(_09622_));
 sky130_fd_sc_hd__o21ai_2 _31255_ (.A1(_09617_),
    .A2(_09622_),
    .B1(_09332_),
    .Y(_09623_));
 sky130_fd_sc_hd__o2bb2ai_2 _31256_ (.A1_N(_09586_),
    .A2_N(_09585_),
    .B1(_09615_),
    .B2(_09612_),
    .Y(_09624_));
 sky130_fd_sc_hd__nand3_2 _31257_ (.A(_09585_),
    .B(_09616_),
    .C(_09586_),
    .Y(_09625_));
 sky130_fd_sc_hd__nand3_2 _31258_ (.A(_09329_),
    .B(_09624_),
    .C(_09625_),
    .Y(_09626_));
 sky130_fd_sc_hd__nand2_2 _31259_ (.A(_07785_),
    .B(_19248_),
    .Y(_09627_));
 sky130_fd_sc_hd__nand2_2 _31260_ (.A(_07787_),
    .B(_06364_),
    .Y(_09628_));
 sky130_fd_sc_hd__nor2_2 _31261_ (.A(_09627_),
    .B(_09628_),
    .Y(_09629_));
 sky130_fd_sc_hd__and2_2 _31262_ (.A(_06665_),
    .B(_07690_),
    .X(_09630_));
 sky130_fd_sc_hd__nand2_2 _31263_ (.A(_09627_),
    .B(_09628_),
    .Y(_09631_));
 sky130_fd_sc_hd__nand3b_2 _31264_ (.A_N(_09629_),
    .B(_09630_),
    .C(_09631_),
    .Y(_09632_));
 sky130_fd_sc_hd__a22oi_2 _31265_ (.A1(_07786_),
    .A2(_07060_),
    .B1(_07788_),
    .B2(_06463_),
    .Y(_09633_));
 sky130_fd_sc_hd__o21bai_2 _31266_ (.A1(_09633_),
    .A2(_09629_),
    .B1_N(_09630_),
    .Y(_09634_));
 sky130_fd_sc_hd__nand2_2 _31267_ (.A(_09632_),
    .B(_09634_),
    .Y(_09635_));
 sky130_fd_sc_hd__nor2_2 _31268_ (.A(_09281_),
    .B(_09282_),
    .Y(_09636_));
 sky130_fd_sc_hd__a21oi_2 _31269_ (.A1(_09283_),
    .A2(_09286_),
    .B1(_09636_),
    .Y(_09637_));
 sky130_fd_sc_hd__nand2_2 _31270_ (.A(_09635_),
    .B(_09637_),
    .Y(_09638_));
 sky130_fd_sc_hd__nand3b_2 _31271_ (.A_N(_09637_),
    .B(_09632_),
    .C(_09634_),
    .Y(_09639_));
 sky130_fd_sc_hd__nand2_2 _31272_ (.A(_09638_),
    .B(_09639_),
    .Y(_09640_));
 sky130_fd_sc_hd__a21oi_2 _31273_ (.A1(_09338_),
    .A2(_09337_),
    .B1(_09336_),
    .Y(_09641_));
 sky130_fd_sc_hd__nand2_2 _31274_ (.A(_09640_),
    .B(_09641_),
    .Y(_09642_));
 sky130_fd_sc_hd__nand3b_2 _31275_ (.A_N(_09641_),
    .B(_09638_),
    .C(_09639_),
    .Y(_09643_));
 sky130_fd_sc_hd__nand2_2 _31276_ (.A(_09642_),
    .B(_09643_),
    .Y(_09644_));
 sky130_fd_sc_hd__a21boi_2 _31277_ (.A1(_09346_),
    .A2(_09349_),
    .B1_N(_09347_),
    .Y(_09645_));
 sky130_fd_sc_hd__nand2_2 _31278_ (.A(_09644_),
    .B(_09645_),
    .Y(_09646_));
 sky130_fd_sc_hd__nand2_2 _31279_ (.A(_09351_),
    .B(_09347_),
    .Y(_09647_));
 sky130_fd_sc_hd__nand3_2 _31280_ (.A(_09647_),
    .B(_09642_),
    .C(_09643_),
    .Y(_09648_));
 sky130_fd_sc_hd__nand2_2 _31281_ (.A(_09646_),
    .B(_09648_),
    .Y(_09649_));
 sky130_fd_sc_hd__nand2_2 _31282_ (.A(_18797_),
    .B(_06606_),
    .Y(_09650_));
 sky130_fd_sc_hd__nand2_2 _31283_ (.A(_07192_),
    .B(_07694_),
    .Y(_09651_));
 sky130_fd_sc_hd__nor2_2 _31284_ (.A(_09650_),
    .B(_09651_),
    .Y(_09652_));
 sky130_fd_sc_hd__and2_2 _31285_ (.A(_08038_),
    .B(_06734_),
    .X(_09653_));
 sky130_fd_sc_hd__nand2_2 _31286_ (.A(_09650_),
    .B(_09651_),
    .Y(_09654_));
 sky130_fd_sc_hd__nand3b_2 _31287_ (.A_N(_09652_),
    .B(_09653_),
    .C(_09654_),
    .Y(_09655_));
 sky130_fd_sc_hd__a22oi_2 _31288_ (.A1(_07199_),
    .A2(_07699_),
    .B1(_07201_),
    .B2(_07906_),
    .Y(_09656_));
 sky130_fd_sc_hd__o21bai_2 _31289_ (.A1(_09656_),
    .A2(_09652_),
    .B1_N(_09653_),
    .Y(_09657_));
 sky130_fd_sc_hd__a21oi_2 _31290_ (.A1(_09372_),
    .A2(_09371_),
    .B1(_09370_),
    .Y(_09658_));
 sky130_fd_sc_hd__a21boi_2 _31291_ (.A1(_09655_),
    .A2(_09657_),
    .B1_N(_09658_),
    .Y(_09659_));
 sky130_fd_sc_hd__nand2_2 _31292_ (.A(_06670_),
    .B(_07605_),
    .Y(_09660_));
 sky130_fd_sc_hd__nand2_2 _31293_ (.A(_06673_),
    .B(_07325_),
    .Y(_09661_));
 sky130_fd_sc_hd__nand2_2 _31294_ (.A(_09660_),
    .B(_09661_),
    .Y(_09662_));
 sky130_fd_sc_hd__nor2_2 _31295_ (.A(_09660_),
    .B(_09661_),
    .Y(_09663_));
 sky130_vsdinv _31296_ (.A(_09663_),
    .Y(_09664_));
 sky130_fd_sc_hd__buf_1 _31297_ (.A(_19204_),
    .X(_09665_));
 sky130_fd_sc_hd__o2bb2ai_2 _31298_ (.A1_N(_09662_),
    .A2_N(_09664_),
    .B1(_18824_),
    .B2(_09665_),
    .Y(_09666_));
 sky130_fd_sc_hd__and2_2 _31299_ (.A(_05895_),
    .B(_08292_),
    .X(_09667_));
 sky130_fd_sc_hd__nand3b_2 _31300_ (.A_N(_09663_),
    .B(_09667_),
    .C(_09662_),
    .Y(_09668_));
 sky130_fd_sc_hd__nand2_2 _31301_ (.A(_09666_),
    .B(_09668_),
    .Y(_09669_));
 sky130_vsdinv _31302_ (.A(_09669_),
    .Y(_09670_));
 sky130_fd_sc_hd__nand3b_2 _31303_ (.A_N(_09658_),
    .B(_09655_),
    .C(_09657_),
    .Y(_09671_));
 sky130_fd_sc_hd__nand3b_2 _31304_ (.A_N(_09659_),
    .B(_09670_),
    .C(_09671_),
    .Y(_09672_));
 sky130_vsdinv _31305_ (.A(_09671_),
    .Y(_09673_));
 sky130_fd_sc_hd__o21ai_2 _31306_ (.A1(_09659_),
    .A2(_09673_),
    .B1(_09669_),
    .Y(_09674_));
 sky130_fd_sc_hd__nand2_2 _31307_ (.A(_09672_),
    .B(_09674_),
    .Y(_09675_));
 sky130_fd_sc_hd__nand2_2 _31308_ (.A(_09649_),
    .B(_09675_),
    .Y(_09676_));
 sky130_fd_sc_hd__nand3b_2 _31309_ (.A_N(_09675_),
    .B(_09646_),
    .C(_09648_),
    .Y(_09677_));
 sky130_fd_sc_hd__o21ai_2 _31310_ (.A1(_09298_),
    .A2(_09294_),
    .B1(_09301_),
    .Y(_09678_));
 sky130_fd_sc_hd__a21oi_2 _31311_ (.A1(_09676_),
    .A2(_09677_),
    .B1(_09678_),
    .Y(_09679_));
 sky130_fd_sc_hd__nand3_2 _31312_ (.A(_09676_),
    .B(_09678_),
    .C(_09677_),
    .Y(_09680_));
 sky130_vsdinv _31313_ (.A(_09680_),
    .Y(_09681_));
 sky130_fd_sc_hd__a21boi_2 _31314_ (.A1(_09382_),
    .A2(_09354_),
    .B1_N(_09356_),
    .Y(_09682_));
 sky130_fd_sc_hd__o21ai_2 _31315_ (.A1(_09679_),
    .A2(_09681_),
    .B1(_09682_),
    .Y(_09683_));
 sky130_fd_sc_hd__buf_1 _31316_ (.A(_09683_),
    .X(_09684_));
 sky130_fd_sc_hd__a21o_2 _31317_ (.A1(_09676_),
    .A2(_09677_),
    .B1(_09678_),
    .X(_09685_));
 sky130_fd_sc_hd__nand3b_2 _31318_ (.A_N(_09682_),
    .B(_09685_),
    .C(_09680_),
    .Y(_09686_));
 sky130_fd_sc_hd__buf_1 _31319_ (.A(_09686_),
    .X(_09687_));
 sky130_fd_sc_hd__a22oi_2 _31320_ (.A1(_09623_),
    .A2(_09626_),
    .B1(_09684_),
    .B2(_09687_),
    .Y(_09688_));
 sky130_fd_sc_hd__nand2_2 _31321_ (.A(_09623_),
    .B(_09626_),
    .Y(_09689_));
 sky130_fd_sc_hd__nand2_2 _31322_ (.A(_09683_),
    .B(_09686_),
    .Y(_09690_));
 sky130_fd_sc_hd__nor2_2 _31323_ (.A(_09689_),
    .B(_09690_),
    .Y(_09691_));
 sky130_fd_sc_hd__a31oi_2 _31324_ (.A1(_09392_),
    .A2(_09330_),
    .A3(_09396_),
    .B1(_09404_),
    .Y(_09692_));
 sky130_fd_sc_hd__o21ai_2 _31325_ (.A1(_09688_),
    .A2(_09691_),
    .B1(_09692_),
    .Y(_09693_));
 sky130_fd_sc_hd__buf_1 _31326_ (.A(_09693_),
    .X(_09694_));
 sky130_fd_sc_hd__a31o_2 _31327_ (.A1(_09392_),
    .A2(_09330_),
    .A3(_09396_),
    .B1(_09404_),
    .X(_09695_));
 sky130_fd_sc_hd__a21oi_2 _31328_ (.A1(_09624_),
    .A2(_09625_),
    .B1(_09329_),
    .Y(_09696_));
 sky130_fd_sc_hd__nor3_2 _31329_ (.A(_09332_),
    .B(_09617_),
    .C(_09622_),
    .Y(_09697_));
 sky130_fd_sc_hd__nor2_2 _31330_ (.A(_09696_),
    .B(_09697_),
    .Y(_09698_));
 sky130_fd_sc_hd__nand3_2 _31331_ (.A(_09698_),
    .B(_09687_),
    .C(_09684_),
    .Y(_09699_));
 sky130_fd_sc_hd__nand2_2 _31332_ (.A(_09690_),
    .B(_09689_),
    .Y(_09700_));
 sky130_fd_sc_hd__nand3_2 _31333_ (.A(_09695_),
    .B(_09699_),
    .C(_09700_),
    .Y(_09701_));
 sky130_fd_sc_hd__a22oi_2 _31334_ (.A1(_09544_),
    .A2(_09547_),
    .B1(_09694_),
    .B2(_09701_),
    .Y(_09702_));
 sky130_fd_sc_hd__nand2_2 _31335_ (.A(_09544_),
    .B(_09546_),
    .Y(_09703_));
 sky130_fd_sc_hd__nand2_2 _31336_ (.A(_09694_),
    .B(_09701_),
    .Y(_09704_));
 sky130_fd_sc_hd__nor2_2 _31337_ (.A(_09703_),
    .B(_09704_),
    .Y(_09705_));
 sky130_fd_sc_hd__a21oi_2 _31338_ (.A1(_09406_),
    .A2(_09407_),
    .B1(_09401_),
    .Y(_09706_));
 sky130_fd_sc_hd__o21a_2 _31339_ (.A1(_09706_),
    .A2(_09411_),
    .B1(_09409_),
    .X(_09707_));
 sky130_fd_sc_hd__o21ai_2 _31340_ (.A1(_09702_),
    .A2(_09705_),
    .B1(_09707_),
    .Y(_09708_));
 sky130_fd_sc_hd__a21boi_2 _31341_ (.A1(_09538_),
    .A2(_09545_),
    .B1_N(_09543_),
    .Y(_09709_));
 sky130_fd_sc_hd__nor2_2 _31342_ (.A(_09543_),
    .B(_09542_),
    .Y(_09710_));
 sky130_fd_sc_hd__nor2_2 _31343_ (.A(_09709_),
    .B(_09710_),
    .Y(_09711_));
 sky130_fd_sc_hd__nand3_2 _31344_ (.A(_09711_),
    .B(_09701_),
    .C(_09694_),
    .Y(_09712_));
 sky130_fd_sc_hd__o21ai_2 _31345_ (.A1(_09706_),
    .A2(_09411_),
    .B1(_09409_),
    .Y(_09713_));
 sky130_fd_sc_hd__nand2_2 _31346_ (.A(_09704_),
    .B(_09703_),
    .Y(_09714_));
 sky130_fd_sc_hd__nand3_2 _31347_ (.A(_09712_),
    .B(_09713_),
    .C(_09714_),
    .Y(_09715_));
 sky130_fd_sc_hd__nand2_2 _31348_ (.A(_09708_),
    .B(_09715_),
    .Y(_09716_));
 sky130_fd_sc_hd__a21boi_2 _31349_ (.A1(_09238_),
    .A2(_09244_),
    .B1_N(_09239_),
    .Y(_09717_));
 sky130_fd_sc_hd__nand2_2 _31350_ (.A(_09262_),
    .B(_09256_),
    .Y(_09718_));
 sky130_fd_sc_hd__xnor2_2 _31351_ (.A(_09717_),
    .B(_09718_),
    .Y(_09719_));
 sky130_vsdinv _31352_ (.A(_09719_),
    .Y(_09720_));
 sky130_fd_sc_hd__nand2_2 _31353_ (.A(_09716_),
    .B(_09720_),
    .Y(_09721_));
 sky130_fd_sc_hd__nand3_2 _31354_ (.A(_09708_),
    .B(_09715_),
    .C(_09719_),
    .Y(_09722_));
 sky130_fd_sc_hd__nand2_2 _31355_ (.A(_09429_),
    .B(_09423_),
    .Y(_09723_));
 sky130_fd_sc_hd__a21oi_2 _31356_ (.A1(_09721_),
    .A2(_09722_),
    .B1(_09723_),
    .Y(_09724_));
 sky130_fd_sc_hd__a21boi_2 _31357_ (.A1(_09415_),
    .A2(_09427_),
    .B1_N(_09423_),
    .Y(_09725_));
 sky130_fd_sc_hd__nand2_2 _31358_ (.A(_09721_),
    .B(_09722_),
    .Y(_09726_));
 sky130_fd_sc_hd__nor2_2 _31359_ (.A(_09725_),
    .B(_09726_),
    .Y(_09727_));
 sky130_fd_sc_hd__buf_1 _31360_ (.A(_09425_),
    .X(_09728_));
 sky130_fd_sc_hd__o21bai_2 _31361_ (.A1(_09724_),
    .A2(_09727_),
    .B1_N(_09728_),
    .Y(_09729_));
 sky130_fd_sc_hd__nand2_2 _31362_ (.A(_09726_),
    .B(_09725_),
    .Y(_09730_));
 sky130_fd_sc_hd__nand3_2 _31363_ (.A(_09723_),
    .B(_09722_),
    .C(_09721_),
    .Y(_09731_));
 sky130_fd_sc_hd__nand3_2 _31364_ (.A(_09730_),
    .B(_09728_),
    .C(_09731_),
    .Y(_09732_));
 sky130_vsdinv _31365_ (.A(_09437_),
    .Y(_09733_));
 sky130_fd_sc_hd__o21ai_2 _31366_ (.A1(_09733_),
    .A2(_09445_),
    .B1(_09436_),
    .Y(_09734_));
 sky130_fd_sc_hd__a21oi_2 _31367_ (.A1(_09729_),
    .A2(_09732_),
    .B1(_09734_),
    .Y(_09735_));
 sky130_fd_sc_hd__a21oi_2 _31368_ (.A1(_09730_),
    .A2(_09731_),
    .B1(_09728_),
    .Y(_09736_));
 sky130_fd_sc_hd__a21boi_2 _31369_ (.A1(_09433_),
    .A2(_09438_),
    .B1_N(_09436_),
    .Y(_09737_));
 sky130_vsdinv _31370_ (.A(_09425_),
    .Y(_09738_));
 sky130_fd_sc_hd__nor3_2 _31371_ (.A(_09738_),
    .B(_09724_),
    .C(_09727_),
    .Y(_09739_));
 sky130_fd_sc_hd__nor3_2 _31372_ (.A(_09736_),
    .B(_09737_),
    .C(_09739_),
    .Y(_09740_));
 sky130_fd_sc_hd__nor2_2 _31373_ (.A(_09735_),
    .B(_09740_),
    .Y(_09741_));
 sky130_fd_sc_hd__nand2_2 _31374_ (.A(_09452_),
    .B(_09166_),
    .Y(_09742_));
 sky130_fd_sc_hd__nor2_2 _31375_ (.A(_09742_),
    .B(_09449_),
    .Y(_09743_));
 sky130_fd_sc_hd__nor2_2 _31376_ (.A(_08649_),
    .B(_08899_),
    .Y(_09744_));
 sky130_fd_sc_hd__nand2_2 _31377_ (.A(_09743_),
    .B(_09744_),
    .Y(_09745_));
 sky130_fd_sc_hd__a21oi_2 _31378_ (.A1(_09447_),
    .A2(_09440_),
    .B1(_09443_),
    .Y(_09746_));
 sky130_vsdinv _31379_ (.A(_09448_),
    .Y(_09747_));
 sky130_fd_sc_hd__nor2_2 _31380_ (.A(_09746_),
    .B(_09747_),
    .Y(_09748_));
 sky130_fd_sc_hd__nand3_2 _31381_ (.A(_09748_),
    .B(_09168_),
    .C(_09170_),
    .Y(_09749_));
 sky130_fd_sc_hd__a21oi_2 _31382_ (.A1(_09167_),
    .A2(_09444_),
    .B1(_09747_),
    .Y(_09750_));
 sky130_fd_sc_hd__nand2_2 _31383_ (.A(_09749_),
    .B(_09750_),
    .Y(_09751_));
 sky130_fd_sc_hd__o21bai_2 _31384_ (.A1(_09745_),
    .A2(_08657_),
    .B1_N(_09751_),
    .Y(_09752_));
 sky130_fd_sc_hd__xor2_2 _31385_ (.A(_09741_),
    .B(_09752_),
    .X(_02647_));
 sky130_fd_sc_hd__a22oi_2 _31386_ (.A1(_07548_),
    .A2(_09456_),
    .B1(_06226_),
    .B2(_19185_),
    .Y(_09753_));
 sky130_fd_sc_hd__nand2_2 _31387_ (.A(_06881_),
    .B(_07733_),
    .Y(_09754_));
 sky130_fd_sc_hd__buf_1 _31388_ (.A(_08825_),
    .X(_09755_));
 sky130_fd_sc_hd__nand2_2 _31389_ (.A(_05768_),
    .B(_09755_),
    .Y(_09756_));
 sky130_fd_sc_hd__nor2_2 _31390_ (.A(_09754_),
    .B(_09756_),
    .Y(_09757_));
 sky130_fd_sc_hd__and2_2 _31391_ (.A(_05586_),
    .B(_09495_),
    .X(_09758_));
 sky130_fd_sc_hd__o21bai_2 _31392_ (.A1(_09753_),
    .A2(_09757_),
    .B1_N(_09758_),
    .Y(_09759_));
 sky130_fd_sc_hd__nand3b_2 _31393_ (.A_N(_09754_),
    .B(_05993_),
    .C(_09079_),
    .Y(_09760_));
 sky130_fd_sc_hd__nand3b_2 _31394_ (.A_N(_09753_),
    .B(_09760_),
    .C(_09758_),
    .Y(_09761_));
 sky130_fd_sc_hd__nand2_2 _31395_ (.A(_09759_),
    .B(_09761_),
    .Y(_09762_));
 sky130_fd_sc_hd__a21oi_2 _31396_ (.A1(_09662_),
    .A2(_09667_),
    .B1(_09663_),
    .Y(_09763_));
 sky130_fd_sc_hd__nand2_2 _31397_ (.A(_09762_),
    .B(_09763_),
    .Y(_09764_));
 sky130_fd_sc_hd__nand3b_2 _31398_ (.A_N(_09763_),
    .B(_09759_),
    .C(_09761_),
    .Y(_09765_));
 sky130_fd_sc_hd__a21oi_2 _31399_ (.A1(_09462_),
    .A2(_09459_),
    .B1(_09458_),
    .Y(_09766_));
 sky130_vsdinv _31400_ (.A(_09766_),
    .Y(_09767_));
 sky130_fd_sc_hd__a21oi_2 _31401_ (.A1(_09764_),
    .A2(_09765_),
    .B1(_09767_),
    .Y(_09768_));
 sky130_fd_sc_hd__nand3_2 _31402_ (.A(_09764_),
    .B(_09767_),
    .C(_09765_),
    .Y(_09769_));
 sky130_vsdinv _31403_ (.A(_09769_),
    .Y(_09770_));
 sky130_fd_sc_hd__o21ai_2 _31404_ (.A1(_09669_),
    .A2(_09659_),
    .B1(_09671_),
    .Y(_09771_));
 sky130_fd_sc_hd__o21bai_2 _31405_ (.A1(_09768_),
    .A2(_09770_),
    .B1_N(_09771_),
    .Y(_09772_));
 sky130_fd_sc_hd__nand2_2 _31406_ (.A(_09764_),
    .B(_09765_),
    .Y(_09773_));
 sky130_fd_sc_hd__nand2_2 _31407_ (.A(_09773_),
    .B(_09766_),
    .Y(_09774_));
 sky130_fd_sc_hd__nand3_2 _31408_ (.A(_09774_),
    .B(_09771_),
    .C(_09769_),
    .Y(_09775_));
 sky130_fd_sc_hd__nand2_2 _31409_ (.A(_09772_),
    .B(_09775_),
    .Y(_09776_));
 sky130_fd_sc_hd__a21boi_2 _31410_ (.A1(_09466_),
    .A2(_09469_),
    .B1_N(_09467_),
    .Y(_09777_));
 sky130_fd_sc_hd__nand2_2 _31411_ (.A(_09776_),
    .B(_09777_),
    .Y(_09778_));
 sky130_fd_sc_hd__nand3b_2 _31412_ (.A_N(_09777_),
    .B(_09772_),
    .C(_09775_),
    .Y(_09779_));
 sky130_fd_sc_hd__nand2_2 _31413_ (.A(_09778_),
    .B(_09779_),
    .Y(_09780_));
 sky130_fd_sc_hd__a21boi_2 _31414_ (.A1(_09475_),
    .A2(_09481_),
    .B1_N(_09478_),
    .Y(_09781_));
 sky130_fd_sc_hd__nand2_2 _31415_ (.A(_09780_),
    .B(_09781_),
    .Y(_09782_));
 sky130_fd_sc_hd__nand3b_2 _31416_ (.A_N(_09781_),
    .B(_09779_),
    .C(_09778_),
    .Y(_09783_));
 sky130_fd_sc_hd__nand2_2 _31417_ (.A(_09782_),
    .B(_09783_),
    .Y(_09784_));
 sky130_fd_sc_hd__buf_1 _31418_ (.A(_09493_),
    .X(_09785_));
 sky130_fd_sc_hd__buf_1 _31419_ (.A(_19166_),
    .X(_09786_));
 sky130_fd_sc_hd__buf_1 _31420_ (.A(_09786_),
    .X(_09787_));
 sky130_fd_sc_hd__a22oi_2 _31421_ (.A1(_05566_),
    .A2(_09785_),
    .B1(_05940_),
    .B2(_09787_),
    .Y(_09788_));
 sky130_fd_sc_hd__nand2_2 _31422_ (.A(_18844_),
    .B(_08557_),
    .Y(_09789_));
 sky130_fd_sc_hd__buf_1 _31423_ (.A(_09086_),
    .X(_09790_));
 sky130_fd_sc_hd__nand2_2 _31424_ (.A(_05939_),
    .B(_09790_),
    .Y(_09791_));
 sky130_fd_sc_hd__nor2_2 _31425_ (.A(_09789_),
    .B(_09791_),
    .Y(_09792_));
 sky130_fd_sc_hd__buf_1 _31426_ (.A(_19143_),
    .X(_09793_));
 sky130_fd_sc_hd__and2_2 _31427_ (.A(_06732_),
    .B(_09793_),
    .X(_09794_));
 sky130_fd_sc_hd__o21bai_2 _31428_ (.A1(_09788_),
    .A2(_09792_),
    .B1_N(_09794_),
    .Y(_09795_));
 sky130_fd_sc_hd__nand2_2 _31429_ (.A(_09789_),
    .B(_09791_),
    .Y(_09796_));
 sky130_fd_sc_hd__nand3b_2 _31430_ (.A_N(_09792_),
    .B(_09796_),
    .C(_09794_),
    .Y(_09797_));
 sky130_fd_sc_hd__nand2_2 _31431_ (.A(_09502_),
    .B(_09498_),
    .Y(_09798_));
 sky130_fd_sc_hd__a21o_2 _31432_ (.A1(_09795_),
    .A2(_09797_),
    .B1(_09798_),
    .X(_09799_));
 sky130_fd_sc_hd__nand3_2 _31433_ (.A(_09798_),
    .B(_09795_),
    .C(_09797_),
    .Y(_09800_));
 sky130_fd_sc_hd__nand2_2 _31434_ (.A(_09799_),
    .B(_09800_),
    .Y(_09801_));
 sky130_fd_sc_hd__buf_1 _31435_ (.A(_09212_),
    .X(_09802_));
 sky130_fd_sc_hd__nand2_2 _31436_ (.A(_05662_),
    .B(_09802_),
    .Y(_09803_));
 sky130_fd_sc_hd__buf_1 _31437_ (.A(\pcpi_mul.rs1[28] ),
    .X(_09804_));
 sky130_fd_sc_hd__buf_1 _31438_ (.A(_09804_),
    .X(_09805_));
 sky130_fd_sc_hd__nand2_2 _31439_ (.A(_18872_),
    .B(_09805_),
    .Y(_09806_));
 sky130_fd_sc_hd__xor2_2 _31440_ (.A(_09803_),
    .B(_09806_),
    .X(_09807_));
 sky130_fd_sc_hd__buf_1 _31441_ (.A(_09224_),
    .X(_09808_));
 sky130_fd_sc_hd__buf_1 _31442_ (.A(_09808_),
    .X(_09809_));
 sky130_fd_sc_hd__and2_2 _31443_ (.A(_07121_),
    .B(_09809_),
    .X(_09810_));
 sky130_fd_sc_hd__nand2_2 _31444_ (.A(_09807_),
    .B(_09810_),
    .Y(_09811_));
 sky130_fd_sc_hd__xnor2_2 _31445_ (.A(_09803_),
    .B(_09806_),
    .Y(_09812_));
 sky130_fd_sc_hd__o21ai_2 _31446_ (.A1(_06923_),
    .A2(_19163_),
    .B1(_09812_),
    .Y(_09813_));
 sky130_fd_sc_hd__nand2_2 _31447_ (.A(_09811_),
    .B(_09813_),
    .Y(_09814_));
 sky130_fd_sc_hd__nand2_2 _31448_ (.A(_09801_),
    .B(_09814_),
    .Y(_09815_));
 sky130_fd_sc_hd__nand3b_2 _31449_ (.A_N(_09814_),
    .B(_09799_),
    .C(_09800_),
    .Y(_09816_));
 sky130_fd_sc_hd__o21ai_2 _31450_ (.A1(_09517_),
    .A2(_09519_),
    .B1(_09507_),
    .Y(_09817_));
 sky130_fd_sc_hd__a21oi_2 _31451_ (.A1(_09815_),
    .A2(_09816_),
    .B1(_09817_),
    .Y(_09818_));
 sky130_fd_sc_hd__nand3_2 _31452_ (.A(_09815_),
    .B(_09816_),
    .C(_09817_),
    .Y(_09819_));
 sky130_vsdinv _31453_ (.A(_09819_),
    .Y(_09820_));
 sky130_fd_sc_hd__o21a_2 _31454_ (.A1(_09508_),
    .A2(_09509_),
    .B1(_09513_),
    .X(_09821_));
 sky130_vsdinv _31455_ (.A(_09821_),
    .Y(_09822_));
 sky130_fd_sc_hd__o21bai_2 _31456_ (.A1(_09818_),
    .A2(_09820_),
    .B1_N(_09822_),
    .Y(_09823_));
 sky130_fd_sc_hd__nand3b_2 _31457_ (.A_N(_09818_),
    .B(_09822_),
    .C(_09819_),
    .Y(_09824_));
 sky130_fd_sc_hd__nand2_2 _31458_ (.A(_09823_),
    .B(_09824_),
    .Y(_09825_));
 sky130_fd_sc_hd__nand2_2 _31459_ (.A(_09784_),
    .B(_09825_),
    .Y(_09826_));
 sky130_fd_sc_hd__nand3b_2 _31460_ (.A_N(_09825_),
    .B(_09783_),
    .C(_09782_),
    .Y(_09827_));
 sky130_fd_sc_hd__o21ai_2 _31461_ (.A1(_09682_),
    .A2(_09679_),
    .B1(_09680_),
    .Y(_09828_));
 sky130_fd_sc_hd__a21oi_2 _31462_ (.A1(_09826_),
    .A2(_09827_),
    .B1(_09828_),
    .Y(_09829_));
 sky130_fd_sc_hd__nand3_2 _31463_ (.A(_09826_),
    .B(_09827_),
    .C(_09828_),
    .Y(_09830_));
 sky130_vsdinv _31464_ (.A(_09830_),
    .Y(_09831_));
 sky130_fd_sc_hd__o21a_2 _31465_ (.A1(_09533_),
    .A2(_09535_),
    .B1(_09491_),
    .X(_09832_));
 sky130_fd_sc_hd__buf_1 _31466_ (.A(_09832_),
    .X(_09833_));
 sky130_fd_sc_hd__o21ai_2 _31467_ (.A1(_09829_),
    .A2(_09831_),
    .B1(_09833_),
    .Y(_09834_));
 sky130_fd_sc_hd__nand2_2 _31468_ (.A(_09826_),
    .B(_09827_),
    .Y(_09835_));
 sky130_vsdinv _31469_ (.A(_09828_),
    .Y(_09836_));
 sky130_fd_sc_hd__nand2_2 _31470_ (.A(_09835_),
    .B(_09836_),
    .Y(_09837_));
 sky130_fd_sc_hd__buf_1 _31471_ (.A(_09830_),
    .X(_09838_));
 sky130_fd_sc_hd__nand3b_2 _31472_ (.A_N(_09832_),
    .B(_09837_),
    .C(_09838_),
    .Y(_09839_));
 sky130_fd_sc_hd__a22oi_2 _31473_ (.A1(_18779_),
    .A2(_06186_),
    .B1(_18784_),
    .B2(_07099_),
    .Y(_09840_));
 sky130_fd_sc_hd__nand2_2 _31474_ (.A(_07164_),
    .B(_06462_),
    .Y(_09841_));
 sky130_fd_sc_hd__nand2_2 _31475_ (.A(_07394_),
    .B(_07690_),
    .Y(_09842_));
 sky130_fd_sc_hd__nor2_2 _31476_ (.A(_09841_),
    .B(_09842_),
    .Y(_09843_));
 sky130_fd_sc_hd__and2_2 _31477_ (.A(_18789_),
    .B(_19230_),
    .X(_09844_));
 sky130_fd_sc_hd__o21bai_2 _31478_ (.A1(_09840_),
    .A2(_09843_),
    .B1_N(_09844_),
    .Y(_09845_));
 sky130_fd_sc_hd__nand3b_2 _31479_ (.A_N(_09841_),
    .B(_08012_),
    .C(_19237_),
    .Y(_09846_));
 sky130_fd_sc_hd__nand3b_2 _31480_ (.A_N(_09840_),
    .B(_09846_),
    .C(_09844_),
    .Y(_09847_));
 sky130_fd_sc_hd__nand2_2 _31481_ (.A(_09845_),
    .B(_09847_),
    .Y(_09848_));
 sky130_fd_sc_hd__a21oi_2 _31482_ (.A1(_09568_),
    .A2(_09570_),
    .B1(_09567_),
    .Y(_09849_));
 sky130_fd_sc_hd__nand2_2 _31483_ (.A(_09848_),
    .B(_09849_),
    .Y(_09850_));
 sky130_fd_sc_hd__nand3b_2 _31484_ (.A_N(_09849_),
    .B(_09847_),
    .C(_09845_),
    .Y(_09851_));
 sky130_fd_sc_hd__buf_1 _31485_ (.A(_09851_),
    .X(_09852_));
 sky130_fd_sc_hd__a21oi_2 _31486_ (.A1(_09631_),
    .A2(_09630_),
    .B1(_09629_),
    .Y(_09853_));
 sky130_vsdinv _31487_ (.A(_09853_),
    .Y(_09854_));
 sky130_fd_sc_hd__a21oi_2 _31488_ (.A1(_09850_),
    .A2(_09852_),
    .B1(_09854_),
    .Y(_09855_));
 sky130_fd_sc_hd__nand3_2 _31489_ (.A(_09850_),
    .B(_09854_),
    .C(_09852_),
    .Y(_09856_));
 sky130_vsdinv _31490_ (.A(_09856_),
    .Y(_09857_));
 sky130_fd_sc_hd__a21boi_2 _31491_ (.A1(_09632_),
    .A2(_09634_),
    .B1_N(_09637_),
    .Y(_09858_));
 sky130_fd_sc_hd__o21ai_2 _31492_ (.A1(_09641_),
    .A2(_09858_),
    .B1(_09639_),
    .Y(_09859_));
 sky130_fd_sc_hd__o21bai_2 _31493_ (.A1(_09855_),
    .A2(_09857_),
    .B1_N(_09859_),
    .Y(_09860_));
 sky130_fd_sc_hd__nand2_2 _31494_ (.A(_09850_),
    .B(_09851_),
    .Y(_09861_));
 sky130_fd_sc_hd__nand2_2 _31495_ (.A(_09861_),
    .B(_09853_),
    .Y(_09862_));
 sky130_fd_sc_hd__nand3_2 _31496_ (.A(_09862_),
    .B(_09859_),
    .C(_09856_),
    .Y(_09863_));
 sky130_fd_sc_hd__nand2_2 _31497_ (.A(_06533_),
    .B(_06744_),
    .Y(_09864_));
 sky130_fd_sc_hd__nand2_2 _31498_ (.A(_06536_),
    .B(_07115_),
    .Y(_09865_));
 sky130_fd_sc_hd__nor2_2 _31499_ (.A(_09864_),
    .B(_09865_),
    .Y(_09866_));
 sky130_fd_sc_hd__and2_2 _31500_ (.A(_08038_),
    .B(_07946_),
    .X(_09867_));
 sky130_fd_sc_hd__nand2_2 _31501_ (.A(_09864_),
    .B(_09865_),
    .Y(_09868_));
 sky130_fd_sc_hd__nand3b_2 _31502_ (.A_N(_09866_),
    .B(_09867_),
    .C(_09868_),
    .Y(_09869_));
 sky130_fd_sc_hd__buf_1 _31503_ (.A(_06536_),
    .X(_09870_));
 sky130_fd_sc_hd__a22oi_2 _31504_ (.A1(_08414_),
    .A2(_08262_),
    .B1(_09870_),
    .B2(_08510_),
    .Y(_09871_));
 sky130_fd_sc_hd__o21bai_2 _31505_ (.A1(_09871_),
    .A2(_09866_),
    .B1_N(_09867_),
    .Y(_09872_));
 sky130_fd_sc_hd__a21oi_2 _31506_ (.A1(_09654_),
    .A2(_09653_),
    .B1(_09652_),
    .Y(_09873_));
 sky130_fd_sc_hd__a21boi_2 _31507_ (.A1(_09869_),
    .A2(_09872_),
    .B1_N(_09873_),
    .Y(_09874_));
 sky130_fd_sc_hd__nand2_2 _31508_ (.A(_06810_),
    .B(_07105_),
    .Y(_09875_));
 sky130_fd_sc_hd__nand2_2 _31509_ (.A(_08180_),
    .B(_07743_),
    .Y(_09876_));
 sky130_fd_sc_hd__nand2_2 _31510_ (.A(_09875_),
    .B(_09876_),
    .Y(_09877_));
 sky130_fd_sc_hd__nor2_2 _31511_ (.A(_09875_),
    .B(_09876_),
    .Y(_09878_));
 sky130_vsdinv _31512_ (.A(_09878_),
    .Y(_09879_));
 sky130_fd_sc_hd__o2bb2ai_2 _31513_ (.A1_N(_09877_),
    .A2_N(_09879_),
    .B1(_07214_),
    .B2(_19197_),
    .Y(_09880_));
 sky130_fd_sc_hd__and2_2 _31514_ (.A(_06137_),
    .B(_08812_),
    .X(_09881_));
 sky130_fd_sc_hd__nand3b_2 _31515_ (.A_N(_09878_),
    .B(_09881_),
    .C(_09877_),
    .Y(_09882_));
 sky130_fd_sc_hd__nand2_2 _31516_ (.A(_09880_),
    .B(_09882_),
    .Y(_09883_));
 sky130_vsdinv _31517_ (.A(_09883_),
    .Y(_09884_));
 sky130_fd_sc_hd__nand3b_2 _31518_ (.A_N(_09873_),
    .B(_09869_),
    .C(_09872_),
    .Y(_09885_));
 sky130_fd_sc_hd__nand3b_2 _31519_ (.A_N(_09874_),
    .B(_09884_),
    .C(_09885_),
    .Y(_09886_));
 sky130_vsdinv _31520_ (.A(_09885_),
    .Y(_09887_));
 sky130_fd_sc_hd__o21ai_2 _31521_ (.A1(_09874_),
    .A2(_09887_),
    .B1(_09883_),
    .Y(_09888_));
 sky130_fd_sc_hd__nand2_2 _31522_ (.A(_09886_),
    .B(_09888_),
    .Y(_09889_));
 sky130_fd_sc_hd__buf_1 _31523_ (.A(_09889_),
    .X(_09890_));
 sky130_fd_sc_hd__a21boi_2 _31524_ (.A1(_09860_),
    .A2(_09863_),
    .B1_N(_09890_),
    .Y(_09891_));
 sky130_fd_sc_hd__a21oi_2 _31525_ (.A1(_09862_),
    .A2(_09856_),
    .B1(_09859_),
    .Y(_09892_));
 sky130_vsdinv _31526_ (.A(_09863_),
    .Y(_09893_));
 sky130_fd_sc_hd__nor3_2 _31527_ (.A(_09890_),
    .B(_09892_),
    .C(_09893_),
    .Y(_09894_));
 sky130_fd_sc_hd__a21oi_2 _31528_ (.A1(_09580_),
    .A2(_09581_),
    .B1(_09578_),
    .Y(_09895_));
 sky130_fd_sc_hd__o21ai_2 _31529_ (.A1(_09584_),
    .A2(_09895_),
    .B1(_09582_),
    .Y(_09896_));
 sky130_fd_sc_hd__o21bai_2 _31530_ (.A1(_09891_),
    .A2(_09894_),
    .B1_N(_09896_),
    .Y(_09897_));
 sky130_fd_sc_hd__o21ai_2 _31531_ (.A1(_09892_),
    .A2(_09893_),
    .B1(_09890_),
    .Y(_09898_));
 sky130_fd_sc_hd__nand3b_2 _31532_ (.A_N(_09889_),
    .B(_09860_),
    .C(_09863_),
    .Y(_09899_));
 sky130_fd_sc_hd__nand3_2 _31533_ (.A(_09898_),
    .B(_09896_),
    .C(_09899_),
    .Y(_09900_));
 sky130_fd_sc_hd__nand2_2 _31534_ (.A(_09897_),
    .B(_09900_),
    .Y(_09901_));
 sky130_fd_sc_hd__o21a_2 _31535_ (.A1(_09644_),
    .A2(_09645_),
    .B1(_09677_),
    .X(_09902_));
 sky130_fd_sc_hd__nand2_2 _31536_ (.A(_09901_),
    .B(_09902_),
    .Y(_09903_));
 sky130_fd_sc_hd__nand3b_2 _31537_ (.A_N(_09902_),
    .B(_09897_),
    .C(_09900_),
    .Y(_09904_));
 sky130_fd_sc_hd__nand2_2 _31538_ (.A(_07537_),
    .B(_06060_),
    .Y(_09905_));
 sky130_fd_sc_hd__nand2_2 _31539_ (.A(_18770_),
    .B(_07382_),
    .Y(_09906_));
 sky130_fd_sc_hd__nor2_2 _31540_ (.A(_09905_),
    .B(_09906_),
    .Y(_09907_));
 sky130_fd_sc_hd__and2_2 _31541_ (.A(_18775_),
    .B(_06588_),
    .X(_09908_));
 sky130_fd_sc_hd__nand2_2 _31542_ (.A(_09905_),
    .B(_09906_),
    .Y(_09909_));
 sky130_fd_sc_hd__and3b_2 _31543_ (.A_N(_09907_),
    .B(_09908_),
    .C(_09909_),
    .X(_09910_));
 sky130_vsdinv _31544_ (.A(_09907_),
    .Y(_09911_));
 sky130_fd_sc_hd__a21oi_2 _31545_ (.A1(_09911_),
    .A2(_09909_),
    .B1(_09908_),
    .Y(_09912_));
 sky130_fd_sc_hd__a22oi_2 _31546_ (.A1(_08729_),
    .A2(_05739_),
    .B1(_08224_),
    .B2(_05741_),
    .Y(_09913_));
 sky130_fd_sc_hd__nand2_2 _31547_ (.A(_18747_),
    .B(_08480_),
    .Y(_09914_));
 sky130_fd_sc_hd__nand2_2 _31548_ (.A(_08224_),
    .B(_05963_),
    .Y(_09915_));
 sky130_fd_sc_hd__nor2_2 _31549_ (.A(_09914_),
    .B(_09915_),
    .Y(_09916_));
 sky130_fd_sc_hd__nand2_2 _31550_ (.A(_07844_),
    .B(_05846_),
    .Y(_09917_));
 sky130_vsdinv _31551_ (.A(_09917_),
    .Y(_09918_));
 sky130_fd_sc_hd__o21bai_2 _31552_ (.A1(_09913_),
    .A2(_09916_),
    .B1_N(_09918_),
    .Y(_09919_));
 sky130_fd_sc_hd__nand3b_2 _31553_ (.A_N(_09914_),
    .B(_09548_),
    .C(_06043_),
    .Y(_09920_));
 sky130_fd_sc_hd__nand2_2 _31554_ (.A(_09914_),
    .B(_09915_),
    .Y(_09921_));
 sky130_fd_sc_hd__nand3_2 _31555_ (.A(_09920_),
    .B(_09918_),
    .C(_09921_),
    .Y(_09922_));
 sky130_fd_sc_hd__o21ai_2 _31556_ (.A1(_09553_),
    .A2(_09549_),
    .B1(_09556_),
    .Y(_09923_));
 sky130_fd_sc_hd__a21oi_2 _31557_ (.A1(_09919_),
    .A2(_09922_),
    .B1(_09923_),
    .Y(_09924_));
 sky130_fd_sc_hd__nand3_2 _31558_ (.A(_09919_),
    .B(_09922_),
    .C(_09923_),
    .Y(_09925_));
 sky130_vsdinv _31559_ (.A(_09925_),
    .Y(_09926_));
 sky130_fd_sc_hd__o22ai_2 _31560_ (.A1(_09910_),
    .A2(_09912_),
    .B1(_09924_),
    .B2(_09926_),
    .Y(_09927_));
 sky130_fd_sc_hd__nor2_2 _31561_ (.A(_09912_),
    .B(_09910_),
    .Y(_09928_));
 sky130_fd_sc_hd__a21o_2 _31562_ (.A1(_09919_),
    .A2(_09922_),
    .B1(_09923_),
    .X(_09929_));
 sky130_fd_sc_hd__nand3_2 _31563_ (.A(_09928_),
    .B(_09929_),
    .C(_09925_),
    .Y(_09930_));
 sky130_fd_sc_hd__nand2_2 _31564_ (.A(_09927_),
    .B(_09930_),
    .Y(_09931_));
 sky130_fd_sc_hd__nand2_2 _31565_ (.A(_09931_),
    .B(_09601_),
    .Y(_09932_));
 sky130_fd_sc_hd__nand3b_2 _31566_ (.A_N(_09601_),
    .B(_09927_),
    .C(_09930_),
    .Y(_09933_));
 sky130_fd_sc_hd__nand2_2 _31567_ (.A(_09932_),
    .B(_09933_),
    .Y(_09934_));
 sky130_fd_sc_hd__o21a_2 _31568_ (.A1(_09574_),
    .A2(_09576_),
    .B1(_09564_),
    .X(_09935_));
 sky130_fd_sc_hd__nand2_2 _31569_ (.A(_09934_),
    .B(_09935_),
    .Y(_09936_));
 sky130_vsdinv _31570_ (.A(_09935_),
    .Y(_09937_));
 sky130_fd_sc_hd__nand3_2 _31571_ (.A(_09932_),
    .B(_09937_),
    .C(_09933_),
    .Y(_09938_));
 sky130_fd_sc_hd__buf_1 _31572_ (.A(_09938_),
    .X(_09939_));
 sky130_fd_sc_hd__a22oi_2 _31573_ (.A1(_09587_),
    .A2(_06826_),
    .B1(_09589_),
    .B2(_08725_),
    .Y(_09940_));
 sky130_fd_sc_hd__and4_2 _31574_ (.A(_09303_),
    .B(_09589_),
    .C(_08725_),
    .D(_07171_),
    .X(_09941_));
 sky130_fd_sc_hd__and2_2 _31575_ (.A(_09308_),
    .B(_05668_),
    .X(_09942_));
 sky130_fd_sc_hd__o21bai_2 _31576_ (.A1(_09940_),
    .A2(_09941_),
    .B1_N(_09942_),
    .Y(_09943_));
 sky130_fd_sc_hd__nand2_2 _31577_ (.A(_18727_),
    .B(_05986_),
    .Y(_09944_));
 sky130_fd_sc_hd__nand3b_2 _31578_ (.A_N(_09944_),
    .B(_08755_),
    .C(_07790_),
    .Y(_09945_));
 sky130_fd_sc_hd__nand3b_2 _31579_ (.A_N(_09940_),
    .B(_09945_),
    .C(_09942_),
    .Y(_09946_));
 sky130_fd_sc_hd__nand2_2 _31580_ (.A(_09943_),
    .B(_09946_),
    .Y(_09947_));
 sky130_fd_sc_hd__nor2_2 _31581_ (.A(_09604_),
    .B(_09607_),
    .Y(_09948_));
 sky130_vsdinv _31582_ (.A(_09948_),
    .Y(_09949_));
 sky130_fd_sc_hd__nand2_2 _31583_ (.A(_09947_),
    .B(_09949_),
    .Y(_09950_));
 sky130_fd_sc_hd__nand3_2 _31584_ (.A(_09943_),
    .B(_09946_),
    .C(_09948_),
    .Y(_09951_));
 sky130_fd_sc_hd__a21oi_2 _31585_ (.A1(_09592_),
    .A2(_09594_),
    .B1(_09591_),
    .Y(_09952_));
 sky130_vsdinv _31586_ (.A(_09952_),
    .Y(_09953_));
 sky130_fd_sc_hd__a21o_2 _31587_ (.A1(_09950_),
    .A2(_09951_),
    .B1(_09953_),
    .X(_09954_));
 sky130_fd_sc_hd__and2_2 _31588_ (.A(_09606_),
    .B(_05431_),
    .X(_09955_));
 sky130_fd_sc_hd__nand2_2 _31589_ (.A(_09603_),
    .B(_06143_),
    .Y(_09956_));
 sky130_fd_sc_hd__buf_1 _31590_ (.A(\pcpi_mul.rs2[29] ),
    .X(_09957_));
 sky130_fd_sc_hd__buf_1 _31591_ (.A(_09957_),
    .X(_09958_));
 sky130_fd_sc_hd__nand2_2 _31592_ (.A(_09958_),
    .B(_19301_),
    .Y(_09959_));
 sky130_fd_sc_hd__xnor2_2 _31593_ (.A(_09956_),
    .B(_09959_),
    .Y(_09960_));
 sky130_fd_sc_hd__xnor2_2 _31594_ (.A(_09955_),
    .B(_09960_),
    .Y(_09961_));
 sky130_fd_sc_hd__nand3_2 _31595_ (.A(_09950_),
    .B(_09953_),
    .C(_09951_),
    .Y(_09962_));
 sky130_fd_sc_hd__nand3_2 _31596_ (.A(_09954_),
    .B(_09961_),
    .C(_09962_),
    .Y(_09963_));
 sky130_fd_sc_hd__buf_1 _31597_ (.A(_09963_),
    .X(_09964_));
 sky130_fd_sc_hd__a21oi_2 _31598_ (.A1(_09950_),
    .A2(_09951_),
    .B1(_09953_),
    .Y(_09965_));
 sky130_vsdinv _31599_ (.A(_09962_),
    .Y(_09966_));
 sky130_fd_sc_hd__o21bai_2 _31600_ (.A1(_09965_),
    .A2(_09966_),
    .B1_N(_09961_),
    .Y(_09967_));
 sky130_fd_sc_hd__o2bb2ai_2 _31601_ (.A1_N(_09964_),
    .A2_N(_09967_),
    .B1(_09609_),
    .B2(_09602_),
    .Y(_09968_));
 sky130_fd_sc_hd__nand3_2 _31602_ (.A(_09967_),
    .B(_09614_),
    .C(_09963_),
    .Y(_09969_));
 sky130_fd_sc_hd__a22oi_2 _31603_ (.A1(_09936_),
    .A2(_09939_),
    .B1(_09968_),
    .B2(_09969_),
    .Y(_09970_));
 sky130_fd_sc_hd__nand2_2 _31604_ (.A(_09936_),
    .B(_09939_),
    .Y(_09971_));
 sky130_fd_sc_hd__nand2_2 _31605_ (.A(_09968_),
    .B(_09969_),
    .Y(_09972_));
 sky130_fd_sc_hd__nor2_2 _31606_ (.A(_09971_),
    .B(_09972_),
    .Y(_09973_));
 sky130_fd_sc_hd__nand2_2 _31607_ (.A(_09625_),
    .B(_09619_),
    .Y(_09974_));
 sky130_fd_sc_hd__o21bai_2 _31608_ (.A1(_09970_),
    .A2(_09973_),
    .B1_N(_09974_),
    .Y(_09975_));
 sky130_fd_sc_hd__a21oi_2 _31609_ (.A1(_09967_),
    .A2(_09964_),
    .B1(_09614_),
    .Y(_09976_));
 sky130_vsdinv _31610_ (.A(_09969_),
    .Y(_09977_));
 sky130_fd_sc_hd__nor2_2 _31611_ (.A(_09976_),
    .B(_09977_),
    .Y(_09978_));
 sky130_fd_sc_hd__nand3_2 _31612_ (.A(_09978_),
    .B(_09939_),
    .C(_09936_),
    .Y(_09979_));
 sky130_fd_sc_hd__o21ai_2 _31613_ (.A1(_09976_),
    .A2(_09977_),
    .B1(_09971_),
    .Y(_09980_));
 sky130_fd_sc_hd__nand3_2 _31614_ (.A(_09979_),
    .B(_09980_),
    .C(_09974_),
    .Y(_09981_));
 sky130_fd_sc_hd__buf_1 _31615_ (.A(_09981_),
    .X(_09982_));
 sky130_fd_sc_hd__a22oi_2 _31616_ (.A1(_09903_),
    .A2(_09904_),
    .B1(_09975_),
    .B2(_09982_),
    .Y(_09983_));
 sky130_fd_sc_hd__nand2_2 _31617_ (.A(_09903_),
    .B(_09904_),
    .Y(_09984_));
 sky130_fd_sc_hd__buf_1 _31618_ (.A(_09984_),
    .X(_09985_));
 sky130_fd_sc_hd__nand2_2 _31619_ (.A(_09975_),
    .B(_09981_),
    .Y(_09986_));
 sky130_fd_sc_hd__nor2_2 _31620_ (.A(_09985_),
    .B(_09986_),
    .Y(_09987_));
 sky130_fd_sc_hd__a31oi_2 _31621_ (.A1(_09684_),
    .A2(_09623_),
    .A3(_09687_),
    .B1(_09697_),
    .Y(_09988_));
 sky130_fd_sc_hd__o21ai_2 _31622_ (.A1(_09983_),
    .A2(_09987_),
    .B1(_09988_),
    .Y(_09989_));
 sky130_fd_sc_hd__nand3b_2 _31623_ (.A_N(_09984_),
    .B(_09982_),
    .C(_09975_),
    .Y(_09990_));
 sky130_fd_sc_hd__a31o_2 _31624_ (.A1(_09684_),
    .A2(_09623_),
    .A3(_09687_),
    .B1(_09697_),
    .X(_09991_));
 sky130_fd_sc_hd__nand2_2 _31625_ (.A(_09986_),
    .B(_09985_),
    .Y(_09992_));
 sky130_fd_sc_hd__nand3_2 _31626_ (.A(_09990_),
    .B(_09991_),
    .C(_09992_),
    .Y(_09993_));
 sky130_fd_sc_hd__buf_1 _31627_ (.A(_09993_),
    .X(_09994_));
 sky130_fd_sc_hd__a22oi_2 _31628_ (.A1(_09834_),
    .A2(_09839_),
    .B1(_09989_),
    .B2(_09994_),
    .Y(_09995_));
 sky130_fd_sc_hd__nand2_2 _31629_ (.A(_09834_),
    .B(_09839_),
    .Y(_09996_));
 sky130_fd_sc_hd__nand2_2 _31630_ (.A(_09989_),
    .B(_09993_),
    .Y(_09997_));
 sky130_fd_sc_hd__nor2_2 _31631_ (.A(_09996_),
    .B(_09997_),
    .Y(_09998_));
 sky130_fd_sc_hd__nor3_2 _31632_ (.A(_09688_),
    .B(_09691_),
    .C(_09692_),
    .Y(_09999_));
 sky130_fd_sc_hd__a31oi_2 _31633_ (.A1(_09694_),
    .A2(_09544_),
    .A3(_09547_),
    .B1(_09999_),
    .Y(_10000_));
 sky130_fd_sc_hd__o21ai_2 _31634_ (.A1(_09995_),
    .A2(_09998_),
    .B1(_10000_),
    .Y(_10001_));
 sky130_fd_sc_hd__a31o_2 _31635_ (.A1(_09693_),
    .A2(_09546_),
    .A3(_09544_),
    .B1(_09999_),
    .X(_10002_));
 sky130_fd_sc_hd__a21boi_2 _31636_ (.A1(_09837_),
    .A2(_09838_),
    .B1_N(_09833_),
    .Y(_10003_));
 sky130_fd_sc_hd__nor3_2 _31637_ (.A(_09833_),
    .B(_09829_),
    .C(_09831_),
    .Y(_10004_));
 sky130_fd_sc_hd__nor2_2 _31638_ (.A(_10003_),
    .B(_10004_),
    .Y(_10005_));
 sky130_fd_sc_hd__nand3_2 _31639_ (.A(_10005_),
    .B(_09994_),
    .C(_09989_),
    .Y(_10006_));
 sky130_fd_sc_hd__nand2_2 _31640_ (.A(_09997_),
    .B(_09996_),
    .Y(_10007_));
 sky130_fd_sc_hd__nand3_2 _31641_ (.A(_10002_),
    .B(_10006_),
    .C(_10007_),
    .Y(_10008_));
 sky130_fd_sc_hd__nand2_2 _31642_ (.A(_10001_),
    .B(_10008_),
    .Y(_10009_));
 sky130_fd_sc_hd__o21a_2 _31643_ (.A1(_09529_),
    .A2(_09528_),
    .B1(_09527_),
    .X(_10010_));
 sky130_fd_sc_hd__nand2_2 _31644_ (.A(_09547_),
    .B(_09545_),
    .Y(_10011_));
 sky130_fd_sc_hd__xor2_2 _31645_ (.A(_10010_),
    .B(_10011_),
    .X(_10012_));
 sky130_fd_sc_hd__nand2_2 _31646_ (.A(_10009_),
    .B(_10012_),
    .Y(_10013_));
 sky130_fd_sc_hd__nand3b_2 _31647_ (.A_N(_10012_),
    .B(_10001_),
    .C(_10008_),
    .Y(_10014_));
 sky130_fd_sc_hd__nand2_2 _31648_ (.A(_10013_),
    .B(_10014_),
    .Y(_10015_));
 sky130_fd_sc_hd__a21oi_2 _31649_ (.A1(_09712_),
    .A2(_09714_),
    .B1(_09713_),
    .Y(_10016_));
 sky130_fd_sc_hd__o21ai_2 _31650_ (.A1(_09720_),
    .A2(_10016_),
    .B1(_09715_),
    .Y(_10017_));
 sky130_vsdinv _31651_ (.A(_10017_),
    .Y(_10018_));
 sky130_fd_sc_hd__nand2_2 _31652_ (.A(_10015_),
    .B(_10018_),
    .Y(_10019_));
 sky130_fd_sc_hd__nand3_2 _31653_ (.A(_10013_),
    .B(_10017_),
    .C(_10014_),
    .Y(_10020_));
 sky130_fd_sc_hd__a21oi_2 _31654_ (.A1(_09262_),
    .A2(_09256_),
    .B1(_09717_),
    .Y(_10021_));
 sky130_fd_sc_hd__a21oi_2 _31655_ (.A1(_10019_),
    .A2(_10020_),
    .B1(_10021_),
    .Y(_10022_));
 sky130_vsdinv _31656_ (.A(_10021_),
    .Y(_10023_));
 sky130_fd_sc_hd__a21oi_2 _31657_ (.A1(_10013_),
    .A2(_10014_),
    .B1(_10017_),
    .Y(_10024_));
 sky130_vsdinv _31658_ (.A(_10020_),
    .Y(_10025_));
 sky130_fd_sc_hd__nor3_2 _31659_ (.A(_10023_),
    .B(_10024_),
    .C(_10025_),
    .Y(_10026_));
 sky130_fd_sc_hd__o21ai_2 _31660_ (.A1(_09738_),
    .A2(_09724_),
    .B1(_09731_),
    .Y(_10027_));
 sky130_fd_sc_hd__o21bai_2 _31661_ (.A1(_10022_),
    .A2(_10026_),
    .B1_N(_10027_),
    .Y(_10028_));
 sky130_fd_sc_hd__o21bai_2 _31662_ (.A1(_10024_),
    .A2(_10025_),
    .B1_N(_10021_),
    .Y(_10029_));
 sky130_fd_sc_hd__nand3_2 _31663_ (.A(_10019_),
    .B(_10020_),
    .C(_10021_),
    .Y(_10030_));
 sky130_fd_sc_hd__nand3_2 _31664_ (.A(_10029_),
    .B(_10027_),
    .C(_10030_),
    .Y(_10031_));
 sky130_fd_sc_hd__nand2_2 _31665_ (.A(_10028_),
    .B(_10031_),
    .Y(_10032_));
 sky130_fd_sc_hd__o21bai_2 _31666_ (.A1(_09736_),
    .A2(_09739_),
    .B1_N(_09734_),
    .Y(_10033_));
 sky130_fd_sc_hd__a21oi_2 _31667_ (.A1(_09752_),
    .A2(_10033_),
    .B1(_09740_),
    .Y(_10034_));
 sky130_fd_sc_hd__xor2_2 _31668_ (.A(_10032_),
    .B(_10034_),
    .X(_02648_));
 sky130_fd_sc_hd__nand2_2 _31669_ (.A(_05926_),
    .B(_09511_),
    .Y(_10035_));
 sky130_fd_sc_hd__nand2_2 _31670_ (.A(_05929_),
    .B(_09808_),
    .Y(_10036_));
 sky130_fd_sc_hd__nor2_2 _31671_ (.A(_10035_),
    .B(_10036_),
    .Y(_10037_));
 sky130_fd_sc_hd__nand2_2 _31672_ (.A(_10035_),
    .B(_10036_),
    .Y(_10038_));
 sky130_fd_sc_hd__buf_1 _31673_ (.A(\pcpi_mul.rs1[30] ),
    .X(_10039_));
 sky130_fd_sc_hd__and2_2 _31674_ (.A(_05820_),
    .B(_10039_),
    .X(_10040_));
 sky130_fd_sc_hd__nand3b_2 _31675_ (.A_N(_10037_),
    .B(_10038_),
    .C(_10040_),
    .Y(_10041_));
 sky130_fd_sc_hd__buf_1 _31676_ (.A(_19161_),
    .X(_10042_));
 sky130_fd_sc_hd__buf_1 _31677_ (.A(_10042_),
    .X(_10043_));
 sky130_fd_sc_hd__a22oi_2 _31678_ (.A1(_18845_),
    .A2(_09787_),
    .B1(_05464_),
    .B2(_10043_),
    .Y(_10044_));
 sky130_fd_sc_hd__o21bai_2 _31679_ (.A1(_10044_),
    .A2(_10037_),
    .B1_N(_10040_),
    .Y(_10045_));
 sky130_fd_sc_hd__a21oi_2 _31680_ (.A1(_09796_),
    .A2(_09794_),
    .B1(_09792_),
    .Y(_10046_));
 sky130_fd_sc_hd__a21bo_2 _31681_ (.A1(_10041_),
    .A2(_10045_),
    .B1_N(_10046_),
    .X(_10047_));
 sky130_fd_sc_hd__nand3b_2 _31682_ (.A_N(_10046_),
    .B(_10045_),
    .C(_10041_),
    .Y(_10048_));
 sky130_fd_sc_hd__nand2_2 _31683_ (.A(_05835_),
    .B(_09805_),
    .Y(_10049_));
 sky130_fd_sc_hd__nand2_2 _31684_ (.A(_05956_),
    .B(_09793_),
    .Y(_10050_));
 sky130_fd_sc_hd__xor2_2 _31685_ (.A(_10049_),
    .B(_10050_),
    .X(_10051_));
 sky130_fd_sc_hd__buf_1 _31686_ (.A(_09802_),
    .X(_10052_));
 sky130_fd_sc_hd__and2_2 _31687_ (.A(_07121_),
    .B(_10052_),
    .X(_10053_));
 sky130_fd_sc_hd__nand2_2 _31688_ (.A(_10051_),
    .B(_10053_),
    .Y(_10054_));
 sky130_fd_sc_hd__xnor2_2 _31689_ (.A(_10049_),
    .B(_10050_),
    .Y(_10055_));
 sky130_fd_sc_hd__o21ai_2 _31690_ (.A1(_06923_),
    .A2(_19159_),
    .B1(_10055_),
    .Y(_10056_));
 sky130_fd_sc_hd__nand2_2 _31691_ (.A(_10054_),
    .B(_10056_),
    .Y(_10057_));
 sky130_fd_sc_hd__a21boi_2 _31692_ (.A1(_10047_),
    .A2(_10048_),
    .B1_N(_10057_),
    .Y(_10058_));
 sky130_fd_sc_hd__nand3b_2 _31693_ (.A_N(_10057_),
    .B(_10048_),
    .C(_10047_),
    .Y(_10059_));
 sky130_vsdinv _31694_ (.A(_10059_),
    .Y(_10060_));
 sky130_fd_sc_hd__a21oi_2 _31695_ (.A1(_09795_),
    .A2(_09797_),
    .B1(_09798_),
    .Y(_10061_));
 sky130_fd_sc_hd__o21ai_2 _31696_ (.A1(_09814_),
    .A2(_10061_),
    .B1(_09800_),
    .Y(_10062_));
 sky130_fd_sc_hd__o21bai_2 _31697_ (.A1(_10058_),
    .A2(_10060_),
    .B1_N(_10062_),
    .Y(_10063_));
 sky130_fd_sc_hd__o21a_2 _31698_ (.A1(_09803_),
    .A2(_09806_),
    .B1(_09811_),
    .X(_10064_));
 sky130_vsdinv _31699_ (.A(_10064_),
    .Y(_10065_));
 sky130_fd_sc_hd__nand3b_2 _31700_ (.A_N(_10058_),
    .B(_10059_),
    .C(_10062_),
    .Y(_10066_));
 sky130_fd_sc_hd__nand3_2 _31701_ (.A(_10063_),
    .B(_10065_),
    .C(_10066_),
    .Y(_10067_));
 sky130_vsdinv _31702_ (.A(_10067_),
    .Y(_10068_));
 sky130_fd_sc_hd__a21oi_2 _31703_ (.A1(_10063_),
    .A2(_10066_),
    .B1(_10065_),
    .Y(_10069_));
 sky130_fd_sc_hd__buf_1 _31704_ (.A(_09072_),
    .X(_10070_));
 sky130_fd_sc_hd__a22oi_2 _31705_ (.A1(_05870_),
    .A2(_10070_),
    .B1(_06097_),
    .B2(_09089_),
    .Y(_10071_));
 sky130_fd_sc_hd__nand2_2 _31706_ (.A(_07059_),
    .B(_09072_),
    .Y(_10072_));
 sky130_fd_sc_hd__nand2_2 _31707_ (.A(_18833_),
    .B(_09492_),
    .Y(_10073_));
 sky130_fd_sc_hd__nor2_2 _31708_ (.A(_10072_),
    .B(_10073_),
    .Y(_10074_));
 sky130_fd_sc_hd__and2_2 _31709_ (.A(_05778_),
    .B(_19172_),
    .X(_10075_));
 sky130_fd_sc_hd__o21bai_2 _31710_ (.A1(_10071_),
    .A2(_10074_),
    .B1_N(_10075_),
    .Y(_10076_));
 sky130_fd_sc_hd__buf_1 _31711_ (.A(_09495_),
    .X(_10077_));
 sky130_fd_sc_hd__nand3b_2 _31712_ (.A_N(_10072_),
    .B(_06227_),
    .C(_10077_),
    .Y(_10078_));
 sky130_fd_sc_hd__nand2_2 _31713_ (.A(_10072_),
    .B(_10073_),
    .Y(_10079_));
 sky130_fd_sc_hd__nand3_2 _31714_ (.A(_10078_),
    .B(_10079_),
    .C(_10075_),
    .Y(_10080_));
 sky130_fd_sc_hd__nand2_2 _31715_ (.A(_10076_),
    .B(_10080_),
    .Y(_10081_));
 sky130_fd_sc_hd__a21oi_2 _31716_ (.A1(_09877_),
    .A2(_09881_),
    .B1(_09878_),
    .Y(_10082_));
 sky130_fd_sc_hd__nand2_2 _31717_ (.A(_10081_),
    .B(_10082_),
    .Y(_10083_));
 sky130_fd_sc_hd__nand3b_2 _31718_ (.A_N(_10082_),
    .B(_10076_),
    .C(_10080_),
    .Y(_10084_));
 sky130_fd_sc_hd__nand2_2 _31719_ (.A(_10083_),
    .B(_10084_),
    .Y(_10085_));
 sky130_fd_sc_hd__o31a_2 _31720_ (.A1(_07920_),
    .A2(_09092_),
    .A3(_09753_),
    .B1(_09760_),
    .X(_10086_));
 sky130_fd_sc_hd__nand2_2 _31721_ (.A(_10085_),
    .B(_10086_),
    .Y(_10087_));
 sky130_vsdinv _31722_ (.A(_10086_),
    .Y(_10088_));
 sky130_fd_sc_hd__nand3_2 _31723_ (.A(_10083_),
    .B(_10088_),
    .C(_10084_),
    .Y(_10089_));
 sky130_fd_sc_hd__nand2_2 _31724_ (.A(_10087_),
    .B(_10089_),
    .Y(_10090_));
 sky130_fd_sc_hd__o21a_2 _31725_ (.A1(_09883_),
    .A2(_09874_),
    .B1(_09885_),
    .X(_10091_));
 sky130_fd_sc_hd__nand2_2 _31726_ (.A(_10090_),
    .B(_10091_),
    .Y(_10092_));
 sky130_fd_sc_hd__o21ai_2 _31727_ (.A1(_09883_),
    .A2(_09874_),
    .B1(_09885_),
    .Y(_10093_));
 sky130_fd_sc_hd__nand3_2 _31728_ (.A(_10093_),
    .B(_10087_),
    .C(_10089_),
    .Y(_10094_));
 sky130_fd_sc_hd__nand2_2 _31729_ (.A(_10092_),
    .B(_10094_),
    .Y(_10095_));
 sky130_fd_sc_hd__a21boi_2 _31730_ (.A1(_09764_),
    .A2(_09767_),
    .B1_N(_09765_),
    .Y(_10096_));
 sky130_fd_sc_hd__nand2_2 _31731_ (.A(_10095_),
    .B(_10096_),
    .Y(_10097_));
 sky130_vsdinv _31732_ (.A(_10096_),
    .Y(_10098_));
 sky130_fd_sc_hd__nand3_2 _31733_ (.A(_10092_),
    .B(_10098_),
    .C(_10094_),
    .Y(_10099_));
 sky130_fd_sc_hd__a21oi_2 _31734_ (.A1(_09774_),
    .A2(_09769_),
    .B1(_09771_),
    .Y(_10100_));
 sky130_fd_sc_hd__o21ai_2 _31735_ (.A1(_09777_),
    .A2(_10100_),
    .B1(_09775_),
    .Y(_10101_));
 sky130_fd_sc_hd__a21oi_2 _31736_ (.A1(_10097_),
    .A2(_10099_),
    .B1(_10101_),
    .Y(_10102_));
 sky130_fd_sc_hd__nand3_2 _31737_ (.A(_10097_),
    .B(_10099_),
    .C(_10101_),
    .Y(_10103_));
 sky130_vsdinv _31738_ (.A(_10103_),
    .Y(_10104_));
 sky130_fd_sc_hd__o22ai_2 _31739_ (.A1(_10068_),
    .A2(_10069_),
    .B1(_10102_),
    .B2(_10104_),
    .Y(_10105_));
 sky130_fd_sc_hd__nor2_2 _31740_ (.A(_10069_),
    .B(_10068_),
    .Y(_10106_));
 sky130_fd_sc_hd__a21o_2 _31741_ (.A1(_10097_),
    .A2(_10099_),
    .B1(_10101_),
    .X(_10107_));
 sky130_fd_sc_hd__nand3_2 _31742_ (.A(_10106_),
    .B(_10103_),
    .C(_10107_),
    .Y(_10108_));
 sky130_fd_sc_hd__a21oi_2 _31743_ (.A1(_09898_),
    .A2(_09899_),
    .B1(_09896_),
    .Y(_10109_));
 sky130_fd_sc_hd__o21ai_2 _31744_ (.A1(_09902_),
    .A2(_10109_),
    .B1(_09900_),
    .Y(_10110_));
 sky130_fd_sc_hd__a21oi_2 _31745_ (.A1(_10105_),
    .A2(_10108_),
    .B1(_10110_),
    .Y(_10111_));
 sky130_fd_sc_hd__nand3_2 _31746_ (.A(_10105_),
    .B(_10110_),
    .C(_10108_),
    .Y(_10112_));
 sky130_vsdinv _31747_ (.A(_10112_),
    .Y(_10113_));
 sky130_fd_sc_hd__o21a_2 _31748_ (.A1(_09825_),
    .A2(_09784_),
    .B1(_09783_),
    .X(_10114_));
 sky130_fd_sc_hd__buf_1 _31749_ (.A(_10114_),
    .X(_10115_));
 sky130_fd_sc_hd__o21ai_2 _31750_ (.A1(_10111_),
    .A2(_10113_),
    .B1(_10115_),
    .Y(_10116_));
 sky130_fd_sc_hd__a21o_2 _31751_ (.A1(_10105_),
    .A2(_10108_),
    .B1(_10110_),
    .X(_10117_));
 sky130_fd_sc_hd__buf_1 _31752_ (.A(_10112_),
    .X(_10118_));
 sky130_fd_sc_hd__nand3b_2 _31753_ (.A_N(_10114_),
    .B(_10117_),
    .C(_10118_),
    .Y(_10119_));
 sky130_fd_sc_hd__buf_1 _31754_ (.A(_07165_),
    .X(_10120_));
 sky130_fd_sc_hd__a22oi_2 _31755_ (.A1(_10120_),
    .A2(_07557_),
    .B1(_07395_),
    .B2(_07699_),
    .Y(_10121_));
 sky130_fd_sc_hd__nand2_2 _31756_ (.A(_07468_),
    .B(_07690_),
    .Y(_10122_));
 sky130_fd_sc_hd__nand2_2 _31757_ (.A(_07004_),
    .B(_07688_),
    .Y(_10123_));
 sky130_fd_sc_hd__nor2_2 _31758_ (.A(_10122_),
    .B(_10123_),
    .Y(_10124_));
 sky130_fd_sc_hd__and2_2 _31759_ (.A(_07012_),
    .B(_07694_),
    .X(_10125_));
 sky130_fd_sc_hd__o21bai_2 _31760_ (.A1(_10121_),
    .A2(_10124_),
    .B1_N(_10125_),
    .Y(_10126_));
 sky130_fd_sc_hd__nand3b_2 _31761_ (.A_N(_10122_),
    .B(_07480_),
    .C(_07314_),
    .Y(_10127_));
 sky130_fd_sc_hd__nand2_2 _31762_ (.A(_10122_),
    .B(_10123_),
    .Y(_10128_));
 sky130_fd_sc_hd__nand3_2 _31763_ (.A(_10127_),
    .B(_10125_),
    .C(_10128_),
    .Y(_10129_));
 sky130_fd_sc_hd__nand2_2 _31764_ (.A(_10126_),
    .B(_10129_),
    .Y(_10130_));
 sky130_fd_sc_hd__a21oi_2 _31765_ (.A1(_09909_),
    .A2(_09908_),
    .B1(_09907_),
    .Y(_10131_));
 sky130_fd_sc_hd__nand2_2 _31766_ (.A(_10130_),
    .B(_10131_),
    .Y(_10132_));
 sky130_fd_sc_hd__nand3b_2 _31767_ (.A_N(_10131_),
    .B(_10129_),
    .C(_10126_),
    .Y(_10133_));
 sky130_fd_sc_hd__nand2_2 _31768_ (.A(_10132_),
    .B(_10133_),
    .Y(_10134_));
 sky130_fd_sc_hd__o31a_2 _31769_ (.A1(_07178_),
    .A2(_19233_),
    .A3(_09840_),
    .B1(_09846_),
    .X(_10135_));
 sky130_fd_sc_hd__nand2_2 _31770_ (.A(_10134_),
    .B(_10135_),
    .Y(_10136_));
 sky130_fd_sc_hd__nand3b_2 _31771_ (.A_N(_10135_),
    .B(_10132_),
    .C(_10133_),
    .Y(_10137_));
 sky130_fd_sc_hd__nand2_2 _31772_ (.A(_10136_),
    .B(_10137_),
    .Y(_10138_));
 sky130_fd_sc_hd__a21boi_2 _31773_ (.A1(_09850_),
    .A2(_09854_),
    .B1_N(_09852_),
    .Y(_10139_));
 sky130_fd_sc_hd__nand2_2 _31774_ (.A(_10138_),
    .B(_10139_),
    .Y(_10140_));
 sky130_fd_sc_hd__nand2_2 _31775_ (.A(_09856_),
    .B(_09852_),
    .Y(_10141_));
 sky130_fd_sc_hd__nand3_2 _31776_ (.A(_10141_),
    .B(_10137_),
    .C(_10136_),
    .Y(_10142_));
 sky130_fd_sc_hd__buf_1 _31777_ (.A(_10142_),
    .X(_10143_));
 sky130_fd_sc_hd__nand2_2 _31778_ (.A(_07495_),
    .B(_06734_),
    .Y(_10144_));
 sky130_fd_sc_hd__nand2_2 _31779_ (.A(_06392_),
    .B(_07605_),
    .Y(_10145_));
 sky130_fd_sc_hd__nor2_2 _31780_ (.A(_10144_),
    .B(_10145_),
    .Y(_10146_));
 sky130_fd_sc_hd__and2_2 _31781_ (.A(_07195_),
    .B(_08299_),
    .X(_10147_));
 sky130_fd_sc_hd__nand2_2 _31782_ (.A(_10144_),
    .B(_10145_),
    .Y(_10148_));
 sky130_fd_sc_hd__nand3b_2 _31783_ (.A_N(_10146_),
    .B(_10147_),
    .C(_10148_),
    .Y(_10149_));
 sky130_fd_sc_hd__buf_1 _31784_ (.A(_07115_),
    .X(_10150_));
 sky130_fd_sc_hd__a22oi_2 _31785_ (.A1(_07503_),
    .A2(_10150_),
    .B1(_08688_),
    .B2(_07118_),
    .Y(_10151_));
 sky130_fd_sc_hd__o21bai_2 _31786_ (.A1(_10151_),
    .A2(_10146_),
    .B1_N(_10147_),
    .Y(_10152_));
 sky130_fd_sc_hd__nand2_2 _31787_ (.A(_10149_),
    .B(_10152_),
    .Y(_10153_));
 sky130_fd_sc_hd__a21oi_2 _31788_ (.A1(_09868_),
    .A2(_09867_),
    .B1(_09866_),
    .Y(_10154_));
 sky130_fd_sc_hd__nand2_2 _31789_ (.A(_10153_),
    .B(_10154_),
    .Y(_10155_));
 sky130_fd_sc_hd__nand3b_2 _31790_ (.A_N(_10154_),
    .B(_10149_),
    .C(_10152_),
    .Y(_10156_));
 sky130_fd_sc_hd__nand2_2 _31791_ (.A(_10155_),
    .B(_10156_),
    .Y(_10157_));
 sky130_fd_sc_hd__nand2_2 _31792_ (.A(_06670_),
    .B(_08302_),
    .Y(_10158_));
 sky130_fd_sc_hd__buf_1 _31793_ (.A(_19195_),
    .X(_10159_));
 sky130_fd_sc_hd__nand2_2 _31794_ (.A(_18819_),
    .B(_10159_),
    .Y(_10160_));
 sky130_fd_sc_hd__nand2_2 _31795_ (.A(_10158_),
    .B(_10160_),
    .Y(_10161_));
 sky130_fd_sc_hd__buf_1 _31796_ (.A(_19196_),
    .X(_10162_));
 sky130_fd_sc_hd__nand3b_2 _31797_ (.A_N(_10158_),
    .B(_06268_),
    .C(_10162_),
    .Y(_10163_));
 sky130_fd_sc_hd__o2bb2ai_2 _31798_ (.A1_N(_10161_),
    .A2_N(_10163_),
    .B1(_18824_),
    .B2(_19192_),
    .Y(_10164_));
 sky130_fd_sc_hd__and2_2 _31799_ (.A(_05895_),
    .B(_07963_),
    .X(_10165_));
 sky130_fd_sc_hd__nand3_2 _31800_ (.A(_10163_),
    .B(_10165_),
    .C(_10161_),
    .Y(_10166_));
 sky130_fd_sc_hd__nand2_2 _31801_ (.A(_10164_),
    .B(_10166_),
    .Y(_10167_));
 sky130_fd_sc_hd__nand2_2 _31802_ (.A(_10157_),
    .B(_10167_),
    .Y(_10168_));
 sky130_fd_sc_hd__nand3b_2 _31803_ (.A_N(_10167_),
    .B(_10155_),
    .C(_10156_),
    .Y(_10169_));
 sky130_fd_sc_hd__nand2_2 _31804_ (.A(_10168_),
    .B(_10169_),
    .Y(_10170_));
 sky130_vsdinv _31805_ (.A(_10170_),
    .Y(_10171_));
 sky130_fd_sc_hd__a21oi_2 _31806_ (.A1(_10140_),
    .A2(_10143_),
    .B1(_10171_),
    .Y(_10172_));
 sky130_fd_sc_hd__a21oi_2 _31807_ (.A1(_10136_),
    .A2(_10137_),
    .B1(_10141_),
    .Y(_10173_));
 sky130_fd_sc_hd__nor3b_2 _31808_ (.A(_10170_),
    .B(_10173_),
    .C_N(_10143_),
    .Y(_10174_));
 sky130_fd_sc_hd__a21boi_2 _31809_ (.A1(_09932_),
    .A2(_09937_),
    .B1_N(_09933_),
    .Y(_10175_));
 sky130_fd_sc_hd__o21ai_2 _31810_ (.A1(_10172_),
    .A2(_10174_),
    .B1(_10175_),
    .Y(_10176_));
 sky130_fd_sc_hd__nand2_2 _31811_ (.A(_09938_),
    .B(_09933_),
    .Y(_10177_));
 sky130_fd_sc_hd__a21o_2 _31812_ (.A1(_10140_),
    .A2(_10142_),
    .B1(_10171_),
    .X(_10178_));
 sky130_fd_sc_hd__nand3_2 _31813_ (.A(_10171_),
    .B(_10140_),
    .C(_10143_),
    .Y(_10179_));
 sky130_fd_sc_hd__nand3_2 _31814_ (.A(_10177_),
    .B(_10178_),
    .C(_10179_),
    .Y(_10180_));
 sky130_fd_sc_hd__nand2_2 _31815_ (.A(_10176_),
    .B(_10180_),
    .Y(_10181_));
 sky130_fd_sc_hd__o21a_2 _31816_ (.A1(_09890_),
    .A2(_09892_),
    .B1(_09863_),
    .X(_10182_));
 sky130_fd_sc_hd__nand2_2 _31817_ (.A(_10181_),
    .B(_10182_),
    .Y(_10183_));
 sky130_vsdinv _31818_ (.A(_10182_),
    .Y(_10184_));
 sky130_fd_sc_hd__nand3_2 _31819_ (.A(_10176_),
    .B(_10184_),
    .C(_10180_),
    .Y(_10185_));
 sky130_fd_sc_hd__buf_1 _31820_ (.A(_08462_),
    .X(_10186_));
 sky130_fd_sc_hd__a22oi_2 _31821_ (.A1(_10186_),
    .A2(_05963_),
    .B1(_09263_),
    .B2(_07499_),
    .Y(_10187_));
 sky130_fd_sc_hd__nand2_2 _31822_ (.A(_08462_),
    .B(_05648_),
    .Y(_10188_));
 sky130_fd_sc_hd__nand2_2 _31823_ (.A(_08971_),
    .B(_19261_),
    .Y(_10189_));
 sky130_fd_sc_hd__nor2_2 _31824_ (.A(_10188_),
    .B(_10189_),
    .Y(_10190_));
 sky130_fd_sc_hd__and2_2 _31825_ (.A(_08234_),
    .B(_19257_),
    .X(_10191_));
 sky130_fd_sc_hd__o21bai_2 _31826_ (.A1(_10187_),
    .A2(_10190_),
    .B1_N(_10191_),
    .Y(_10192_));
 sky130_fd_sc_hd__nand3b_2 _31827_ (.A_N(_10188_),
    .B(_18753_),
    .C(_05728_),
    .Y(_10193_));
 sky130_fd_sc_hd__nand2_2 _31828_ (.A(_10188_),
    .B(_10189_),
    .Y(_10194_));
 sky130_fd_sc_hd__nand3_2 _31829_ (.A(_10193_),
    .B(_10191_),
    .C(_10194_),
    .Y(_10195_));
 sky130_fd_sc_hd__nand2_2 _31830_ (.A(_10192_),
    .B(_10195_),
    .Y(_10196_));
 sky130_fd_sc_hd__o21ai_2 _31831_ (.A1(_09917_),
    .A2(_09913_),
    .B1(_09920_),
    .Y(_10197_));
 sky130_vsdinv _31832_ (.A(_10197_),
    .Y(_10198_));
 sky130_fd_sc_hd__nand2_2 _31833_ (.A(_10196_),
    .B(_10198_),
    .Y(_10199_));
 sky130_fd_sc_hd__nand3_2 _31834_ (.A(_10192_),
    .B(_10195_),
    .C(_10197_),
    .Y(_10200_));
 sky130_fd_sc_hd__nand2_2 _31835_ (.A(_08217_),
    .B(_19252_),
    .Y(_10201_));
 sky130_fd_sc_hd__nand2_2 _31836_ (.A(_08985_),
    .B(_08905_),
    .Y(_10202_));
 sky130_fd_sc_hd__nor2_2 _31837_ (.A(_10201_),
    .B(_10202_),
    .Y(_10203_));
 sky130_fd_sc_hd__and2_2 _31838_ (.A(_07532_),
    .B(_19242_),
    .X(_10204_));
 sky130_fd_sc_hd__nand2_2 _31839_ (.A(_10201_),
    .B(_10202_),
    .Y(_10205_));
 sky130_fd_sc_hd__nand3b_2 _31840_ (.A_N(_10203_),
    .B(_10204_),
    .C(_10205_),
    .Y(_10206_));
 sky130_fd_sc_hd__buf_1 _31841_ (.A(_08985_),
    .X(_10207_));
 sky130_fd_sc_hd__a22oi_2 _31842_ (.A1(_07851_),
    .A2(_09340_),
    .B1(_10207_),
    .B2(_09341_),
    .Y(_10208_));
 sky130_fd_sc_hd__o21bai_2 _31843_ (.A1(_10208_),
    .A2(_10203_),
    .B1_N(_10204_),
    .Y(_10209_));
 sky130_fd_sc_hd__nand2_2 _31844_ (.A(_10206_),
    .B(_10209_),
    .Y(_10210_));
 sky130_vsdinv _31845_ (.A(_10210_),
    .Y(_10211_));
 sky130_fd_sc_hd__a21oi_2 _31846_ (.A1(_10199_),
    .A2(_10200_),
    .B1(_10211_),
    .Y(_10212_));
 sky130_fd_sc_hd__a21oi_2 _31847_ (.A1(_10192_),
    .A2(_10195_),
    .B1(_10197_),
    .Y(_10213_));
 sky130_vsdinv _31848_ (.A(_10200_),
    .Y(_10214_));
 sky130_fd_sc_hd__nor3_2 _31849_ (.A(_10210_),
    .B(_10213_),
    .C(_10214_),
    .Y(_10215_));
 sky130_fd_sc_hd__a21oi_2 _31850_ (.A1(_09943_),
    .A2(_09946_),
    .B1(_09948_),
    .Y(_10216_));
 sky130_fd_sc_hd__o21ai_2 _31851_ (.A1(_09952_),
    .A2(_10216_),
    .B1(_09951_),
    .Y(_10217_));
 sky130_fd_sc_hd__o21bai_2 _31852_ (.A1(_10212_),
    .A2(_10215_),
    .B1_N(_10217_),
    .Y(_10218_));
 sky130_fd_sc_hd__o21ai_2 _31853_ (.A1(_10213_),
    .A2(_10214_),
    .B1(_10210_),
    .Y(_10219_));
 sky130_fd_sc_hd__nand3_2 _31854_ (.A(_10211_),
    .B(_10199_),
    .C(_10200_),
    .Y(_10220_));
 sky130_fd_sc_hd__nand3_2 _31855_ (.A(_10219_),
    .B(_10217_),
    .C(_10220_),
    .Y(_10221_));
 sky130_fd_sc_hd__nand2_2 _31856_ (.A(_10218_),
    .B(_10221_),
    .Y(_10222_));
 sky130_fd_sc_hd__a21oi_2 _31857_ (.A1(_09928_),
    .A2(_09929_),
    .B1(_09926_),
    .Y(_10223_));
 sky130_fd_sc_hd__nand2_2 _31858_ (.A(_10222_),
    .B(_10223_),
    .Y(_10224_));
 sky130_vsdinv _31859_ (.A(_10223_),
    .Y(_10225_));
 sky130_fd_sc_hd__nand3_2 _31860_ (.A(_10218_),
    .B(_10225_),
    .C(_10221_),
    .Y(_10226_));
 sky130_fd_sc_hd__buf_1 _31861_ (.A(_10226_),
    .X(_10227_));
 sky130_fd_sc_hd__a22oi_2 _31862_ (.A1(_09312_),
    .A2(_07403_),
    .B1(_09313_),
    .B2(_05746_),
    .Y(_10228_));
 sky130_fd_sc_hd__buf_1 _31863_ (.A(_09005_),
    .X(_10229_));
 sky130_fd_sc_hd__nand2_2 _31864_ (.A(_10229_),
    .B(_07794_),
    .Y(_10230_));
 sky130_fd_sc_hd__buf_1 _31865_ (.A(_08754_),
    .X(_10231_));
 sky130_fd_sc_hd__nand2_2 _31866_ (.A(_10231_),
    .B(_05518_),
    .Y(_10232_));
 sky130_fd_sc_hd__nor2_2 _31867_ (.A(_10230_),
    .B(_10232_),
    .Y(_10233_));
 sky130_fd_sc_hd__and2_2 _31868_ (.A(_08758_),
    .B(_19272_),
    .X(_10234_));
 sky130_fd_sc_hd__o21bai_2 _31869_ (.A1(_10228_),
    .A2(_10233_),
    .B1_N(_10234_),
    .Y(_10235_));
 sky130_fd_sc_hd__nand3b_2 _31870_ (.A_N(_10230_),
    .B(_08756_),
    .C(_05746_),
    .Y(_10236_));
 sky130_fd_sc_hd__nand2_2 _31871_ (.A(_10230_),
    .B(_10232_),
    .Y(_10237_));
 sky130_fd_sc_hd__nand3_2 _31872_ (.A(_10236_),
    .B(_10234_),
    .C(_10237_),
    .Y(_10238_));
 sky130_fd_sc_hd__nand2_2 _31873_ (.A(_10235_),
    .B(_10238_),
    .Y(_10239_));
 sky130_fd_sc_hd__nand2_2 _31874_ (.A(_09956_),
    .B(_09959_),
    .Y(_10240_));
 sky130_fd_sc_hd__nor2_2 _31875_ (.A(_09956_),
    .B(_09959_),
    .Y(_10241_));
 sky130_fd_sc_hd__a21oi_2 _31876_ (.A1(_10240_),
    .A2(_09955_),
    .B1(_10241_),
    .Y(_10242_));
 sky130_fd_sc_hd__nand2_2 _31877_ (.A(_10239_),
    .B(_10242_),
    .Y(_10243_));
 sky130_fd_sc_hd__nand3b_2 _31878_ (.A_N(_10242_),
    .B(_10238_),
    .C(_10235_),
    .Y(_10244_));
 sky130_fd_sc_hd__buf_1 _31879_ (.A(_18740_),
    .X(_10245_));
 sky130_fd_sc_hd__buf_1 _31880_ (.A(_10245_),
    .X(_10246_));
 sky130_fd_sc_hd__o31ai_2 _31881_ (.A1(_10246_),
    .A2(_19279_),
    .A3(_09940_),
    .B1(_09945_),
    .Y(_10247_));
 sky130_fd_sc_hd__a21oi_2 _31882_ (.A1(_10243_),
    .A2(_10244_),
    .B1(_10247_),
    .Y(_10248_));
 sky130_fd_sc_hd__nand3_2 _31883_ (.A(_10243_),
    .B(_10247_),
    .C(_10244_),
    .Y(_10249_));
 sky130_vsdinv _31884_ (.A(_10249_),
    .Y(_10250_));
 sky130_fd_sc_hd__nand2_2 _31885_ (.A(_09958_),
    .B(_19297_),
    .Y(_10251_));
 sky130_fd_sc_hd__buf_1 _31886_ (.A(\pcpi_mul.rs2[28] ),
    .X(_10252_));
 sky130_fd_sc_hd__buf_1 _31887_ (.A(_10252_),
    .X(_10253_));
 sky130_fd_sc_hd__nand2_2 _31888_ (.A(_10253_),
    .B(_07013_),
    .Y(_10254_));
 sky130_fd_sc_hd__nor2_2 _31889_ (.A(_10251_),
    .B(_10254_),
    .Y(_10255_));
 sky130_fd_sc_hd__and2_2 _31890_ (.A(_18723_),
    .B(_05644_),
    .X(_10256_));
 sky130_fd_sc_hd__nand2_2 _31891_ (.A(_10251_),
    .B(_10254_),
    .Y(_10257_));
 sky130_fd_sc_hd__nand3b_2 _31892_ (.A_N(_10255_),
    .B(_10256_),
    .C(_10257_),
    .Y(_10258_));
 sky130_fd_sc_hd__buf_1 _31893_ (.A(\pcpi_mul.rs2[29] ),
    .X(_10259_));
 sky130_fd_sc_hd__buf_1 _31894_ (.A(_10259_),
    .X(_10260_));
 sky130_fd_sc_hd__buf_1 _31895_ (.A(_10260_),
    .X(_10261_));
 sky130_fd_sc_hd__buf_1 _31896_ (.A(_10252_),
    .X(_10262_));
 sky130_fd_sc_hd__buf_1 _31897_ (.A(_10262_),
    .X(_10263_));
 sky130_fd_sc_hd__a22oi_2 _31898_ (.A1(_10261_),
    .A2(_05402_),
    .B1(_10263_),
    .B2(_05494_),
    .Y(_10264_));
 sky130_fd_sc_hd__o21bai_2 _31899_ (.A1(_10264_),
    .A2(_10255_),
    .B1_N(_10256_),
    .Y(_10265_));
 sky130_fd_sc_hd__buf_1 _31900_ (.A(\pcpi_mul.rs2[30] ),
    .X(_10266_));
 sky130_fd_sc_hd__buf_1 _31901_ (.A(_10266_),
    .X(_10267_));
 sky130_fd_sc_hd__buf_1 _31902_ (.A(_10267_),
    .X(_10268_));
 sky130_fd_sc_hd__and2_2 _31903_ (.A(_10268_),
    .B(_05239_),
    .X(_10269_));
 sky130_fd_sc_hd__a21oi_2 _31904_ (.A1(_10258_),
    .A2(_10265_),
    .B1(_10269_),
    .Y(_10270_));
 sky130_fd_sc_hd__nand3_2 _31905_ (.A(_10258_),
    .B(_10265_),
    .C(_10269_),
    .Y(_10271_));
 sky130_vsdinv _31906_ (.A(_10271_),
    .Y(_10272_));
 sky130_fd_sc_hd__nor2_2 _31907_ (.A(_10270_),
    .B(_10272_),
    .Y(_10273_));
 sky130_fd_sc_hd__o21bai_2 _31908_ (.A1(_10248_),
    .A2(_10250_),
    .B1_N(_10273_),
    .Y(_10274_));
 sky130_fd_sc_hd__a21o_2 _31909_ (.A1(_10243_),
    .A2(_10244_),
    .B1(_10247_),
    .X(_10275_));
 sky130_fd_sc_hd__nand3_2 _31910_ (.A(_10275_),
    .B(_10273_),
    .C(_10249_),
    .Y(_10276_));
 sky130_fd_sc_hd__nand3b_2 _31911_ (.A_N(_09964_),
    .B(_10274_),
    .C(_10276_),
    .Y(_10277_));
 sky130_fd_sc_hd__nand2_2 _31912_ (.A(_10274_),
    .B(_10276_),
    .Y(_10278_));
 sky130_fd_sc_hd__nand2_2 _31913_ (.A(_10278_),
    .B(_09964_),
    .Y(_10279_));
 sky130_fd_sc_hd__a22oi_2 _31914_ (.A1(_10224_),
    .A2(_10227_),
    .B1(_10277_),
    .B2(_10279_),
    .Y(_10280_));
 sky130_fd_sc_hd__nand2_2 _31915_ (.A(_10224_),
    .B(_10227_),
    .Y(_10281_));
 sky130_fd_sc_hd__nand2_2 _31916_ (.A(_10279_),
    .B(_10277_),
    .Y(_10282_));
 sky130_fd_sc_hd__nor2_2 _31917_ (.A(_10281_),
    .B(_10282_),
    .Y(_10283_));
 sky130_fd_sc_hd__a31oi_2 _31918_ (.A1(_09968_),
    .A2(_09936_),
    .A3(_09939_),
    .B1(_09977_),
    .Y(_10284_));
 sky130_fd_sc_hd__o21ai_2 _31919_ (.A1(_10280_),
    .A2(_10283_),
    .B1(_10284_),
    .Y(_10285_));
 sky130_fd_sc_hd__o21bai_2 _31920_ (.A1(_09976_),
    .A2(_09971_),
    .B1_N(_09977_),
    .Y(_10286_));
 sky130_fd_sc_hd__a21oi_2 _31921_ (.A1(_10218_),
    .A2(_10221_),
    .B1(_10225_),
    .Y(_10287_));
 sky130_vsdinv _31922_ (.A(_10227_),
    .Y(_10288_));
 sky130_fd_sc_hd__nor2_2 _31923_ (.A(_10287_),
    .B(_10288_),
    .Y(_10289_));
 sky130_fd_sc_hd__nand3_2 _31924_ (.A(_10289_),
    .B(_10277_),
    .C(_10279_),
    .Y(_10290_));
 sky130_fd_sc_hd__nand2_2 _31925_ (.A(_10282_),
    .B(_10281_),
    .Y(_10291_));
 sky130_fd_sc_hd__nand3_2 _31926_ (.A(_10286_),
    .B(_10290_),
    .C(_10291_),
    .Y(_10292_));
 sky130_fd_sc_hd__buf_1 _31927_ (.A(_10292_),
    .X(_10293_));
 sky130_fd_sc_hd__a22oi_2 _31928_ (.A1(_10183_),
    .A2(_10185_),
    .B1(_10285_),
    .B2(_10293_),
    .Y(_10294_));
 sky130_fd_sc_hd__nand2_2 _31929_ (.A(_10183_),
    .B(_10185_),
    .Y(_10295_));
 sky130_fd_sc_hd__nand2_2 _31930_ (.A(_10285_),
    .B(_10292_),
    .Y(_10296_));
 sky130_fd_sc_hd__nor2_2 _31931_ (.A(_10295_),
    .B(_10296_),
    .Y(_10297_));
 sky130_fd_sc_hd__a21oi_2 _31932_ (.A1(_09979_),
    .A2(_09980_),
    .B1(_09974_),
    .Y(_10298_));
 sky130_fd_sc_hd__o21a_2 _31933_ (.A1(_10298_),
    .A2(_09985_),
    .B1(_09982_),
    .X(_10299_));
 sky130_fd_sc_hd__o21ai_2 _31934_ (.A1(_10294_),
    .A2(_10297_),
    .B1(_10299_),
    .Y(_10300_));
 sky130_fd_sc_hd__o21ai_2 _31935_ (.A1(_10298_),
    .A2(_09985_),
    .B1(_09982_),
    .Y(_10301_));
 sky130_fd_sc_hd__a21oi_2 _31936_ (.A1(_10176_),
    .A2(_10180_),
    .B1(_10184_),
    .Y(_10302_));
 sky130_vsdinv _31937_ (.A(_10185_),
    .Y(_10303_));
 sky130_fd_sc_hd__nor2_2 _31938_ (.A(_10302_),
    .B(_10303_),
    .Y(_10304_));
 sky130_fd_sc_hd__nand3_2 _31939_ (.A(_10304_),
    .B(_10293_),
    .C(_10285_),
    .Y(_10305_));
 sky130_fd_sc_hd__nand2_2 _31940_ (.A(_10296_),
    .B(_10295_),
    .Y(_10306_));
 sky130_fd_sc_hd__nand3_2 _31941_ (.A(_10301_),
    .B(_10305_),
    .C(_10306_),
    .Y(_10307_));
 sky130_fd_sc_hd__buf_1 _31942_ (.A(_10307_),
    .X(_10308_));
 sky130_fd_sc_hd__a22oi_2 _31943_ (.A1(_10116_),
    .A2(_10119_),
    .B1(_10300_),
    .B2(_10308_),
    .Y(_10309_));
 sky130_fd_sc_hd__nand2_2 _31944_ (.A(_10116_),
    .B(_10119_),
    .Y(_10310_));
 sky130_fd_sc_hd__nand2_2 _31945_ (.A(_10300_),
    .B(_10307_),
    .Y(_10311_));
 sky130_fd_sc_hd__nor2_2 _31946_ (.A(_10310_),
    .B(_10311_),
    .Y(_10312_));
 sky130_fd_sc_hd__a21boi_2 _31947_ (.A1(_10005_),
    .A2(_09989_),
    .B1_N(_09994_),
    .Y(_10313_));
 sky130_fd_sc_hd__o21ai_2 _31948_ (.A1(_10309_),
    .A2(_10312_),
    .B1(_10313_),
    .Y(_10314_));
 sky130_fd_sc_hd__a21oi_2 _31949_ (.A1(_09990_),
    .A2(_09992_),
    .B1(_09991_),
    .Y(_10315_));
 sky130_fd_sc_hd__o21ai_2 _31950_ (.A1(_10315_),
    .A2(_09996_),
    .B1(_09994_),
    .Y(_10316_));
 sky130_fd_sc_hd__a21boi_2 _31951_ (.A1(_10117_),
    .A2(_10118_),
    .B1_N(_10115_),
    .Y(_10317_));
 sky130_fd_sc_hd__nor3_2 _31952_ (.A(_10115_),
    .B(_10111_),
    .C(_10113_),
    .Y(_10318_));
 sky130_fd_sc_hd__nor2_2 _31953_ (.A(_10317_),
    .B(_10318_),
    .Y(_10319_));
 sky130_fd_sc_hd__nand3_2 _31954_ (.A(_10319_),
    .B(_10308_),
    .C(_10300_),
    .Y(_10320_));
 sky130_fd_sc_hd__nand2_2 _31955_ (.A(_10311_),
    .B(_10310_),
    .Y(_10321_));
 sky130_fd_sc_hd__nand3_2 _31956_ (.A(_10316_),
    .B(_10320_),
    .C(_10321_),
    .Y(_10322_));
 sky130_fd_sc_hd__o21a_2 _31957_ (.A1(_09821_),
    .A2(_09818_),
    .B1(_09819_),
    .X(_10323_));
 sky130_fd_sc_hd__o21ai_2 _31958_ (.A1(_09833_),
    .A2(_09829_),
    .B1(_09838_),
    .Y(_10324_));
 sky130_fd_sc_hd__xnor2_2 _31959_ (.A(_10323_),
    .B(_10324_),
    .Y(_10325_));
 sky130_fd_sc_hd__a21oi_2 _31960_ (.A1(_10314_),
    .A2(_10322_),
    .B1(_10325_),
    .Y(_10326_));
 sky130_fd_sc_hd__nand3_2 _31961_ (.A(_10314_),
    .B(_10325_),
    .C(_10322_),
    .Y(_10327_));
 sky130_vsdinv _31962_ (.A(_10327_),
    .Y(_10328_));
 sky130_fd_sc_hd__a21oi_2 _31963_ (.A1(_10006_),
    .A2(_10007_),
    .B1(_10002_),
    .Y(_10329_));
 sky130_fd_sc_hd__o21ai_2 _31964_ (.A1(_10012_),
    .A2(_10329_),
    .B1(_10008_),
    .Y(_10330_));
 sky130_fd_sc_hd__o21bai_2 _31965_ (.A1(_10326_),
    .A2(_10328_),
    .B1_N(_10330_),
    .Y(_10331_));
 sky130_fd_sc_hd__nand2_2 _31966_ (.A(_10314_),
    .B(_10322_),
    .Y(_10332_));
 sky130_vsdinv _31967_ (.A(_10325_),
    .Y(_10333_));
 sky130_fd_sc_hd__nand2_2 _31968_ (.A(_10332_),
    .B(_10333_),
    .Y(_10334_));
 sky130_fd_sc_hd__nand3_2 _31969_ (.A(_10334_),
    .B(_10330_),
    .C(_10327_),
    .Y(_10335_));
 sky130_fd_sc_hd__a21oi_2 _31970_ (.A1(_09547_),
    .A2(_09545_),
    .B1(_10010_),
    .Y(_10336_));
 sky130_fd_sc_hd__buf_1 _31971_ (.A(_10336_),
    .X(_10337_));
 sky130_fd_sc_hd__a21oi_2 _31972_ (.A1(_10331_),
    .A2(_10335_),
    .B1(_10337_),
    .Y(_10338_));
 sky130_vsdinv _31973_ (.A(_10336_),
    .Y(_10339_));
 sky130_fd_sc_hd__a21oi_2 _31974_ (.A1(_10334_),
    .A2(_10327_),
    .B1(_10330_),
    .Y(_10340_));
 sky130_vsdinv _31975_ (.A(_10335_),
    .Y(_10341_));
 sky130_fd_sc_hd__nor3_2 _31976_ (.A(_10339_),
    .B(_10340_),
    .C(_10341_),
    .Y(_10342_));
 sky130_fd_sc_hd__o21ai_2 _31977_ (.A1(_10023_),
    .A2(_10024_),
    .B1(_10020_),
    .Y(_10343_));
 sky130_fd_sc_hd__o21bai_2 _31978_ (.A1(_10338_),
    .A2(_10342_),
    .B1_N(_10343_),
    .Y(_10344_));
 sky130_fd_sc_hd__o21bai_2 _31979_ (.A1(_10340_),
    .A2(_10341_),
    .B1_N(_10337_),
    .Y(_10345_));
 sky130_fd_sc_hd__nand3_2 _31980_ (.A(_10331_),
    .B(_10337_),
    .C(_10335_),
    .Y(_10346_));
 sky130_fd_sc_hd__nand3_2 _31981_ (.A(_10345_),
    .B(_10346_),
    .C(_10343_),
    .Y(_10347_));
 sky130_fd_sc_hd__nand2_2 _31982_ (.A(_10344_),
    .B(_10347_),
    .Y(_10348_));
 sky130_fd_sc_hd__nand3_2 _31983_ (.A(_09729_),
    .B(_09732_),
    .C(_09734_),
    .Y(_10349_));
 sky130_fd_sc_hd__nand2_2 _31984_ (.A(_10033_),
    .B(_10349_),
    .Y(_10350_));
 sky130_fd_sc_hd__nor2_2 _31985_ (.A(_10350_),
    .B(_10032_),
    .Y(_10351_));
 sky130_fd_sc_hd__a21oi_2 _31986_ (.A1(_10029_),
    .A2(_10030_),
    .B1(_10027_),
    .Y(_10352_));
 sky130_fd_sc_hd__a21oi_2 _31987_ (.A1(_10349_),
    .A2(_10031_),
    .B1(_10352_),
    .Y(_10353_));
 sky130_fd_sc_hd__a21oi_2 _31988_ (.A1(_09752_),
    .A2(_10351_),
    .B1(_10353_),
    .Y(_10354_));
 sky130_fd_sc_hd__xor2_2 _31989_ (.A(_10348_),
    .B(_10354_),
    .X(_02649_));
 sky130_fd_sc_hd__a22oi_2 _31990_ (.A1(_10120_),
    .A2(_06607_),
    .B1(_08391_),
    .B2(_08256_),
    .Y(_10355_));
 sky130_fd_sc_hd__buf_1 _31991_ (.A(_07468_),
    .X(_10356_));
 sky130_fd_sc_hd__and4_2 _31992_ (.A(_10356_),
    .B(_08908_),
    .C(_08256_),
    .D(_07102_),
    .X(_10357_));
 sky130_fd_sc_hd__and2_2 _31993_ (.A(_07477_),
    .B(_08510_),
    .X(_10358_));
 sky130_fd_sc_hd__o21bai_2 _31994_ (.A1(_10355_),
    .A2(_10357_),
    .B1_N(_10358_),
    .Y(_10359_));
 sky130_fd_sc_hd__nand2_2 _31995_ (.A(_18780_),
    .B(_06453_),
    .Y(_10360_));
 sky130_fd_sc_hd__nand3b_2 _31996_ (.A_N(_10360_),
    .B(_08142_),
    .C(_06596_),
    .Y(_10361_));
 sky130_fd_sc_hd__nand3b_2 _31997_ (.A_N(_10355_),
    .B(_10361_),
    .C(_10358_),
    .Y(_10362_));
 sky130_fd_sc_hd__nand2_2 _31998_ (.A(_10359_),
    .B(_10362_),
    .Y(_10363_));
 sky130_fd_sc_hd__a21oi_2 _31999_ (.A1(_10205_),
    .A2(_10204_),
    .B1(_10203_),
    .Y(_10364_));
 sky130_fd_sc_hd__nand2_2 _32000_ (.A(_10363_),
    .B(_10364_),
    .Y(_10365_));
 sky130_fd_sc_hd__nand3b_2 _32001_ (.A_N(_10364_),
    .B(_10359_),
    .C(_10362_),
    .Y(_10366_));
 sky130_fd_sc_hd__nand2_2 _32002_ (.A(_10365_),
    .B(_10366_),
    .Y(_10367_));
 sky130_fd_sc_hd__a21oi_2 _32003_ (.A1(_10128_),
    .A2(_10125_),
    .B1(_10124_),
    .Y(_10368_));
 sky130_fd_sc_hd__nand2_2 _32004_ (.A(_10367_),
    .B(_10368_),
    .Y(_10369_));
 sky130_fd_sc_hd__nand3b_2 _32005_ (.A_N(_10368_),
    .B(_10365_),
    .C(_10366_),
    .Y(_10370_));
 sky130_fd_sc_hd__nand2_2 _32006_ (.A(_10137_),
    .B(_10133_),
    .Y(_10371_));
 sky130_fd_sc_hd__a21o_2 _32007_ (.A1(_10369_),
    .A2(_10370_),
    .B1(_10371_),
    .X(_10372_));
 sky130_fd_sc_hd__nand3_2 _32008_ (.A(_10371_),
    .B(_10369_),
    .C(_10370_),
    .Y(_10373_));
 sky130_fd_sc_hd__buf_1 _32009_ (.A(_10373_),
    .X(_10374_));
 sky130_fd_sc_hd__nand2_2 _32010_ (.A(_08032_),
    .B(_08258_),
    .Y(_10375_));
 sky130_fd_sc_hd__buf_1 _32011_ (.A(_07105_),
    .X(_10376_));
 sky130_fd_sc_hd__nand2_2 _32012_ (.A(_07824_),
    .B(_10376_),
    .Y(_10377_));
 sky130_fd_sc_hd__nand2_2 _32013_ (.A(_10375_),
    .B(_10377_),
    .Y(_10378_));
 sky130_fd_sc_hd__buf_1 _32014_ (.A(_09364_),
    .X(_10379_));
 sky130_fd_sc_hd__nand3b_2 _32015_ (.A_N(_10375_),
    .B(_08043_),
    .C(_10379_),
    .Y(_10380_));
 sky130_fd_sc_hd__o2bb2ai_2 _32016_ (.A1_N(_10378_),
    .A2_N(_10380_),
    .B1(_18810_),
    .B2(_09665_),
    .Y(_10381_));
 sky130_fd_sc_hd__buf_1 _32017_ (.A(_06274_),
    .X(_10382_));
 sky130_fd_sc_hd__buf_1 _32018_ (.A(_07743_),
    .X(_10383_));
 sky130_fd_sc_hd__and2_2 _32019_ (.A(_10382_),
    .B(_10383_),
    .X(_10384_));
 sky130_fd_sc_hd__nand3_2 _32020_ (.A(_10380_),
    .B(_10384_),
    .C(_10378_),
    .Y(_10385_));
 sky130_fd_sc_hd__a21oi_2 _32021_ (.A1(_10148_),
    .A2(_10147_),
    .B1(_10146_),
    .Y(_10386_));
 sky130_vsdinv _32022_ (.A(_10386_),
    .Y(_10387_));
 sky130_fd_sc_hd__a21oi_2 _32023_ (.A1(_10381_),
    .A2(_10385_),
    .B1(_10387_),
    .Y(_10388_));
 sky130_fd_sc_hd__nand3_2 _32024_ (.A(_10381_),
    .B(_10387_),
    .C(_10385_),
    .Y(_10389_));
 sky130_vsdinv _32025_ (.A(_10389_),
    .Y(_10390_));
 sky130_fd_sc_hd__and2_2 _32026_ (.A(_06815_),
    .B(_07951_),
    .X(_10391_));
 sky130_fd_sc_hd__buf_1 _32027_ (.A(_10391_),
    .X(_10392_));
 sky130_fd_sc_hd__buf_1 _32028_ (.A(_08178_),
    .X(_10393_));
 sky130_fd_sc_hd__nand2_2 _32029_ (.A(_10393_),
    .B(_07752_),
    .Y(_10394_));
 sky130_fd_sc_hd__nand2_2 _32030_ (.A(_06812_),
    .B(_07963_),
    .Y(_10395_));
 sky130_fd_sc_hd__xnor2_2 _32031_ (.A(_10394_),
    .B(_10395_),
    .Y(_10396_));
 sky130_fd_sc_hd__xor2_2 _32032_ (.A(_10392_),
    .B(_10396_),
    .X(_10397_));
 sky130_fd_sc_hd__o21ai_2 _32033_ (.A1(_10388_),
    .A2(_10390_),
    .B1(_10397_),
    .Y(_10398_));
 sky130_fd_sc_hd__xnor2_2 _32034_ (.A(_10392_),
    .B(_10396_),
    .Y(_10399_));
 sky130_fd_sc_hd__nand3b_2 _32035_ (.A_N(_10388_),
    .B(_10399_),
    .C(_10389_),
    .Y(_10400_));
 sky130_fd_sc_hd__nand2_2 _32036_ (.A(_10398_),
    .B(_10400_),
    .Y(_10401_));
 sky130_fd_sc_hd__buf_1 _32037_ (.A(_10401_),
    .X(_10402_));
 sky130_fd_sc_hd__a21boi_2 _32038_ (.A1(_10372_),
    .A2(_10374_),
    .B1_N(_10402_),
    .Y(_10403_));
 sky130_fd_sc_hd__a21oi_2 _32039_ (.A1(_10369_),
    .A2(_10370_),
    .B1(_10371_),
    .Y(_10404_));
 sky130_fd_sc_hd__nor3b_2 _32040_ (.A(_10402_),
    .B(_10404_),
    .C_N(_10374_),
    .Y(_10405_));
 sky130_fd_sc_hd__nand2_2 _32041_ (.A(_10226_),
    .B(_10221_),
    .Y(_10406_));
 sky130_fd_sc_hd__o21bai_2 _32042_ (.A1(_10403_),
    .A2(_10405_),
    .B1_N(_10406_),
    .Y(_10407_));
 sky130_fd_sc_hd__a21bo_2 _32043_ (.A1(_10372_),
    .A2(_10373_),
    .B1_N(_10402_),
    .X(_10408_));
 sky130_fd_sc_hd__nand3b_2 _32044_ (.A_N(_10401_),
    .B(_10372_),
    .C(_10374_),
    .Y(_10409_));
 sky130_fd_sc_hd__nand3_2 _32045_ (.A(_10408_),
    .B(_10406_),
    .C(_10409_),
    .Y(_10410_));
 sky130_fd_sc_hd__nand2_2 _32046_ (.A(_10407_),
    .B(_10410_),
    .Y(_10411_));
 sky130_fd_sc_hd__a21boi_2 _32047_ (.A1(_10171_),
    .A2(_10140_),
    .B1_N(_10143_),
    .Y(_10412_));
 sky130_fd_sc_hd__nand2_2 _32048_ (.A(_10411_),
    .B(_10412_),
    .Y(_10413_));
 sky130_fd_sc_hd__nand3b_2 _32049_ (.A_N(_10412_),
    .B(_10407_),
    .C(_10410_),
    .Y(_10414_));
 sky130_fd_sc_hd__buf_1 _32050_ (.A(_09266_),
    .X(_10415_));
 sky130_fd_sc_hd__a22oi_2 _32051_ (.A1(_08730_),
    .A2(_06075_),
    .B1(_10415_),
    .B2(_06343_),
    .Y(_10416_));
 sky130_fd_sc_hd__buf_1 _32052_ (.A(_08729_),
    .X(_10417_));
 sky130_fd_sc_hd__and4_2 _32053_ (.A(_10417_),
    .B(_08731_),
    .C(_06061_),
    .D(_05847_),
    .X(_10418_));
 sky130_fd_sc_hd__and2_2 _32054_ (.A(_07845_),
    .B(_06199_),
    .X(_10419_));
 sky130_fd_sc_hd__o21bai_2 _32055_ (.A1(_10416_),
    .A2(_10418_),
    .B1_N(_10419_),
    .Y(_10420_));
 sky130_fd_sc_hd__buf_1 _32056_ (.A(_08463_),
    .X(_10421_));
 sky130_fd_sc_hd__nand2_2 _32057_ (.A(_10421_),
    .B(_06075_),
    .Y(_10422_));
 sky130_fd_sc_hd__nand3b_2 _32058_ (.A_N(_10422_),
    .B(_18754_),
    .C(_05951_),
    .Y(_10423_));
 sky130_fd_sc_hd__nand3b_2 _32059_ (.A_N(_10416_),
    .B(_10423_),
    .C(_10419_),
    .Y(_10424_));
 sky130_fd_sc_hd__nand2_2 _32060_ (.A(_10420_),
    .B(_10424_),
    .Y(_10425_));
 sky130_fd_sc_hd__a21oi_2 _32061_ (.A1(_10194_),
    .A2(_10191_),
    .B1(_10190_),
    .Y(_10426_));
 sky130_fd_sc_hd__nand2_2 _32062_ (.A(_10425_),
    .B(_10426_),
    .Y(_10427_));
 sky130_fd_sc_hd__nand3b_2 _32063_ (.A_N(_10426_),
    .B(_10420_),
    .C(_10424_),
    .Y(_10428_));
 sky130_fd_sc_hd__buf_1 _32064_ (.A(_07851_),
    .X(_10429_));
 sky130_fd_sc_hd__buf_1 _32065_ (.A(_10207_),
    .X(_10430_));
 sky130_fd_sc_hd__a22oi_2 _32066_ (.A1(_10429_),
    .A2(_06197_),
    .B1(_10430_),
    .B2(_06366_),
    .Y(_10431_));
 sky130_fd_sc_hd__nand2_2 _32067_ (.A(_18765_),
    .B(_06589_),
    .Y(_10432_));
 sky130_fd_sc_hd__buf_1 _32068_ (.A(_07535_),
    .X(_10433_));
 sky130_fd_sc_hd__nand2_2 _32069_ (.A(_10433_),
    .B(_06729_),
    .Y(_10434_));
 sky130_fd_sc_hd__nor2_2 _32070_ (.A(_10432_),
    .B(_10434_),
    .Y(_10435_));
 sky130_fd_sc_hd__buf_1 _32071_ (.A(_08990_),
    .X(_10436_));
 sky130_fd_sc_hd__and2_2 _32072_ (.A(_10436_),
    .B(_08054_),
    .X(_10437_));
 sky130_vsdinv _32073_ (.A(_10437_),
    .Y(_10438_));
 sky130_fd_sc_hd__nor3_2 _32074_ (.A(_10431_),
    .B(_10435_),
    .C(_10438_),
    .Y(_10439_));
 sky130_fd_sc_hd__o21a_2 _32075_ (.A1(_10431_),
    .A2(_10435_),
    .B1(_10438_),
    .X(_10440_));
 sky130_fd_sc_hd__nor2_2 _32076_ (.A(_10439_),
    .B(_10440_),
    .Y(_10441_));
 sky130_fd_sc_hd__a21oi_2 _32077_ (.A1(_10427_),
    .A2(_10428_),
    .B1(_10441_),
    .Y(_10442_));
 sky130_fd_sc_hd__nand3_2 _32078_ (.A(_10427_),
    .B(_10441_),
    .C(_10428_),
    .Y(_10443_));
 sky130_vsdinv _32079_ (.A(_10443_),
    .Y(_10444_));
 sky130_fd_sc_hd__nand2_2 _32080_ (.A(_10249_),
    .B(_10244_),
    .Y(_10445_));
 sky130_fd_sc_hd__o21bai_2 _32081_ (.A1(_10442_),
    .A2(_10444_),
    .B1_N(_10445_),
    .Y(_10446_));
 sky130_fd_sc_hd__nand3b_2 _32082_ (.A_N(_10442_),
    .B(_10445_),
    .C(_10443_),
    .Y(_10447_));
 sky130_fd_sc_hd__nand2_2 _32083_ (.A(_10446_),
    .B(_10447_),
    .Y(_10448_));
 sky130_fd_sc_hd__a21oi_2 _32084_ (.A1(_10211_),
    .A2(_10199_),
    .B1(_10214_),
    .Y(_10449_));
 sky130_fd_sc_hd__nand2_2 _32085_ (.A(_10448_),
    .B(_10449_),
    .Y(_10450_));
 sky130_fd_sc_hd__nand3b_2 _32086_ (.A_N(_10449_),
    .B(_10446_),
    .C(_10447_),
    .Y(_10451_));
 sky130_fd_sc_hd__buf_1 _32087_ (.A(_09587_),
    .X(_10452_));
 sky130_fd_sc_hd__buf_1 _32088_ (.A(_08754_),
    .X(_10453_));
 sky130_fd_sc_hd__a22oi_2 _32089_ (.A1(_10452_),
    .A2(_05518_),
    .B1(_10453_),
    .B2(_05931_),
    .Y(_10454_));
 sky130_fd_sc_hd__nand2_2 _32090_ (.A(_09006_),
    .B(_08003_),
    .Y(_10455_));
 sky130_fd_sc_hd__buf_1 _32091_ (.A(_09305_),
    .X(_10456_));
 sky130_fd_sc_hd__nand2_2 _32092_ (.A(_10456_),
    .B(_06052_),
    .Y(_10457_));
 sky130_fd_sc_hd__nor2_2 _32093_ (.A(_10455_),
    .B(_10457_),
    .Y(_10458_));
 sky130_fd_sc_hd__and2_2 _32094_ (.A(_08758_),
    .B(_06043_),
    .X(_10459_));
 sky130_fd_sc_hd__o21bai_2 _32095_ (.A1(_10454_),
    .A2(_10458_),
    .B1_N(_10459_),
    .Y(_10460_));
 sky130_fd_sc_hd__nand3b_2 _32096_ (.A_N(_10455_),
    .B(_08756_),
    .C(_19273_),
    .Y(_10461_));
 sky130_fd_sc_hd__nand3b_2 _32097_ (.A_N(_10454_),
    .B(_10461_),
    .C(_10459_),
    .Y(_10462_));
 sky130_fd_sc_hd__nand2_2 _32098_ (.A(_10460_),
    .B(_10462_),
    .Y(_10463_));
 sky130_fd_sc_hd__a21oi_2 _32099_ (.A1(_10257_),
    .A2(_10256_),
    .B1(_10255_),
    .Y(_10464_));
 sky130_fd_sc_hd__nand2_2 _32100_ (.A(_10463_),
    .B(_10464_),
    .Y(_10465_));
 sky130_fd_sc_hd__nand3b_2 _32101_ (.A_N(_10464_),
    .B(_10462_),
    .C(_10460_),
    .Y(_10466_));
 sky130_fd_sc_hd__nand2_2 _32102_ (.A(_10465_),
    .B(_10466_),
    .Y(_10467_));
 sky130_fd_sc_hd__a21oi_2 _32103_ (.A1(_10237_),
    .A2(_10234_),
    .B1(_10233_),
    .Y(_10468_));
 sky130_fd_sc_hd__nand2_2 _32104_ (.A(_10467_),
    .B(_10468_),
    .Y(_10469_));
 sky130_fd_sc_hd__nand3b_2 _32105_ (.A_N(_10468_),
    .B(_10465_),
    .C(_10466_),
    .Y(_10470_));
 sky130_fd_sc_hd__nand2_2 _32106_ (.A(_09958_),
    .B(_07013_),
    .Y(_10471_));
 sky130_fd_sc_hd__nand2_2 _32107_ (.A(_10262_),
    .B(_05540_),
    .Y(_10472_));
 sky130_fd_sc_hd__nor2_2 _32108_ (.A(_10471_),
    .B(_10472_),
    .Y(_10473_));
 sky130_fd_sc_hd__buf_1 _32109_ (.A(_18722_),
    .X(_10474_));
 sky130_fd_sc_hd__and2_2 _32110_ (.A(_10474_),
    .B(_05555_),
    .X(_10475_));
 sky130_fd_sc_hd__nand2_2 _32111_ (.A(_10471_),
    .B(_10472_),
    .Y(_10476_));
 sky130_fd_sc_hd__nand3b_2 _32112_ (.A_N(_10473_),
    .B(_10475_),
    .C(_10476_),
    .Y(_10477_));
 sky130_fd_sc_hd__a22oi_2 _32113_ (.A1(_10261_),
    .A2(_05494_),
    .B1(_10263_),
    .B2(_05880_),
    .Y(_10478_));
 sky130_fd_sc_hd__o21bai_2 _32114_ (.A1(_10478_),
    .A2(_10473_),
    .B1_N(_10475_),
    .Y(_10479_));
 sky130_fd_sc_hd__buf_1 _32115_ (.A(\pcpi_mul.rs2[31] ),
    .X(_10480_));
 sky130_fd_sc_hd__buf_1 _32116_ (.A(_10480_),
    .X(_10481_));
 sky130_fd_sc_hd__buf_1 _32117_ (.A(_10481_),
    .X(_10482_));
 sky130_fd_sc_hd__buf_1 _32118_ (.A(_10266_),
    .X(_10483_));
 sky130_fd_sc_hd__buf_1 _32119_ (.A(_10483_),
    .X(_10484_));
 sky130_fd_sc_hd__a22oi_2 _32120_ (.A1(_10482_),
    .A2(_06546_),
    .B1(_10484_),
    .B2(_06144_),
    .Y(_10485_));
 sky130_fd_sc_hd__buf_1 _32121_ (.A(_18693_),
    .X(_10486_));
 sky130_fd_sc_hd__buf_1 _32122_ (.A(_10486_),
    .X(_10487_));
 sky130_fd_sc_hd__nand2_2 _32123_ (.A(_10487_),
    .B(_05465_),
    .Y(_10488_));
 sky130_fd_sc_hd__nand2_2 _32124_ (.A(_18704_),
    .B(_05424_),
    .Y(_10489_));
 sky130_fd_sc_hd__nor2_2 _32125_ (.A(_10488_),
    .B(_10489_),
    .Y(_10490_));
 sky130_fd_sc_hd__o2bb2ai_2 _32126_ (.A1_N(_10477_),
    .A2_N(_10479_),
    .B1(_10485_),
    .B2(_10490_),
    .Y(_10491_));
 sky130_fd_sc_hd__nor2_2 _32127_ (.A(_10485_),
    .B(_10490_),
    .Y(_10492_));
 sky130_fd_sc_hd__nand3_2 _32128_ (.A(_10477_),
    .B(_10479_),
    .C(_10492_),
    .Y(_10493_));
 sky130_fd_sc_hd__nand3_2 _32129_ (.A(_10272_),
    .B(_10491_),
    .C(_10493_),
    .Y(_10494_));
 sky130_fd_sc_hd__a21oi_2 _32130_ (.A1(_10477_),
    .A2(_10479_),
    .B1(_10492_),
    .Y(_10495_));
 sky130_vsdinv _32131_ (.A(_10493_),
    .Y(_10496_));
 sky130_fd_sc_hd__o21ai_2 _32132_ (.A1(_10495_),
    .A2(_10496_),
    .B1(_10271_),
    .Y(_10497_));
 sky130_fd_sc_hd__a22oi_2 _32133_ (.A1(_10469_),
    .A2(_10470_),
    .B1(_10494_),
    .B2(_10497_),
    .Y(_10498_));
 sky130_fd_sc_hd__nand2_2 _32134_ (.A(_10469_),
    .B(_10470_),
    .Y(_10499_));
 sky130_fd_sc_hd__nand2_2 _32135_ (.A(_10497_),
    .B(_10494_),
    .Y(_10500_));
 sky130_fd_sc_hd__nor2_2 _32136_ (.A(_10499_),
    .B(_10500_),
    .Y(_10501_));
 sky130_vsdinv _32137_ (.A(_10276_),
    .Y(_10502_));
 sky130_fd_sc_hd__o21bai_2 _32138_ (.A1(_10498_),
    .A2(_10501_),
    .B1_N(_10502_),
    .Y(_10503_));
 sky130_fd_sc_hd__nand3b_2 _32139_ (.A_N(_10499_),
    .B(_10494_),
    .C(_10497_),
    .Y(_10504_));
 sky130_fd_sc_hd__nand2_2 _32140_ (.A(_10500_),
    .B(_10499_),
    .Y(_10505_));
 sky130_fd_sc_hd__nand3_2 _32141_ (.A(_10504_),
    .B(_10502_),
    .C(_10505_),
    .Y(_10506_));
 sky130_fd_sc_hd__buf_1 _32142_ (.A(_10506_),
    .X(_10507_));
 sky130_fd_sc_hd__a22oi_2 _32143_ (.A1(_10450_),
    .A2(_10451_),
    .B1(_10503_),
    .B2(_10507_),
    .Y(_10508_));
 sky130_fd_sc_hd__nand2_2 _32144_ (.A(_10450_),
    .B(_10451_),
    .Y(_10509_));
 sky130_fd_sc_hd__nand2_2 _32145_ (.A(_10503_),
    .B(_10506_),
    .Y(_10510_));
 sky130_fd_sc_hd__nor2_2 _32146_ (.A(_10509_),
    .B(_10510_),
    .Y(_10511_));
 sky130_vsdinv _32147_ (.A(_10277_),
    .Y(_10512_));
 sky130_fd_sc_hd__a31oi_2 _32148_ (.A1(_10279_),
    .A2(_10224_),
    .A3(_10227_),
    .B1(_10512_),
    .Y(_10513_));
 sky130_fd_sc_hd__o21ai_2 _32149_ (.A1(_10508_),
    .A2(_10511_),
    .B1(_10513_),
    .Y(_10514_));
 sky130_fd_sc_hd__and2_2 _32150_ (.A(_10450_),
    .B(_10451_),
    .X(_10515_));
 sky130_fd_sc_hd__nand3_2 _32151_ (.A(_10515_),
    .B(_10507_),
    .C(_10503_),
    .Y(_10516_));
 sky130_fd_sc_hd__o21bai_2 _32152_ (.A1(_10281_),
    .A2(_10282_),
    .B1_N(_10512_),
    .Y(_10517_));
 sky130_fd_sc_hd__nand2_2 _32153_ (.A(_10510_),
    .B(_10509_),
    .Y(_10518_));
 sky130_fd_sc_hd__nand3_2 _32154_ (.A(_10516_),
    .B(_10517_),
    .C(_10518_),
    .Y(_10519_));
 sky130_fd_sc_hd__a22oi_2 _32155_ (.A1(_10413_),
    .A2(_10414_),
    .B1(_10514_),
    .B2(_10519_),
    .Y(_10520_));
 sky130_fd_sc_hd__nand2_2 _32156_ (.A(_10413_),
    .B(_10414_),
    .Y(_10521_));
 sky130_fd_sc_hd__nand2_2 _32157_ (.A(_10514_),
    .B(_10519_),
    .Y(_10522_));
 sky130_fd_sc_hd__nor2_2 _32158_ (.A(_10521_),
    .B(_10522_),
    .Y(_10523_));
 sky130_fd_sc_hd__a21boi_2 _32159_ (.A1(_10304_),
    .A2(_10285_),
    .B1_N(_10293_),
    .Y(_10524_));
 sky130_fd_sc_hd__o21ai_2 _32160_ (.A1(_10520_),
    .A2(_10523_),
    .B1(_10524_),
    .Y(_10525_));
 sky130_fd_sc_hd__nand3b_2 _32161_ (.A_N(_10521_),
    .B(_10519_),
    .C(_10514_),
    .Y(_10526_));
 sky130_fd_sc_hd__o21ai_2 _32162_ (.A1(_10295_),
    .A2(_10296_),
    .B1(_10293_),
    .Y(_10527_));
 sky130_fd_sc_hd__nand2_2 _32163_ (.A(_10522_),
    .B(_10521_),
    .Y(_10528_));
 sky130_fd_sc_hd__nand3_2 _32164_ (.A(_10526_),
    .B(_10527_),
    .C(_10528_),
    .Y(_10529_));
 sky130_fd_sc_hd__nand2_2 _32165_ (.A(_10525_),
    .B(_10529_),
    .Y(_10530_));
 sky130_fd_sc_hd__buf_1 _32166_ (.A(_19161_),
    .X(_10531_));
 sky130_fd_sc_hd__buf_1 _32167_ (.A(\pcpi_mul.rs1[27] ),
    .X(_10532_));
 sky130_fd_sc_hd__buf_1 _32168_ (.A(_10532_),
    .X(_10533_));
 sky130_fd_sc_hd__a22o_2 _32169_ (.A1(_06586_),
    .A2(_10531_),
    .B1(_05463_),
    .B2(_10533_),
    .X(_10534_));
 sky130_fd_sc_hd__buf_1 _32170_ (.A(\pcpi_mul.rs1[27] ),
    .X(_10535_));
 sky130_fd_sc_hd__nand2_2 _32171_ (.A(_08291_),
    .B(_10535_),
    .Y(_10536_));
 sky130_fd_sc_hd__buf_1 _32172_ (.A(\pcpi_mul.rs1[26] ),
    .X(_10537_));
 sky130_fd_sc_hd__buf_1 _32173_ (.A(_10537_),
    .X(_10538_));
 sky130_fd_sc_hd__nand3b_2 _32174_ (.A_N(_10536_),
    .B(_05825_),
    .C(_10538_),
    .Y(_10539_));
 sky130_fd_sc_hd__buf_1 _32175_ (.A(\pcpi_mul.rs1[31] ),
    .X(_10540_));
 sky130_vsdinv _32176_ (.A(_10540_),
    .Y(_10541_));
 sky130_fd_sc_hd__o2bb2ai_2 _32177_ (.A1_N(_10534_),
    .A2_N(_10539_),
    .B1(_06346_),
    .B2(_10541_),
    .Y(_10542_));
 sky130_fd_sc_hd__and2_2 _32178_ (.A(_06349_),
    .B(_10540_),
    .X(_10543_));
 sky130_fd_sc_hd__nand3_2 _32179_ (.A(_10539_),
    .B(_10534_),
    .C(_10543_),
    .Y(_10544_));
 sky130_fd_sc_hd__a21oi_2 _32180_ (.A1(_10038_),
    .A2(_10040_),
    .B1(_10037_),
    .Y(_10545_));
 sky130_vsdinv _32181_ (.A(_10545_),
    .Y(_10546_));
 sky130_fd_sc_hd__a21o_2 _32182_ (.A1(_10542_),
    .A2(_10544_),
    .B1(_10546_),
    .X(_10547_));
 sky130_fd_sc_hd__buf_1 _32183_ (.A(_10547_),
    .X(_10548_));
 sky130_fd_sc_hd__nand3_2 _32184_ (.A(_10542_),
    .B(_10546_),
    .C(_10544_),
    .Y(_10549_));
 sky130_fd_sc_hd__buf_1 _32185_ (.A(_10549_),
    .X(_10550_));
 sky130_fd_sc_hd__buf_1 _32186_ (.A(_09804_),
    .X(_10551_));
 sky130_fd_sc_hd__and2_2 _32187_ (.A(_06073_),
    .B(_10551_),
    .X(_10552_));
 sky130_vsdinv _32188_ (.A(_10552_),
    .Y(_10553_));
 sky130_fd_sc_hd__buf_1 _32189_ (.A(\pcpi_mul.rs1[29] ),
    .X(_10554_));
 sky130_fd_sc_hd__buf_1 _32190_ (.A(_10554_),
    .X(_10555_));
 sky130_fd_sc_hd__nand2_2 _32191_ (.A(_05421_),
    .B(_10555_),
    .Y(_10556_));
 sky130_fd_sc_hd__nand2_2 _32192_ (.A(_05526_),
    .B(_10039_),
    .Y(_10557_));
 sky130_fd_sc_hd__xnor2_2 _32193_ (.A(_10556_),
    .B(_10557_),
    .Y(_10558_));
 sky130_fd_sc_hd__xor2_2 _32194_ (.A(_10553_),
    .B(_10558_),
    .X(_10559_));
 sky130_fd_sc_hd__buf_1 _32195_ (.A(_10559_),
    .X(_10560_));
 sky130_fd_sc_hd__a21oi_2 _32196_ (.A1(_10548_),
    .A2(_10550_),
    .B1(_10560_),
    .Y(_10561_));
 sky130_fd_sc_hd__and3_2 _32197_ (.A(_10559_),
    .B(_10547_),
    .C(_10549_),
    .X(_10562_));
 sky130_fd_sc_hd__a21boi_2 _32198_ (.A1(_10041_),
    .A2(_10045_),
    .B1_N(_10046_),
    .Y(_10563_));
 sky130_fd_sc_hd__o21ai_2 _32199_ (.A1(_10563_),
    .A2(_10057_),
    .B1(_10048_),
    .Y(_10564_));
 sky130_fd_sc_hd__o21bai_2 _32200_ (.A1(_10561_),
    .A2(_10562_),
    .B1_N(_10564_),
    .Y(_10565_));
 sky130_fd_sc_hd__o21a_2 _32201_ (.A1(_10049_),
    .A2(_10050_),
    .B1(_10054_),
    .X(_10566_));
 sky130_vsdinv _32202_ (.A(_10566_),
    .Y(_10567_));
 sky130_fd_sc_hd__a21o_2 _32203_ (.A1(_10548_),
    .A2(_10550_),
    .B1(_10560_),
    .X(_10568_));
 sky130_fd_sc_hd__nand3_2 _32204_ (.A(_10560_),
    .B(_10548_),
    .C(_10550_),
    .Y(_10569_));
 sky130_fd_sc_hd__nand3_2 _32205_ (.A(_10568_),
    .B(_10564_),
    .C(_10569_),
    .Y(_10570_));
 sky130_fd_sc_hd__nand3_2 _32206_ (.A(_10565_),
    .B(_10567_),
    .C(_10570_),
    .Y(_10571_));
 sky130_vsdinv _32207_ (.A(_10571_),
    .Y(_10572_));
 sky130_fd_sc_hd__a21oi_2 _32208_ (.A1(_10565_),
    .A2(_10570_),
    .B1(_10567_),
    .Y(_10573_));
 sky130_fd_sc_hd__buf_1 _32209_ (.A(_19179_),
    .X(_10574_));
 sky130_fd_sc_hd__buf_1 _32210_ (.A(_10574_),
    .X(_10575_));
 sky130_fd_sc_hd__buf_1 _32211_ (.A(_19172_),
    .X(_10576_));
 sky130_fd_sc_hd__a22oi_2 _32212_ (.A1(_05983_),
    .A2(_10575_),
    .B1(_05769_),
    .B2(_10576_),
    .Y(_10577_));
 sky130_fd_sc_hd__nand2_2 _32213_ (.A(_05982_),
    .B(_09492_),
    .Y(_10578_));
 sky130_fd_sc_hd__nand2_2 _32214_ (.A(_05993_),
    .B(_08833_),
    .Y(_10579_));
 sky130_fd_sc_hd__nor2_2 _32215_ (.A(_10578_),
    .B(_10579_),
    .Y(_10580_));
 sky130_fd_sc_hd__and2_2 _32216_ (.A(_06771_),
    .B(_09786_),
    .X(_10581_));
 sky130_fd_sc_hd__o21bai_2 _32217_ (.A1(_10577_),
    .A2(_10580_),
    .B1_N(_10581_),
    .Y(_10582_));
 sky130_fd_sc_hd__buf_1 _32218_ (.A(_08557_),
    .X(_10583_));
 sky130_fd_sc_hd__nand3b_2 _32219_ (.A_N(_10578_),
    .B(_06231_),
    .C(_10583_),
    .Y(_10584_));
 sky130_fd_sc_hd__nand2_2 _32220_ (.A(_10578_),
    .B(_10579_),
    .Y(_10585_));
 sky130_fd_sc_hd__nand3_2 _32221_ (.A(_10584_),
    .B(_10585_),
    .C(_10581_),
    .Y(_10586_));
 sky130_fd_sc_hd__nand2_2 _32222_ (.A(_10582_),
    .B(_10586_),
    .Y(_10587_));
 sky130_fd_sc_hd__nor2_2 _32223_ (.A(_10158_),
    .B(_10160_),
    .Y(_10588_));
 sky130_fd_sc_hd__a21oi_2 _32224_ (.A1(_10161_),
    .A2(_10165_),
    .B1(_10588_),
    .Y(_10589_));
 sky130_fd_sc_hd__nand2_2 _32225_ (.A(_10587_),
    .B(_10589_),
    .Y(_10590_));
 sky130_fd_sc_hd__nand3b_2 _32226_ (.A_N(_10589_),
    .B(_10582_),
    .C(_10586_),
    .Y(_10591_));
 sky130_fd_sc_hd__a21oi_2 _32227_ (.A1(_10079_),
    .A2(_10075_),
    .B1(_10074_),
    .Y(_10592_));
 sky130_vsdinv _32228_ (.A(_10592_),
    .Y(_10593_));
 sky130_fd_sc_hd__a21oi_2 _32229_ (.A1(_10590_),
    .A2(_10591_),
    .B1(_10593_),
    .Y(_10594_));
 sky130_fd_sc_hd__nand3_2 _32230_ (.A(_10590_),
    .B(_10593_),
    .C(_10591_),
    .Y(_10595_));
 sky130_vsdinv _32231_ (.A(_10595_),
    .Y(_10596_));
 sky130_fd_sc_hd__a21boi_2 _32232_ (.A1(_10149_),
    .A2(_10152_),
    .B1_N(_10154_),
    .Y(_10597_));
 sky130_fd_sc_hd__o21ai_2 _32233_ (.A1(_10167_),
    .A2(_10597_),
    .B1(_10156_),
    .Y(_10598_));
 sky130_fd_sc_hd__o21bai_2 _32234_ (.A1(_10594_),
    .A2(_10596_),
    .B1_N(_10598_),
    .Y(_10599_));
 sky130_fd_sc_hd__nand3b_2 _32235_ (.A_N(_10594_),
    .B(_10598_),
    .C(_10595_),
    .Y(_10600_));
 sky130_fd_sc_hd__nand2_2 _32236_ (.A(_10599_),
    .B(_10600_),
    .Y(_10601_));
 sky130_fd_sc_hd__a21boi_2 _32237_ (.A1(_10083_),
    .A2(_10088_),
    .B1_N(_10084_),
    .Y(_10602_));
 sky130_fd_sc_hd__nand2_2 _32238_ (.A(_10601_),
    .B(_10602_),
    .Y(_10603_));
 sky130_fd_sc_hd__nand3b_2 _32239_ (.A_N(_10602_),
    .B(_10599_),
    .C(_10600_),
    .Y(_10604_));
 sky130_fd_sc_hd__a21oi_2 _32240_ (.A1(_10087_),
    .A2(_10089_),
    .B1(_10093_),
    .Y(_10605_));
 sky130_fd_sc_hd__o21ai_2 _32241_ (.A1(_10096_),
    .A2(_10605_),
    .B1(_10094_),
    .Y(_10606_));
 sky130_fd_sc_hd__a21oi_2 _32242_ (.A1(_10603_),
    .A2(_10604_),
    .B1(_10606_),
    .Y(_10607_));
 sky130_fd_sc_hd__nand3_2 _32243_ (.A(_10603_),
    .B(_10604_),
    .C(_10606_),
    .Y(_10608_));
 sky130_vsdinv _32244_ (.A(_10608_),
    .Y(_10609_));
 sky130_fd_sc_hd__o22ai_2 _32245_ (.A1(_10572_),
    .A2(_10573_),
    .B1(_10607_),
    .B2(_10609_),
    .Y(_10610_));
 sky130_fd_sc_hd__nor2_2 _32246_ (.A(_10573_),
    .B(_10572_),
    .Y(_10611_));
 sky130_fd_sc_hd__a21o_2 _32247_ (.A1(_10603_),
    .A2(_10604_),
    .B1(_10606_),
    .X(_10612_));
 sky130_fd_sc_hd__nand3_2 _32248_ (.A(_10611_),
    .B(_10608_),
    .C(_10612_),
    .Y(_10613_));
 sky130_fd_sc_hd__a21oi_2 _32249_ (.A1(_10178_),
    .A2(_10179_),
    .B1(_10177_),
    .Y(_10614_));
 sky130_fd_sc_hd__o21ai_2 _32250_ (.A1(_10182_),
    .A2(_10614_),
    .B1(_10180_),
    .Y(_10615_));
 sky130_fd_sc_hd__a21oi_2 _32251_ (.A1(_10610_),
    .A2(_10613_),
    .B1(_10615_),
    .Y(_10616_));
 sky130_fd_sc_hd__nand3_2 _32252_ (.A(_10610_),
    .B(_10615_),
    .C(_10613_),
    .Y(_10617_));
 sky130_vsdinv _32253_ (.A(_10617_),
    .Y(_10618_));
 sky130_fd_sc_hd__a21oi_2 _32254_ (.A1(_10106_),
    .A2(_10107_),
    .B1(_10104_),
    .Y(_10619_));
 sky130_fd_sc_hd__buf_1 _32255_ (.A(_10619_),
    .X(_10620_));
 sky130_fd_sc_hd__o21ai_2 _32256_ (.A1(_10616_),
    .A2(_10618_),
    .B1(_10620_),
    .Y(_10621_));
 sky130_fd_sc_hd__nand2_2 _32257_ (.A(_10610_),
    .B(_10613_),
    .Y(_10622_));
 sky130_vsdinv _32258_ (.A(_10615_),
    .Y(_10623_));
 sky130_fd_sc_hd__nand2_2 _32259_ (.A(_10622_),
    .B(_10623_),
    .Y(_10624_));
 sky130_fd_sc_hd__buf_1 _32260_ (.A(_10617_),
    .X(_10625_));
 sky130_fd_sc_hd__nand3b_2 _32261_ (.A_N(_10620_),
    .B(_10624_),
    .C(_10625_),
    .Y(_10626_));
 sky130_fd_sc_hd__nand2_2 _32262_ (.A(_10621_),
    .B(_10626_),
    .Y(_10627_));
 sky130_fd_sc_hd__nand2_2 _32263_ (.A(_10530_),
    .B(_10627_),
    .Y(_10628_));
 sky130_fd_sc_hd__a21boi_2 _32264_ (.A1(_10624_),
    .A2(_10625_),
    .B1_N(_10619_),
    .Y(_10629_));
 sky130_fd_sc_hd__nor3_2 _32265_ (.A(_10620_),
    .B(_10616_),
    .C(_10618_),
    .Y(_10630_));
 sky130_fd_sc_hd__nor2_2 _32266_ (.A(_10629_),
    .B(_10630_),
    .Y(_10631_));
 sky130_fd_sc_hd__nand3_2 _32267_ (.A(_10631_),
    .B(_10529_),
    .C(_10525_),
    .Y(_10632_));
 sky130_fd_sc_hd__nand2_2 _32268_ (.A(_10628_),
    .B(_10632_),
    .Y(_10633_));
 sky130_fd_sc_hd__a21oi_2 _32269_ (.A1(_10305_),
    .A2(_10306_),
    .B1(_10301_),
    .Y(_10634_));
 sky130_fd_sc_hd__o21a_2 _32270_ (.A1(_10634_),
    .A2(_10310_),
    .B1(_10308_),
    .X(_10635_));
 sky130_fd_sc_hd__nand2_2 _32271_ (.A(_10633_),
    .B(_10635_),
    .Y(_10636_));
 sky130_fd_sc_hd__o21ai_2 _32272_ (.A1(_10634_),
    .A2(_10310_),
    .B1(_10308_),
    .Y(_10637_));
 sky130_fd_sc_hd__nand3_2 _32273_ (.A(_10637_),
    .B(_10628_),
    .C(_10632_),
    .Y(_10638_));
 sky130_fd_sc_hd__nand2_2 _32274_ (.A(_10636_),
    .B(_10638_),
    .Y(_10639_));
 sky130_fd_sc_hd__a21boi_2 _32275_ (.A1(_10063_),
    .A2(_10065_),
    .B1_N(_10066_),
    .Y(_10640_));
 sky130_fd_sc_hd__o21ai_2 _32276_ (.A1(_10115_),
    .A2(_10111_),
    .B1(_10118_),
    .Y(_10641_));
 sky130_fd_sc_hd__xnor2_2 _32277_ (.A(_10640_),
    .B(_10641_),
    .Y(_10642_));
 sky130_vsdinv _32278_ (.A(_10642_),
    .Y(_10643_));
 sky130_fd_sc_hd__nand2_2 _32279_ (.A(_10639_),
    .B(_10643_),
    .Y(_10644_));
 sky130_fd_sc_hd__nand3_2 _32280_ (.A(_10636_),
    .B(_10642_),
    .C(_10638_),
    .Y(_10645_));
 sky130_fd_sc_hd__a21oi_2 _32281_ (.A1(_10320_),
    .A2(_10321_),
    .B1(_10316_),
    .Y(_10646_));
 sky130_fd_sc_hd__o21ai_2 _32282_ (.A1(_10333_),
    .A2(_10646_),
    .B1(_10322_),
    .Y(_10647_));
 sky130_fd_sc_hd__a21oi_2 _32283_ (.A1(_10644_),
    .A2(_10645_),
    .B1(_10647_),
    .Y(_10648_));
 sky130_fd_sc_hd__nand3_2 _32284_ (.A(_10644_),
    .B(_10645_),
    .C(_10647_),
    .Y(_10649_));
 sky130_vsdinv _32285_ (.A(_10649_),
    .Y(_10650_));
 sky130_fd_sc_hd__a21oi_2 _32286_ (.A1(_09839_),
    .A2(_09838_),
    .B1(_10323_),
    .Y(_10651_));
 sky130_fd_sc_hd__o21bai_2 _32287_ (.A1(_10648_),
    .A2(_10650_),
    .B1_N(_10651_),
    .Y(_10652_));
 sky130_fd_sc_hd__a21oi_2 _32288_ (.A1(_10636_),
    .A2(_10638_),
    .B1(_10642_),
    .Y(_10653_));
 sky130_fd_sc_hd__a21oi_2 _32289_ (.A1(_10628_),
    .A2(_10632_),
    .B1(_10637_),
    .Y(_10654_));
 sky130_fd_sc_hd__nor2_2 _32290_ (.A(_10635_),
    .B(_10633_),
    .Y(_10655_));
 sky130_fd_sc_hd__nor3_2 _32291_ (.A(_10643_),
    .B(_10654_),
    .C(_10655_),
    .Y(_10656_));
 sky130_fd_sc_hd__o21bai_2 _32292_ (.A1(_10653_),
    .A2(_10656_),
    .B1_N(_10647_),
    .Y(_10657_));
 sky130_fd_sc_hd__nand3_2 _32293_ (.A(_10657_),
    .B(_10651_),
    .C(_10649_),
    .Y(_10658_));
 sky130_fd_sc_hd__o21ai_2 _32294_ (.A1(_10339_),
    .A2(_10340_),
    .B1(_10335_),
    .Y(_10659_));
 sky130_fd_sc_hd__a21oi_2 _32295_ (.A1(_10652_),
    .A2(_10658_),
    .B1(_10659_),
    .Y(_10660_));
 sky130_fd_sc_hd__a21oi_2 _32296_ (.A1(_10331_),
    .A2(_10337_),
    .B1(_10341_),
    .Y(_10661_));
 sky130_fd_sc_hd__a21oi_2 _32297_ (.A1(_10657_),
    .A2(_10649_),
    .B1(_10651_),
    .Y(_10662_));
 sky130_vsdinv _32298_ (.A(_10651_),
    .Y(_10663_));
 sky130_fd_sc_hd__nor3_2 _32299_ (.A(_10663_),
    .B(_10648_),
    .C(_10650_),
    .Y(_10664_));
 sky130_fd_sc_hd__nor3_2 _32300_ (.A(_10661_),
    .B(_10662_),
    .C(_10664_),
    .Y(_10665_));
 sky130_fd_sc_hd__nor2_2 _32301_ (.A(_10660_),
    .B(_10665_),
    .Y(_10666_));
 sky130_vsdinv _32302_ (.A(_10347_),
    .Y(_10667_));
 sky130_fd_sc_hd__o21bai_2 _32303_ (.A1(_10348_),
    .A2(_10354_),
    .B1_N(_10667_),
    .Y(_10668_));
 sky130_fd_sc_hd__xor2_2 _32304_ (.A(_10666_),
    .B(_10668_),
    .X(_02650_));
 sky130_fd_sc_hd__buf_1 _32305_ (.A(_18693_),
    .X(_10669_));
 sky130_fd_sc_hd__nand2_2 _32306_ (.A(_10669_),
    .B(_05510_),
    .Y(_10670_));
 sky130_fd_sc_hd__buf_1 _32307_ (.A(\pcpi_mul.rs2[32] ),
    .X(_10671_));
 sky130_fd_sc_hd__buf_1 _32308_ (.A(_10671_),
    .X(_10672_));
 sky130_fd_sc_hd__buf_1 _32309_ (.A(_10672_),
    .X(_10673_));
 sky130_fd_sc_hd__nand3b_2 _32310_ (.A_N(_10670_),
    .B(_10673_),
    .C(_19302_),
    .Y(_10674_));
 sky130_fd_sc_hd__buf_1 _32311_ (.A(_16968_),
    .X(_10675_));
 sky130_fd_sc_hd__o21ai_2 _32312_ (.A1(_05465_),
    .A2(_10675_),
    .B1(_10670_),
    .Y(_10676_));
 sky130_fd_sc_hd__and2_2 _32313_ (.A(_10267_),
    .B(_05431_),
    .X(_10677_));
 sky130_fd_sc_hd__a21o_2 _32314_ (.A1(_10674_),
    .A2(_10676_),
    .B1(_10677_),
    .X(_10678_));
 sky130_fd_sc_hd__nand3_2 _32315_ (.A(_10674_),
    .B(_10677_),
    .C(_10676_),
    .Y(_10679_));
 sky130_fd_sc_hd__a21oi_2 _32316_ (.A1(_10678_),
    .A2(_10679_),
    .B1(_10490_),
    .Y(_10680_));
 sky130_fd_sc_hd__nand3_2 _32317_ (.A(_10678_),
    .B(_10490_),
    .C(_10679_),
    .Y(_10681_));
 sky130_vsdinv _32318_ (.A(_10681_),
    .Y(_10682_));
 sky130_fd_sc_hd__buf_1 _32319_ (.A(_18710_),
    .X(_10683_));
 sky130_fd_sc_hd__and4_2 _32320_ (.A(_10683_),
    .B(_09603_),
    .C(_05814_),
    .D(_05987_),
    .X(_10684_));
 sky130_fd_sc_hd__and2_2 _32321_ (.A(_09606_),
    .B(_05927_),
    .X(_10685_));
 sky130_fd_sc_hd__buf_1 _32322_ (.A(\pcpi_mul.rs2[28] ),
    .X(_10686_));
 sky130_fd_sc_hd__buf_1 _32323_ (.A(_10686_),
    .X(_10687_));
 sky130_fd_sc_hd__a22oi_2 _32324_ (.A1(_18711_),
    .A2(_05639_),
    .B1(_10687_),
    .B2(_07403_),
    .Y(_10688_));
 sky130_vsdinv _32325_ (.A(_10688_),
    .Y(_10689_));
 sky130_fd_sc_hd__nand3b_2 _32326_ (.A_N(_10684_),
    .B(_10685_),
    .C(_10689_),
    .Y(_10690_));
 sky130_fd_sc_hd__o21bai_2 _32327_ (.A1(_10688_),
    .A2(_10684_),
    .B1_N(_10685_),
    .Y(_10691_));
 sky130_fd_sc_hd__nand2_2 _32328_ (.A(_10690_),
    .B(_10691_),
    .Y(_10692_));
 sky130_vsdinv _32329_ (.A(_10692_),
    .Y(_10693_));
 sky130_fd_sc_hd__o21bai_2 _32330_ (.A1(_10680_),
    .A2(_10682_),
    .B1_N(_10693_),
    .Y(_10694_));
 sky130_fd_sc_hd__o2bb2ai_2 _32331_ (.A1_N(_10679_),
    .A2_N(_10678_),
    .B1(_10488_),
    .B2(_10489_),
    .Y(_10695_));
 sky130_fd_sc_hd__nand3_2 _32332_ (.A(_10695_),
    .B(_10693_),
    .C(_10681_),
    .Y(_10696_));
 sky130_fd_sc_hd__nand2_2 _32333_ (.A(_10694_),
    .B(_10696_),
    .Y(_10697_));
 sky130_fd_sc_hd__nand2_2 _32334_ (.A(_10697_),
    .B(_10493_),
    .Y(_10698_));
 sky130_fd_sc_hd__nand3_2 _32335_ (.A(_10694_),
    .B(_10496_),
    .C(_10696_),
    .Y(_10699_));
 sky130_fd_sc_hd__nand2_2 _32336_ (.A(_09303_),
    .B(_07365_),
    .Y(_10700_));
 sky130_fd_sc_hd__nand2_2 _32337_ (.A(_18734_),
    .B(_05741_),
    .Y(_10701_));
 sky130_fd_sc_hd__xor2_2 _32338_ (.A(_10700_),
    .B(_10701_),
    .X(_10702_));
 sky130_fd_sc_hd__buf_1 _32339_ (.A(_09308_),
    .X(_10703_));
 sky130_fd_sc_hd__and2_2 _32340_ (.A(_10703_),
    .B(_05847_),
    .X(_10704_));
 sky130_fd_sc_hd__nand2_2 _32341_ (.A(_10702_),
    .B(_10704_),
    .Y(_10705_));
 sky130_fd_sc_hd__xnor2_2 _32342_ (.A(_10700_),
    .B(_10701_),
    .Y(_10706_));
 sky130_fd_sc_hd__o21ai_2 _32343_ (.A1(_18741_),
    .A2(_19263_),
    .B1(_10706_),
    .Y(_10707_));
 sky130_fd_sc_hd__nand2_2 _32344_ (.A(_10705_),
    .B(_10707_),
    .Y(_10708_));
 sky130_fd_sc_hd__a21oi_2 _32345_ (.A1(_10476_),
    .A2(_10475_),
    .B1(_10473_),
    .Y(_10709_));
 sky130_fd_sc_hd__nand2_2 _32346_ (.A(_10708_),
    .B(_10709_),
    .Y(_10710_));
 sky130_fd_sc_hd__nand3b_2 _32347_ (.A_N(_10709_),
    .B(_10705_),
    .C(_10707_),
    .Y(_10711_));
 sky130_fd_sc_hd__o31a_2 _32348_ (.A1(_18741_),
    .A2(_19268_),
    .A3(_10454_),
    .B1(_10461_),
    .X(_10712_));
 sky130_vsdinv _32349_ (.A(_10712_),
    .Y(_10713_));
 sky130_fd_sc_hd__a21oi_2 _32350_ (.A1(_10710_),
    .A2(_10711_),
    .B1(_10713_),
    .Y(_10714_));
 sky130_fd_sc_hd__nand3_2 _32351_ (.A(_10710_),
    .B(_10713_),
    .C(_10711_),
    .Y(_10715_));
 sky130_vsdinv _32352_ (.A(_10715_),
    .Y(_10716_));
 sky130_fd_sc_hd__nor2_2 _32353_ (.A(_10714_),
    .B(_10716_),
    .Y(_10717_));
 sky130_fd_sc_hd__a21oi_2 _32354_ (.A1(_10698_),
    .A2(_10699_),
    .B1(_10717_),
    .Y(_10718_));
 sky130_fd_sc_hd__a21o_2 _32355_ (.A1(_10710_),
    .A2(_10711_),
    .B1(_10713_),
    .X(_10719_));
 sky130_fd_sc_hd__nand2_2 _32356_ (.A(_10719_),
    .B(_10715_),
    .Y(_10720_));
 sky130_fd_sc_hd__a21oi_2 _32357_ (.A1(_10694_),
    .A2(_10696_),
    .B1(_10496_),
    .Y(_10721_));
 sky130_vsdinv _32358_ (.A(_10699_),
    .Y(_10722_));
 sky130_fd_sc_hd__nor3_2 _32359_ (.A(_10720_),
    .B(_10721_),
    .C(_10722_),
    .Y(_10723_));
 sky130_vsdinv _32360_ (.A(_10494_),
    .Y(_10724_));
 sky130_fd_sc_hd__a31oi_2 _32361_ (.A1(_10497_),
    .A2(_10469_),
    .A3(_10470_),
    .B1(_10724_),
    .Y(_10725_));
 sky130_vsdinv _32362_ (.A(_10725_),
    .Y(_10726_));
 sky130_fd_sc_hd__o21bai_2 _32363_ (.A1(_10718_),
    .A2(_10723_),
    .B1_N(_10726_),
    .Y(_10727_));
 sky130_fd_sc_hd__o21bai_2 _32364_ (.A1(_10721_),
    .A2(_10722_),
    .B1_N(_10717_),
    .Y(_10728_));
 sky130_fd_sc_hd__nand3_2 _32365_ (.A(_10698_),
    .B(_10717_),
    .C(_10699_),
    .Y(_10729_));
 sky130_fd_sc_hd__nand3_2 _32366_ (.A(_10728_),
    .B(_10729_),
    .C(_10726_),
    .Y(_10730_));
 sky130_fd_sc_hd__nand2_2 _32367_ (.A(_08472_),
    .B(_08035_),
    .Y(_10731_));
 sky130_fd_sc_hd__nand2_2 _32368_ (.A(_09272_),
    .B(_09340_),
    .Y(_10732_));
 sky130_fd_sc_hd__nand2_2 _32369_ (.A(_10731_),
    .B(_10732_),
    .Y(_10733_));
 sky130_fd_sc_hd__buf_1 _32370_ (.A(_10415_),
    .X(_10734_));
 sky130_fd_sc_hd__nand3b_2 _32371_ (.A_N(_10731_),
    .B(_10734_),
    .C(_06358_),
    .Y(_10735_));
 sky130_fd_sc_hd__buf_1 _32372_ (.A(_08231_),
    .X(_10736_));
 sky130_fd_sc_hd__o2bb2ai_2 _32373_ (.A1_N(_10733_),
    .A2_N(_10735_),
    .B1(_10736_),
    .B2(_19250_),
    .Y(_10737_));
 sky130_fd_sc_hd__and2_2 _32374_ (.A(_08084_),
    .B(_09341_),
    .X(_10738_));
 sky130_fd_sc_hd__nand3_2 _32375_ (.A(_10735_),
    .B(_10738_),
    .C(_10733_),
    .Y(_10739_));
 sky130_fd_sc_hd__o31ai_2 _32376_ (.A1(_10736_),
    .A2(_19254_),
    .A3(_10416_),
    .B1(_10423_),
    .Y(_10740_));
 sky130_fd_sc_hd__a21o_2 _32377_ (.A1(_10737_),
    .A2(_10739_),
    .B1(_10740_),
    .X(_10741_));
 sky130_fd_sc_hd__nand3_2 _32378_ (.A(_10740_),
    .B(_10737_),
    .C(_10739_),
    .Y(_10742_));
 sky130_fd_sc_hd__buf_1 _32379_ (.A(_07304_),
    .X(_10743_));
 sky130_fd_sc_hd__and2_2 _32380_ (.A(_07161_),
    .B(_10743_),
    .X(_10744_));
 sky130_fd_sc_hd__buf_1 _32381_ (.A(_18764_),
    .X(_10745_));
 sky130_fd_sc_hd__nand2_2 _32382_ (.A(_10745_),
    .B(_06478_),
    .Y(_10746_));
 sky130_fd_sc_hd__nand2_2 _32383_ (.A(_18771_),
    .B(_06616_),
    .Y(_10747_));
 sky130_fd_sc_hd__xnor2_2 _32384_ (.A(_10746_),
    .B(_10747_),
    .Y(_10748_));
 sky130_fd_sc_hd__xnor2_2 _32385_ (.A(_10744_),
    .B(_10748_),
    .Y(_10749_));
 sky130_fd_sc_hd__a21oi_2 _32386_ (.A1(_10741_),
    .A2(_10742_),
    .B1(_10749_),
    .Y(_10750_));
 sky130_fd_sc_hd__nand3_2 _32387_ (.A(_10749_),
    .B(_10741_),
    .C(_10742_),
    .Y(_10751_));
 sky130_vsdinv _32388_ (.A(_10751_),
    .Y(_10752_));
 sky130_fd_sc_hd__nand2_2 _32389_ (.A(_10470_),
    .B(_10466_),
    .Y(_10753_));
 sky130_fd_sc_hd__o21bai_2 _32390_ (.A1(_10750_),
    .A2(_10752_),
    .B1_N(_10753_),
    .Y(_10754_));
 sky130_fd_sc_hd__nand3b_2 _32391_ (.A_N(_10750_),
    .B(_10753_),
    .C(_10751_),
    .Y(_10755_));
 sky130_fd_sc_hd__buf_1 _32392_ (.A(_10755_),
    .X(_10756_));
 sky130_fd_sc_hd__a21boi_2 _32393_ (.A1(_10427_),
    .A2(_10441_),
    .B1_N(_10428_),
    .Y(_10757_));
 sky130_vsdinv _32394_ (.A(_10757_),
    .Y(_10758_));
 sky130_fd_sc_hd__a21oi_2 _32395_ (.A1(_10754_),
    .A2(_10756_),
    .B1(_10758_),
    .Y(_10759_));
 sky130_fd_sc_hd__nand3_2 _32396_ (.A(_10754_),
    .B(_10758_),
    .C(_10755_),
    .Y(_10760_));
 sky130_vsdinv _32397_ (.A(_10760_),
    .Y(_10761_));
 sky130_fd_sc_hd__nor2_2 _32398_ (.A(_10759_),
    .B(_10761_),
    .Y(_10762_));
 sky130_fd_sc_hd__a21oi_2 _32399_ (.A1(_10727_),
    .A2(_10730_),
    .B1(_10762_),
    .Y(_10763_));
 sky130_fd_sc_hd__a21o_2 _32400_ (.A1(_10754_),
    .A2(_10756_),
    .B1(_10758_),
    .X(_10764_));
 sky130_fd_sc_hd__nand2_2 _32401_ (.A(_10764_),
    .B(_10760_),
    .Y(_10765_));
 sky130_fd_sc_hd__a21oi_2 _32402_ (.A1(_10728_),
    .A2(_10729_),
    .B1(_10726_),
    .Y(_10766_));
 sky130_fd_sc_hd__nor3_2 _32403_ (.A(_10725_),
    .B(_10718_),
    .C(_10723_),
    .Y(_10767_));
 sky130_fd_sc_hd__nor3_2 _32404_ (.A(_10765_),
    .B(_10766_),
    .C(_10767_),
    .Y(_10768_));
 sky130_fd_sc_hd__o21ai_2 _32405_ (.A1(_10509_),
    .A2(_10510_),
    .B1(_10507_),
    .Y(_10769_));
 sky130_fd_sc_hd__o21bai_2 _32406_ (.A1(_10763_),
    .A2(_10768_),
    .B1_N(_10769_),
    .Y(_10770_));
 sky130_fd_sc_hd__o21bai_2 _32407_ (.A1(_10766_),
    .A2(_10767_),
    .B1_N(_10762_),
    .Y(_10771_));
 sky130_fd_sc_hd__nand3_2 _32408_ (.A(_10727_),
    .B(_10762_),
    .C(_10730_),
    .Y(_10772_));
 sky130_fd_sc_hd__nand3_2 _32409_ (.A(_10771_),
    .B(_10772_),
    .C(_10769_),
    .Y(_10773_));
 sky130_fd_sc_hd__buf_1 _32410_ (.A(_07474_),
    .X(_10774_));
 sky130_fd_sc_hd__buf_1 _32411_ (.A(_08255_),
    .X(_10775_));
 sky130_fd_sc_hd__a22o_2 _32412_ (.A1(_18781_),
    .A2(_06746_),
    .B1(_10774_),
    .B2(_10775_),
    .X(_10776_));
 sky130_fd_sc_hd__buf_1 _32413_ (.A(_07006_),
    .X(_10777_));
 sky130_fd_sc_hd__nand2_2 _32414_ (.A(_10777_),
    .B(_07913_),
    .Y(_10778_));
 sky130_fd_sc_hd__nand3b_2 _32415_ (.A_N(_10778_),
    .B(_10774_),
    .C(_10775_),
    .Y(_10779_));
 sky130_fd_sc_hd__buf_1 _32416_ (.A(_07178_),
    .X(_10780_));
 sky130_fd_sc_hd__o2bb2ai_2 _32417_ (.A1_N(_10776_),
    .A2_N(_10779_),
    .B1(_10780_),
    .B2(_19213_),
    .Y(_10781_));
 sky130_fd_sc_hd__and2_2 _32418_ (.A(_06667_),
    .B(_07948_),
    .X(_10782_));
 sky130_fd_sc_hd__nand3_2 _32419_ (.A(_10779_),
    .B(_10776_),
    .C(_10782_),
    .Y(_10783_));
 sky130_fd_sc_hd__nand2_2 _32420_ (.A(_10432_),
    .B(_10434_),
    .Y(_10784_));
 sky130_fd_sc_hd__a21oi_2 _32421_ (.A1(_10784_),
    .A2(_10437_),
    .B1(_10435_),
    .Y(_10785_));
 sky130_vsdinv _32422_ (.A(_10785_),
    .Y(_10786_));
 sky130_fd_sc_hd__a21o_2 _32423_ (.A1(_10781_),
    .A2(_10783_),
    .B1(_10786_),
    .X(_10787_));
 sky130_fd_sc_hd__nand3_2 _32424_ (.A(_10781_),
    .B(_10786_),
    .C(_10783_),
    .Y(_10788_));
 sky130_fd_sc_hd__o31a_2 _32425_ (.A1(_10780_),
    .A2(_19218_),
    .A3(_10355_),
    .B1(_10361_),
    .X(_10789_));
 sky130_vsdinv _32426_ (.A(_10789_),
    .Y(_10790_));
 sky130_fd_sc_hd__a21oi_2 _32427_ (.A1(_10787_),
    .A2(_10788_),
    .B1(_10790_),
    .Y(_10791_));
 sky130_fd_sc_hd__nand3_2 _32428_ (.A(_10787_),
    .B(_10790_),
    .C(_10788_),
    .Y(_10792_));
 sky130_fd_sc_hd__nand2_2 _32429_ (.A(_10370_),
    .B(_10366_),
    .Y(_10793_));
 sky130_fd_sc_hd__nand3b_2 _32430_ (.A_N(_10791_),
    .B(_10792_),
    .C(_10793_),
    .Y(_10794_));
 sky130_vsdinv _32431_ (.A(_10792_),
    .Y(_10795_));
 sky130_fd_sc_hd__o21bai_2 _32432_ (.A1(_10791_),
    .A2(_10795_),
    .B1_N(_10793_),
    .Y(_10796_));
 sky130_fd_sc_hd__nand2_2 _32433_ (.A(_07503_),
    .B(_07944_),
    .Y(_10797_));
 sky130_fd_sc_hd__nand2_2 _32434_ (.A(_07824_),
    .B(_08292_),
    .Y(_10798_));
 sky130_fd_sc_hd__nand2_2 _32435_ (.A(_10797_),
    .B(_10798_),
    .Y(_10799_));
 sky130_fd_sc_hd__nand3b_2 _32436_ (.A_N(_10797_),
    .B(_06394_),
    .C(_08304_),
    .Y(_10800_));
 sky130_fd_sc_hd__o2bb2ai_2 _32437_ (.A1_N(_10799_),
    .A2_N(_10800_),
    .B1(_18811_),
    .B2(_19198_),
    .Y(_10801_));
 sky130_fd_sc_hd__and2_2 _32438_ (.A(_10382_),
    .B(_07752_),
    .X(_10802_));
 sky130_fd_sc_hd__nand3_2 _32439_ (.A(_10800_),
    .B(_10802_),
    .C(_10799_),
    .Y(_10803_));
 sky130_fd_sc_hd__nor2_2 _32440_ (.A(_10375_),
    .B(_10377_),
    .Y(_10804_));
 sky130_fd_sc_hd__a21oi_2 _32441_ (.A1(_10378_),
    .A2(_10384_),
    .B1(_10804_),
    .Y(_10805_));
 sky130_vsdinv _32442_ (.A(_10805_),
    .Y(_10806_));
 sky130_fd_sc_hd__a21oi_2 _32443_ (.A1(_10801_),
    .A2(_10803_),
    .B1(_10806_),
    .Y(_10807_));
 sky130_fd_sc_hd__and2_2 _32444_ (.A(_06137_),
    .B(_10574_),
    .X(_10808_));
 sky130_fd_sc_hd__nand2_2 _32445_ (.A(_06670_),
    .B(_09456_),
    .Y(_10809_));
 sky130_fd_sc_hd__nand2_2 _32446_ (.A(_06141_),
    .B(_08565_),
    .Y(_10810_));
 sky130_fd_sc_hd__xnor2_2 _32447_ (.A(_10809_),
    .B(_10810_),
    .Y(_10811_));
 sky130_fd_sc_hd__xor2_2 _32448_ (.A(_10808_),
    .B(_10811_),
    .X(_10812_));
 sky130_fd_sc_hd__nand3_2 _32449_ (.A(_10801_),
    .B(_10806_),
    .C(_10803_),
    .Y(_10813_));
 sky130_fd_sc_hd__nor3b_2 _32450_ (.A(_10807_),
    .B(_10812_),
    .C_N(_10813_),
    .Y(_10814_));
 sky130_fd_sc_hd__or2b_2 _32451_ (.A(_10807_),
    .B_N(_10813_),
    .X(_10815_));
 sky130_fd_sc_hd__and2_2 _32452_ (.A(_10815_),
    .B(_10812_),
    .X(_10816_));
 sky130_fd_sc_hd__o2bb2ai_2 _32453_ (.A1_N(_10794_),
    .A2_N(_10796_),
    .B1(_10814_),
    .B2(_10816_),
    .Y(_10817_));
 sky130_fd_sc_hd__xor2_2 _32454_ (.A(_10812_),
    .B(_10815_),
    .X(_10818_));
 sky130_fd_sc_hd__nand3_2 _32455_ (.A(_10818_),
    .B(_10794_),
    .C(_10796_),
    .Y(_10819_));
 sky130_fd_sc_hd__nand2_2 _32456_ (.A(_10451_),
    .B(_10447_),
    .Y(_10820_));
 sky130_fd_sc_hd__a21o_2 _32457_ (.A1(_10817_),
    .A2(_10819_),
    .B1(_10820_),
    .X(_10821_));
 sky130_fd_sc_hd__nand3_2 _32458_ (.A(_10817_),
    .B(_10819_),
    .C(_10820_),
    .Y(_10822_));
 sky130_fd_sc_hd__buf_1 _32459_ (.A(_10822_),
    .X(_10823_));
 sky130_fd_sc_hd__o21a_2 _32460_ (.A1(_10402_),
    .A2(_10404_),
    .B1(_10374_),
    .X(_10824_));
 sky130_vsdinv _32461_ (.A(_10824_),
    .Y(_10825_));
 sky130_fd_sc_hd__a21oi_2 _32462_ (.A1(_10821_),
    .A2(_10823_),
    .B1(_10825_),
    .Y(_10826_));
 sky130_fd_sc_hd__a21oi_2 _32463_ (.A1(_10817_),
    .A2(_10819_),
    .B1(_10820_),
    .Y(_10827_));
 sky130_fd_sc_hd__nor3b_2 _32464_ (.A(_10824_),
    .B(_10827_),
    .C_N(_10822_),
    .Y(_10828_));
 sky130_fd_sc_hd__nor2_2 _32465_ (.A(_10826_),
    .B(_10828_),
    .Y(_10829_));
 sky130_fd_sc_hd__a21oi_2 _32466_ (.A1(_10770_),
    .A2(_10773_),
    .B1(_10829_),
    .Y(_10830_));
 sky130_fd_sc_hd__a21o_2 _32467_ (.A1(_10821_),
    .A2(_10823_),
    .B1(_10825_),
    .X(_10831_));
 sky130_fd_sc_hd__nand3_2 _32468_ (.A(_10821_),
    .B(_10825_),
    .C(_10823_),
    .Y(_10832_));
 sky130_fd_sc_hd__nand2_2 _32469_ (.A(_10831_),
    .B(_10832_),
    .Y(_10833_));
 sky130_fd_sc_hd__a21oi_2 _32470_ (.A1(_10771_),
    .A2(_10772_),
    .B1(_10769_),
    .Y(_10834_));
 sky130_vsdinv _32471_ (.A(_10507_),
    .Y(_10835_));
 sky130_fd_sc_hd__o211a_2 _32472_ (.A1(_10835_),
    .A2(_10511_),
    .B1(_10772_),
    .C1(_10771_),
    .X(_10836_));
 sky130_fd_sc_hd__nor3_2 _32473_ (.A(_10833_),
    .B(_10834_),
    .C(_10836_),
    .Y(_10837_));
 sky130_fd_sc_hd__o21ai_2 _32474_ (.A1(_10521_),
    .A2(_10522_),
    .B1(_10519_),
    .Y(_10838_));
 sky130_fd_sc_hd__o21bai_2 _32475_ (.A1(_10830_),
    .A2(_10837_),
    .B1_N(_10838_),
    .Y(_10839_));
 sky130_fd_sc_hd__o21bai_2 _32476_ (.A1(_10834_),
    .A2(_10836_),
    .B1_N(_10829_),
    .Y(_10840_));
 sky130_fd_sc_hd__nand3_2 _32477_ (.A(_10770_),
    .B(_10829_),
    .C(_10773_),
    .Y(_10841_));
 sky130_fd_sc_hd__nand3_2 _32478_ (.A(_10840_),
    .B(_10841_),
    .C(_10838_),
    .Y(_10842_));
 sky130_fd_sc_hd__buf_1 _32479_ (.A(_08832_),
    .X(_10843_));
 sky130_fd_sc_hd__buf_1 _32480_ (.A(_09511_),
    .X(_10844_));
 sky130_fd_sc_hd__a22o_2 _32481_ (.A1(_06311_),
    .A2(_10843_),
    .B1(_18834_),
    .B2(_10844_),
    .X(_10845_));
 sky130_fd_sc_hd__nand2_2 _32482_ (.A(_05768_),
    .B(_09790_),
    .Y(_10846_));
 sky130_fd_sc_hd__nand3b_2 _32483_ (.A_N(_10846_),
    .B(_05773_),
    .C(_09785_),
    .Y(_10847_));
 sky130_fd_sc_hd__o2bb2ai_2 _32484_ (.A1_N(_10845_),
    .A2_N(_10847_),
    .B1(_06114_),
    .B2(_19163_),
    .Y(_10848_));
 sky130_fd_sc_hd__buf_1 _32485_ (.A(_09808_),
    .X(_10849_));
 sky130_fd_sc_hd__and2_2 _32486_ (.A(_05779_),
    .B(_10849_),
    .X(_10850_));
 sky130_fd_sc_hd__nand3_2 _32487_ (.A(_10847_),
    .B(_10845_),
    .C(_10850_),
    .Y(_10851_));
 sky130_fd_sc_hd__nand2_2 _32488_ (.A(_10394_),
    .B(_10395_),
    .Y(_10852_));
 sky130_fd_sc_hd__nor2_2 _32489_ (.A(_10394_),
    .B(_10395_),
    .Y(_10853_));
 sky130_fd_sc_hd__a21oi_2 _32490_ (.A1(_10852_),
    .A2(_10392_),
    .B1(_10853_),
    .Y(_10854_));
 sky130_vsdinv _32491_ (.A(_10854_),
    .Y(_10855_));
 sky130_fd_sc_hd__a21o_2 _32492_ (.A1(_10848_),
    .A2(_10851_),
    .B1(_10855_),
    .X(_10856_));
 sky130_fd_sc_hd__nand3_2 _32493_ (.A(_10848_),
    .B(_10855_),
    .C(_10851_),
    .Y(_10857_));
 sky130_fd_sc_hd__a21oi_2 _32494_ (.A1(_10585_),
    .A2(_10581_),
    .B1(_10580_),
    .Y(_10858_));
 sky130_vsdinv _32495_ (.A(_10858_),
    .Y(_10859_));
 sky130_fd_sc_hd__a21oi_2 _32496_ (.A1(_10856_),
    .A2(_10857_),
    .B1(_10859_),
    .Y(_10860_));
 sky130_fd_sc_hd__nand3_2 _32497_ (.A(_10856_),
    .B(_10859_),
    .C(_10857_),
    .Y(_10861_));
 sky130_vsdinv _32498_ (.A(_10861_),
    .Y(_10862_));
 sky130_fd_sc_hd__o21ai_2 _32499_ (.A1(_10388_),
    .A2(_10397_),
    .B1(_10389_),
    .Y(_10863_));
 sky130_fd_sc_hd__o21bai_2 _32500_ (.A1(_10860_),
    .A2(_10862_),
    .B1_N(_10863_),
    .Y(_10864_));
 sky130_fd_sc_hd__a21o_2 _32501_ (.A1(_10856_),
    .A2(_10857_),
    .B1(_10859_),
    .X(_10865_));
 sky130_fd_sc_hd__nand3_2 _32502_ (.A(_10865_),
    .B(_10863_),
    .C(_10861_),
    .Y(_10866_));
 sky130_fd_sc_hd__a21boi_2 _32503_ (.A1(_10590_),
    .A2(_10593_),
    .B1_N(_10591_),
    .Y(_10867_));
 sky130_vsdinv _32504_ (.A(_10867_),
    .Y(_10868_));
 sky130_fd_sc_hd__a21oi_2 _32505_ (.A1(_10864_),
    .A2(_10866_),
    .B1(_10868_),
    .Y(_10869_));
 sky130_fd_sc_hd__nand3_2 _32506_ (.A(_10864_),
    .B(_10868_),
    .C(_10866_),
    .Y(_10870_));
 sky130_vsdinv _32507_ (.A(_10870_),
    .Y(_10871_));
 sky130_fd_sc_hd__nand2_2 _32508_ (.A(_10604_),
    .B(_10600_),
    .Y(_10872_));
 sky130_fd_sc_hd__o21bai_2 _32509_ (.A1(_10869_),
    .A2(_10871_),
    .B1_N(_10872_),
    .Y(_10873_));
 sky130_fd_sc_hd__nand3b_2 _32510_ (.A_N(_10869_),
    .B(_10870_),
    .C(_10872_),
    .Y(_10874_));
 sky130_fd_sc_hd__buf_1 _32511_ (.A(_09212_),
    .X(_10875_));
 sky130_fd_sc_hd__nand2_2 _32512_ (.A(_05492_),
    .B(_10875_),
    .Y(_10876_));
 sky130_fd_sc_hd__buf_1 _32513_ (.A(_19149_),
    .X(_10877_));
 sky130_fd_sc_hd__nand2_2 _32514_ (.A(_05732_),
    .B(_10877_),
    .Y(_10878_));
 sky130_fd_sc_hd__xor2_2 _32515_ (.A(_10876_),
    .B(_10878_),
    .X(_10879_));
 sky130_fd_sc_hd__buf_1 _32516_ (.A(\pcpi_mul.rs1[32] ),
    .X(_10880_));
 sky130_fd_sc_hd__buf_1 _32517_ (.A(_10880_),
    .X(_10881_));
 sky130_fd_sc_hd__and2_2 _32518_ (.A(_10881_),
    .B(_18877_),
    .X(_10882_));
 sky130_fd_sc_hd__buf_1 _32519_ (.A(_10882_),
    .X(_10883_));
 sky130_fd_sc_hd__buf_1 _32520_ (.A(_10883_),
    .X(_10884_));
 sky130_fd_sc_hd__nand2_2 _32521_ (.A(_10879_),
    .B(_10884_),
    .Y(_10885_));
 sky130_fd_sc_hd__xnor2_2 _32522_ (.A(_10876_),
    .B(_10878_),
    .Y(_10886_));
 sky130_vsdinv _32523_ (.A(_10882_),
    .Y(_10887_));
 sky130_fd_sc_hd__buf_1 _32524_ (.A(_10887_),
    .X(_10888_));
 sky130_fd_sc_hd__nand2_2 _32525_ (.A(_10886_),
    .B(_10888_),
    .Y(_10889_));
 sky130_fd_sc_hd__nand2_2 _32526_ (.A(_10885_),
    .B(_10889_),
    .Y(_10890_));
 sky130_fd_sc_hd__a21boi_2 _32527_ (.A1(_10534_),
    .A2(_10543_),
    .B1_N(_10539_),
    .Y(_10891_));
 sky130_fd_sc_hd__nand2_2 _32528_ (.A(_10890_),
    .B(_10891_),
    .Y(_10892_));
 sky130_fd_sc_hd__nand3b_2 _32529_ (.A_N(_10891_),
    .B(_10889_),
    .C(_10885_),
    .Y(_10893_));
 sky130_fd_sc_hd__buf_1 _32530_ (.A(_19143_),
    .X(_10894_));
 sky130_fd_sc_hd__buf_1 _32531_ (.A(_10894_),
    .X(_10895_));
 sky130_fd_sc_hd__and2_2 _32532_ (.A(_05439_),
    .B(_10895_),
    .X(_10896_));
 sky130_fd_sc_hd__buf_1 _32533_ (.A(_10039_),
    .X(_10897_));
 sky130_fd_sc_hd__nand2_2 _32534_ (.A(_18867_),
    .B(_10897_),
    .Y(_10898_));
 sky130_fd_sc_hd__buf_1 _32535_ (.A(\pcpi_mul.rs1[31] ),
    .X(_10899_));
 sky130_fd_sc_hd__buf_1 _32536_ (.A(_10899_),
    .X(_10900_));
 sky130_fd_sc_hd__nand2_2 _32537_ (.A(_06363_),
    .B(_10900_),
    .Y(_10901_));
 sky130_fd_sc_hd__xnor2_2 _32538_ (.A(_10898_),
    .B(_10901_),
    .Y(_10902_));
 sky130_fd_sc_hd__xnor2_2 _32539_ (.A(_10896_),
    .B(_10902_),
    .Y(_10903_));
 sky130_fd_sc_hd__a21oi_2 _32540_ (.A1(_10892_),
    .A2(_10893_),
    .B1(_10903_),
    .Y(_10904_));
 sky130_vsdinv _32541_ (.A(_10550_),
    .Y(_10905_));
 sky130_fd_sc_hd__a21oi_2 _32542_ (.A1(_10560_),
    .A2(_10548_),
    .B1(_10905_),
    .Y(_10906_));
 sky130_vsdinv _32543_ (.A(_10906_),
    .Y(_10907_));
 sky130_fd_sc_hd__nand3_2 _32544_ (.A(_10892_),
    .B(_10903_),
    .C(_10893_),
    .Y(_10908_));
 sky130_fd_sc_hd__nand3b_2 _32545_ (.A_N(_10904_),
    .B(_10907_),
    .C(_10908_),
    .Y(_10909_));
 sky130_vsdinv _32546_ (.A(_10908_),
    .Y(_10910_));
 sky130_fd_sc_hd__o21ai_2 _32547_ (.A1(_10904_),
    .A2(_10910_),
    .B1(_10906_),
    .Y(_10911_));
 sky130_fd_sc_hd__buf_1 _32548_ (.A(\pcpi_mul.rs1[30] ),
    .X(_10912_));
 sky130_fd_sc_hd__buf_1 _32549_ (.A(_10912_),
    .X(_10913_));
 sky130_fd_sc_hd__buf_1 _32550_ (.A(_10913_),
    .X(_10914_));
 sky130_fd_sc_hd__buf_1 _32551_ (.A(_10914_),
    .X(_10915_));
 sky130_fd_sc_hd__buf_1 _32552_ (.A(_10915_),
    .X(_10916_));
 sky130_fd_sc_hd__nand3b_2 _32553_ (.A_N(_10556_),
    .B(_18875_),
    .C(_10916_),
    .Y(_10917_));
 sky130_fd_sc_hd__o21a_2 _32554_ (.A1(_10553_),
    .A2(_10558_),
    .B1(_10917_),
    .X(_10918_));
 sky130_fd_sc_hd__a21bo_2 _32555_ (.A1(_10909_),
    .A2(_10911_),
    .B1_N(_10918_),
    .X(_10919_));
 sky130_fd_sc_hd__nand3b_2 _32556_ (.A_N(_10918_),
    .B(_10909_),
    .C(_10911_),
    .Y(_10920_));
 sky130_fd_sc_hd__nand2_2 _32557_ (.A(_10919_),
    .B(_10920_),
    .Y(_10921_));
 sky130_fd_sc_hd__buf_1 _32558_ (.A(_10921_),
    .X(_10922_));
 sky130_fd_sc_hd__a21boi_2 _32559_ (.A1(_10873_),
    .A2(_10874_),
    .B1_N(_10922_),
    .Y(_10923_));
 sky130_fd_sc_hd__nand2_2 _32560_ (.A(_10873_),
    .B(_10874_),
    .Y(_10924_));
 sky130_fd_sc_hd__nor2_2 _32561_ (.A(_10922_),
    .B(_10924_),
    .Y(_10925_));
 sky130_fd_sc_hd__nand2_2 _32562_ (.A(_10414_),
    .B(_10410_),
    .Y(_10926_));
 sky130_fd_sc_hd__o21bai_2 _32563_ (.A1(_10923_),
    .A2(_10925_),
    .B1_N(_10926_),
    .Y(_10927_));
 sky130_fd_sc_hd__nand2_2 _32564_ (.A(_10924_),
    .B(_10922_),
    .Y(_10928_));
 sky130_fd_sc_hd__nand3b_2 _32565_ (.A_N(_10921_),
    .B(_10874_),
    .C(_10873_),
    .Y(_10929_));
 sky130_fd_sc_hd__nand3_2 _32566_ (.A(_10926_),
    .B(_10928_),
    .C(_10929_),
    .Y(_10930_));
 sky130_fd_sc_hd__buf_1 _32567_ (.A(_10930_),
    .X(_10931_));
 sky130_fd_sc_hd__a21oi_2 _32568_ (.A1(_10611_),
    .A2(_10612_),
    .B1(_10609_),
    .Y(_10932_));
 sky130_fd_sc_hd__buf_1 _32569_ (.A(_10932_),
    .X(_10933_));
 sky130_fd_sc_hd__a21boi_2 _32570_ (.A1(_10927_),
    .A2(_10931_),
    .B1_N(_10933_),
    .Y(_10934_));
 sky130_fd_sc_hd__a21oi_2 _32571_ (.A1(_10928_),
    .A2(_10929_),
    .B1(_10926_),
    .Y(_10935_));
 sky130_fd_sc_hd__nor3b_2 _32572_ (.A(_10933_),
    .B(_10935_),
    .C_N(_10930_),
    .Y(_10936_));
 sky130_fd_sc_hd__nor2_2 _32573_ (.A(_10934_),
    .B(_10936_),
    .Y(_10937_));
 sky130_fd_sc_hd__a21oi_2 _32574_ (.A1(_10839_),
    .A2(_10842_),
    .B1(_10937_),
    .Y(_10938_));
 sky130_fd_sc_hd__a21bo_2 _32575_ (.A1(_10927_),
    .A2(_10930_),
    .B1_N(_10933_),
    .X(_10939_));
 sky130_fd_sc_hd__nand3b_2 _32576_ (.A_N(_10932_),
    .B(_10927_),
    .C(_10931_),
    .Y(_10940_));
 sky130_fd_sc_hd__nand2_2 _32577_ (.A(_10939_),
    .B(_10940_),
    .Y(_10941_));
 sky130_fd_sc_hd__a21oi_2 _32578_ (.A1(_10840_),
    .A2(_10841_),
    .B1(_10838_),
    .Y(_10942_));
 sky130_vsdinv _32579_ (.A(_10842_),
    .Y(_10943_));
 sky130_fd_sc_hd__nor3_2 _32580_ (.A(_10941_),
    .B(_10942_),
    .C(_10943_),
    .Y(_10944_));
 sky130_fd_sc_hd__a21boi_2 _32581_ (.A1(_10631_),
    .A2(_10525_),
    .B1_N(_10529_),
    .Y(_10945_));
 sky130_vsdinv _32582_ (.A(_10945_),
    .Y(_10946_));
 sky130_fd_sc_hd__o21bai_2 _32583_ (.A1(_10938_),
    .A2(_10944_),
    .B1_N(_10946_),
    .Y(_10947_));
 sky130_fd_sc_hd__buf_1 _32584_ (.A(_10947_),
    .X(_10948_));
 sky130_fd_sc_hd__o21bai_2 _32585_ (.A1(_10942_),
    .A2(_10943_),
    .B1_N(_10937_),
    .Y(_10949_));
 sky130_fd_sc_hd__nand3_2 _32586_ (.A(_10839_),
    .B(_10937_),
    .C(_10842_),
    .Y(_10950_));
 sky130_fd_sc_hd__nand3_2 _32587_ (.A(_10949_),
    .B(_10950_),
    .C(_10946_),
    .Y(_10951_));
 sky130_vsdinv _32588_ (.A(_10570_),
    .Y(_10952_));
 sky130_fd_sc_hd__o2bb2ai_2 _32589_ (.A1_N(_10625_),
    .A2_N(_10626_),
    .B1(_10952_),
    .B2(_10572_),
    .Y(_10953_));
 sky130_fd_sc_hd__o2111ai_2 _32590_ (.A1(_10620_),
    .A2(_10616_),
    .B1(_10570_),
    .C1(_10571_),
    .D1(_10625_),
    .Y(_10954_));
 sky130_fd_sc_hd__nand2_2 _32591_ (.A(_10953_),
    .B(_10954_),
    .Y(_10955_));
 sky130_fd_sc_hd__xor2_2 _32592_ (.A(_16973_),
    .B(_10955_),
    .X(_10956_));
 sky130_fd_sc_hd__buf_1 _32593_ (.A(_10956_),
    .X(_10957_));
 sky130_fd_sc_hd__a21oi_2 _32594_ (.A1(_10948_),
    .A2(_10951_),
    .B1(_10957_),
    .Y(_10958_));
 sky130_fd_sc_hd__nand3_2 _32595_ (.A(_10947_),
    .B(_10956_),
    .C(_10951_),
    .Y(_10959_));
 sky130_vsdinv _32596_ (.A(_10959_),
    .Y(_10960_));
 sky130_fd_sc_hd__o21ai_2 _32597_ (.A1(_10643_),
    .A2(_10654_),
    .B1(_10638_),
    .Y(_10961_));
 sky130_fd_sc_hd__o21bai_2 _32598_ (.A1(_10958_),
    .A2(_10960_),
    .B1_N(_10961_),
    .Y(_10962_));
 sky130_fd_sc_hd__a21o_2 _32599_ (.A1(_10948_),
    .A2(_10951_),
    .B1(_10957_),
    .X(_10963_));
 sky130_fd_sc_hd__nand3_2 _32600_ (.A(_10963_),
    .B(_10959_),
    .C(_10961_),
    .Y(_10964_));
 sky130_fd_sc_hd__a21oi_2 _32601_ (.A1(_10119_),
    .A2(_10118_),
    .B1(_10640_),
    .Y(_10965_));
 sky130_fd_sc_hd__a21o_2 _32602_ (.A1(_10962_),
    .A2(_10964_),
    .B1(_10965_),
    .X(_10966_));
 sky130_fd_sc_hd__nand3_2 _32603_ (.A(_10962_),
    .B(_10964_),
    .C(_10965_),
    .Y(_10967_));
 sky130_fd_sc_hd__o21ai_2 _32604_ (.A1(_10663_),
    .A2(_10648_),
    .B1(_10649_),
    .Y(_10968_));
 sky130_fd_sc_hd__a21o_2 _32605_ (.A1(_10966_),
    .A2(_10967_),
    .B1(_10968_),
    .X(_10969_));
 sky130_fd_sc_hd__nand3_2 _32606_ (.A(_10966_),
    .B(_10967_),
    .C(_10968_),
    .Y(_10970_));
 sky130_fd_sc_hd__nand2_2 _32607_ (.A(_10969_),
    .B(_10970_),
    .Y(_10971_));
 sky130_fd_sc_hd__o21bai_2 _32608_ (.A1(_10662_),
    .A2(_10664_),
    .B1_N(_10659_),
    .Y(_10972_));
 sky130_fd_sc_hd__nand3_2 _32609_ (.A(_10652_),
    .B(_10658_),
    .C(_10659_),
    .Y(_10973_));
 sky130_fd_sc_hd__nand2_2 _32610_ (.A(_10972_),
    .B(_10973_),
    .Y(_10974_));
 sky130_fd_sc_hd__nor2_2 _32611_ (.A(_10348_),
    .B(_10974_),
    .Y(_10975_));
 sky130_fd_sc_hd__nand2_2 _32612_ (.A(_10975_),
    .B(_10351_),
    .Y(_10976_));
 sky130_fd_sc_hd__nor2_2 _32613_ (.A(_09745_),
    .B(_10976_),
    .Y(_10977_));
 sky130_fd_sc_hd__nand3_2 _32614_ (.A(_06877_),
    .B(_10977_),
    .C(_08651_),
    .Y(_10978_));
 sky130_fd_sc_hd__nand2_2 _32615_ (.A(_08656_),
    .B(_10977_),
    .Y(_10979_));
 sky130_fd_sc_hd__a21oi_2 _32616_ (.A1(_09730_),
    .A2(_09728_),
    .B1(_09727_),
    .Y(_10980_));
 sky130_fd_sc_hd__nor3_2 _32617_ (.A(_10980_),
    .B(_10022_),
    .C(_10026_),
    .Y(_10981_));
 sky130_fd_sc_hd__nor2_2 _32618_ (.A(_10352_),
    .B(_10981_),
    .Y(_10982_));
 sky130_fd_sc_hd__nand2_2 _32619_ (.A(_10982_),
    .B(_09741_),
    .Y(_10983_));
 sky130_fd_sc_hd__a21oi_2 _32620_ (.A1(_10345_),
    .A2(_10346_),
    .B1(_10343_),
    .Y(_10984_));
 sky130_fd_sc_hd__nor2_2 _32621_ (.A(_10984_),
    .B(_10667_),
    .Y(_10985_));
 sky130_fd_sc_hd__nand2_2 _32622_ (.A(_10666_),
    .B(_10985_),
    .Y(_10986_));
 sky130_fd_sc_hd__nor2_2 _32623_ (.A(_10983_),
    .B(_10986_),
    .Y(_10987_));
 sky130_fd_sc_hd__nand3_2 _32624_ (.A(_10666_),
    .B(_10985_),
    .C(_10353_),
    .Y(_10988_));
 sky130_fd_sc_hd__nand2_2 _32625_ (.A(_10667_),
    .B(_10972_),
    .Y(_10989_));
 sky130_fd_sc_hd__nand3_2 _32626_ (.A(_10988_),
    .B(_10973_),
    .C(_10989_),
    .Y(_10990_));
 sky130_fd_sc_hd__a21oi_2 _32627_ (.A1(_10987_),
    .A2(_09751_),
    .B1(_10990_),
    .Y(_10991_));
 sky130_fd_sc_hd__nand3_2 _32628_ (.A(_10978_),
    .B(_10979_),
    .C(_10991_),
    .Y(_10992_));
 sky130_fd_sc_hd__buf_1 _32629_ (.A(_10992_),
    .X(_10993_));
 sky130_fd_sc_hd__xnor2_2 _32630_ (.A(_10971_),
    .B(_10993_),
    .Y(_02651_));
 sky130_fd_sc_hd__buf_1 _32631_ (.A(_18693_),
    .X(_10994_));
 sky130_fd_sc_hd__nand2_2 _32632_ (.A(_10994_),
    .B(_05635_),
    .Y(_10995_));
 sky130_fd_sc_hd__buf_1 _32633_ (.A(\pcpi_mul.rs2[32] ),
    .X(_10996_));
 sky130_fd_sc_hd__buf_1 _32634_ (.A(_10996_),
    .X(_10997_));
 sky130_fd_sc_hd__nand3b_2 _32635_ (.A_N(_10995_),
    .B(_10997_),
    .C(_19298_),
    .Y(_10998_));
 sky130_fd_sc_hd__o21ai_2 _32636_ (.A1(_05424_),
    .A2(_10675_),
    .B1(_10995_),
    .Y(_10999_));
 sky130_fd_sc_hd__and2_2 _32637_ (.A(_10267_),
    .B(_05987_),
    .X(_11000_));
 sky130_fd_sc_hd__a21oi_2 _32638_ (.A1(_10998_),
    .A2(_10999_),
    .B1(_11000_),
    .Y(_11001_));
 sky130_fd_sc_hd__nand3_2 _32639_ (.A(_10998_),
    .B(_11000_),
    .C(_10999_),
    .Y(_11002_));
 sky130_vsdinv _32640_ (.A(_11002_),
    .Y(_11003_));
 sky130_fd_sc_hd__buf_1 _32641_ (.A(_16967_),
    .X(_11004_));
 sky130_fd_sc_hd__buf_1 _32642_ (.A(_11004_),
    .X(_11005_));
 sky130_fd_sc_hd__nor3_2 _32643_ (.A(_06546_),
    .B(_11005_),
    .C(_10670_),
    .Y(_11006_));
 sky130_fd_sc_hd__a21o_2 _32644_ (.A1(_10676_),
    .A2(_10677_),
    .B1(_11006_),
    .X(_11007_));
 sky130_fd_sc_hd__o21bai_2 _32645_ (.A1(_11001_),
    .A2(_11003_),
    .B1_N(_11007_),
    .Y(_11008_));
 sky130_fd_sc_hd__a21o_2 _32646_ (.A1(_10998_),
    .A2(_10999_),
    .B1(_11000_),
    .X(_11009_));
 sky130_fd_sc_hd__nand3_2 _32647_ (.A(_11009_),
    .B(_11007_),
    .C(_11002_),
    .Y(_11010_));
 sky130_fd_sc_hd__buf_1 _32648_ (.A(_10259_),
    .X(_11011_));
 sky130_fd_sc_hd__and4_2 _32649_ (.A(_11011_),
    .B(_10686_),
    .C(_05745_),
    .D(_05674_),
    .X(_11012_));
 sky130_fd_sc_hd__and2_2 _32650_ (.A(_18723_),
    .B(_19272_),
    .X(_11013_));
 sky130_fd_sc_hd__buf_1 _32651_ (.A(_10259_),
    .X(_11014_));
 sky130_fd_sc_hd__buf_1 _32652_ (.A(_10252_),
    .X(_11015_));
 sky130_fd_sc_hd__a22oi_2 _32653_ (.A1(_11014_),
    .A2(_08725_),
    .B1(_11015_),
    .B2(_05745_),
    .Y(_11016_));
 sky130_vsdinv _32654_ (.A(_11016_),
    .Y(_11017_));
 sky130_fd_sc_hd__nand3b_2 _32655_ (.A_N(_11012_),
    .B(_11013_),
    .C(_11017_),
    .Y(_11018_));
 sky130_fd_sc_hd__o21bai_2 _32656_ (.A1(_11016_),
    .A2(_11012_),
    .B1_N(_11013_),
    .Y(_11019_));
 sky130_fd_sc_hd__nand2_2 _32657_ (.A(_11018_),
    .B(_11019_),
    .Y(_11020_));
 sky130_vsdinv _32658_ (.A(_11020_),
    .Y(_11021_));
 sky130_fd_sc_hd__a21oi_2 _32659_ (.A1(_11008_),
    .A2(_11010_),
    .B1(_11021_),
    .Y(_11022_));
 sky130_fd_sc_hd__nand3_2 _32660_ (.A(_11008_),
    .B(_11021_),
    .C(_11010_),
    .Y(_11023_));
 sky130_vsdinv _32661_ (.A(_11023_),
    .Y(_11024_));
 sky130_fd_sc_hd__o21ai_2 _32662_ (.A1(_10692_),
    .A2(_10680_),
    .B1(_10681_),
    .Y(_11025_));
 sky130_fd_sc_hd__o21bai_2 _32663_ (.A1(_11022_),
    .A2(_11024_),
    .B1_N(_11025_),
    .Y(_11026_));
 sky130_fd_sc_hd__a21o_2 _32664_ (.A1(_11008_),
    .A2(_11010_),
    .B1(_11021_),
    .X(_11027_));
 sky130_fd_sc_hd__nand3_2 _32665_ (.A(_11027_),
    .B(_11023_),
    .C(_11025_),
    .Y(_11028_));
 sky130_fd_sc_hd__a21o_2 _32666_ (.A1(_10689_),
    .A2(_10685_),
    .B1(_10684_),
    .X(_11029_));
 sky130_vsdinv _32667_ (.A(_11029_),
    .Y(_11030_));
 sky130_fd_sc_hd__nand2_2 _32668_ (.A(_10229_),
    .B(_05649_),
    .Y(_11031_));
 sky130_fd_sc_hd__nand2_2 _32669_ (.A(_18734_),
    .B(_07499_),
    .Y(_11032_));
 sky130_fd_sc_hd__xor2_2 _32670_ (.A(_11031_),
    .B(_11032_),
    .X(_11033_));
 sky130_fd_sc_hd__and2_2 _32671_ (.A(_10703_),
    .B(_06343_),
    .X(_11034_));
 sky130_fd_sc_hd__nand2_2 _32672_ (.A(_11033_),
    .B(_11034_),
    .Y(_11035_));
 sky130_fd_sc_hd__buf_1 _32673_ (.A(_10245_),
    .X(_11036_));
 sky130_fd_sc_hd__xnor2_2 _32674_ (.A(_11031_),
    .B(_11032_),
    .Y(_11037_));
 sky130_fd_sc_hd__o21ai_2 _32675_ (.A1(_11036_),
    .A2(_19259_),
    .B1(_11037_),
    .Y(_11038_));
 sky130_fd_sc_hd__nand2_2 _32676_ (.A(_11035_),
    .B(_11038_),
    .Y(_11039_));
 sky130_fd_sc_hd__nand2_2 _32677_ (.A(_11030_),
    .B(_11039_),
    .Y(_11040_));
 sky130_fd_sc_hd__nand3_2 _32678_ (.A(_11029_),
    .B(_11035_),
    .C(_11038_),
    .Y(_11041_));
 sky130_fd_sc_hd__buf_1 _32679_ (.A(_10456_),
    .X(_11042_));
 sky130_fd_sc_hd__nand3b_2 _32680_ (.A_N(_10700_),
    .B(_11042_),
    .C(_06317_),
    .Y(_11043_));
 sky130_fd_sc_hd__a21boi_2 _32681_ (.A1(_10702_),
    .A2(_10704_),
    .B1_N(_11043_),
    .Y(_11044_));
 sky130_vsdinv _32682_ (.A(_11044_),
    .Y(_11045_));
 sky130_fd_sc_hd__a21oi_2 _32683_ (.A1(_11040_),
    .A2(_11041_),
    .B1(_11045_),
    .Y(_11046_));
 sky130_fd_sc_hd__nand3_2 _32684_ (.A(_11040_),
    .B(_11045_),
    .C(_11041_),
    .Y(_11047_));
 sky130_vsdinv _32685_ (.A(_11047_),
    .Y(_11048_));
 sky130_fd_sc_hd__nor2_2 _32686_ (.A(_11046_),
    .B(_11048_),
    .Y(_11049_));
 sky130_fd_sc_hd__a21oi_2 _32687_ (.A1(_11026_),
    .A2(_11028_),
    .B1(_11049_),
    .Y(_11050_));
 sky130_fd_sc_hd__a21oi_2 _32688_ (.A1(_11035_),
    .A2(_11038_),
    .B1(_11029_),
    .Y(_11051_));
 sky130_vsdinv _32689_ (.A(_11041_),
    .Y(_11052_));
 sky130_fd_sc_hd__o21bai_2 _32690_ (.A1(_11051_),
    .A2(_11052_),
    .B1_N(_11045_),
    .Y(_11053_));
 sky130_fd_sc_hd__nand2_2 _32691_ (.A(_11053_),
    .B(_11047_),
    .Y(_11054_));
 sky130_fd_sc_hd__a21oi_2 _32692_ (.A1(_11027_),
    .A2(_11023_),
    .B1(_11025_),
    .Y(_11055_));
 sky130_vsdinv _32693_ (.A(_11028_),
    .Y(_11056_));
 sky130_fd_sc_hd__nor3_2 _32694_ (.A(_11054_),
    .B(_11055_),
    .C(_11056_),
    .Y(_11057_));
 sky130_fd_sc_hd__o21ai_2 _32695_ (.A1(_10720_),
    .A2(_10721_),
    .B1(_10699_),
    .Y(_11058_));
 sky130_fd_sc_hd__o21bai_2 _32696_ (.A1(_11050_),
    .A2(_11057_),
    .B1_N(_11058_),
    .Y(_11059_));
 sky130_fd_sc_hd__o22ai_2 _32697_ (.A1(_11048_),
    .A2(_11046_),
    .B1(_11055_),
    .B2(_11056_),
    .Y(_11060_));
 sky130_fd_sc_hd__nand3_2 _32698_ (.A(_11049_),
    .B(_11026_),
    .C(_11028_),
    .Y(_11061_));
 sky130_fd_sc_hd__nand3_2 _32699_ (.A(_11060_),
    .B(_11061_),
    .C(_11058_),
    .Y(_11062_));
 sky130_fd_sc_hd__buf_1 _32700_ (.A(_11062_),
    .X(_11063_));
 sky130_fd_sc_hd__buf_1 _32701_ (.A(_08990_),
    .X(_11064_));
 sky130_fd_sc_hd__and2_2 _32702_ (.A(_11064_),
    .B(_06924_),
    .X(_11065_));
 sky130_fd_sc_hd__nand2_2 _32703_ (.A(_08218_),
    .B(_07557_),
    .Y(_11066_));
 sky130_fd_sc_hd__buf_1 _32704_ (.A(_18770_),
    .X(_11067_));
 sky130_fd_sc_hd__nand2_2 _32705_ (.A(_11067_),
    .B(_07102_),
    .Y(_11068_));
 sky130_fd_sc_hd__xnor2_2 _32706_ (.A(_11066_),
    .B(_11068_),
    .Y(_11069_));
 sky130_fd_sc_hd__xor2_2 _32707_ (.A(_11065_),
    .B(_11069_),
    .X(_11070_));
 sky130_fd_sc_hd__nand2_2 _32708_ (.A(_18748_),
    .B(_06357_),
    .Y(_11071_));
 sky130_fd_sc_hd__nand2_2 _32709_ (.A(_09272_),
    .B(_06886_),
    .Y(_11072_));
 sky130_fd_sc_hd__nand2_2 _32710_ (.A(_11071_),
    .B(_11072_),
    .Y(_11073_));
 sky130_fd_sc_hd__buf_1 _32711_ (.A(_08731_),
    .X(_11074_));
 sky130_fd_sc_hd__nand3b_2 _32712_ (.A_N(_11071_),
    .B(_11074_),
    .C(_06197_),
    .Y(_11075_));
 sky130_fd_sc_hd__o2bb2ai_2 _32713_ (.A1_N(_11073_),
    .A2_N(_11075_),
    .B1(_18760_),
    .B2(_19243_),
    .Y(_11076_));
 sky130_fd_sc_hd__nor2_2 _32714_ (.A(_10731_),
    .B(_10732_),
    .Y(_11077_));
 sky130_fd_sc_hd__a21oi_2 _32715_ (.A1(_10733_),
    .A2(_10738_),
    .B1(_11077_),
    .Y(_11078_));
 sky130_vsdinv _32716_ (.A(_11078_),
    .Y(_11079_));
 sky130_fd_sc_hd__buf_1 _32717_ (.A(_08234_),
    .X(_11080_));
 sky130_fd_sc_hd__and2_2 _32718_ (.A(_11080_),
    .B(_06365_),
    .X(_11081_));
 sky130_fd_sc_hd__nand3_2 _32719_ (.A(_11075_),
    .B(_11081_),
    .C(_11073_),
    .Y(_11082_));
 sky130_fd_sc_hd__nand3_2 _32720_ (.A(_11076_),
    .B(_11079_),
    .C(_11082_),
    .Y(_11083_));
 sky130_fd_sc_hd__a21o_2 _32721_ (.A1(_11076_),
    .A2(_11082_),
    .B1(_11079_),
    .X(_11084_));
 sky130_fd_sc_hd__nand3b_2 _32722_ (.A_N(_11070_),
    .B(_11083_),
    .C(_11084_),
    .Y(_11085_));
 sky130_fd_sc_hd__nand2_2 _32723_ (.A(_11084_),
    .B(_11083_),
    .Y(_11086_));
 sky130_fd_sc_hd__nand2_2 _32724_ (.A(_11086_),
    .B(_11070_),
    .Y(_11087_));
 sky130_fd_sc_hd__nand2_2 _32725_ (.A(_10715_),
    .B(_10711_),
    .Y(_11088_));
 sky130_fd_sc_hd__a21oi_2 _32726_ (.A1(_11085_),
    .A2(_11087_),
    .B1(_11088_),
    .Y(_11089_));
 sky130_fd_sc_hd__nand3_2 _32727_ (.A(_11088_),
    .B(_11085_),
    .C(_11087_),
    .Y(_11090_));
 sky130_vsdinv _32728_ (.A(_11090_),
    .Y(_11091_));
 sky130_vsdinv _32729_ (.A(_10742_),
    .Y(_11092_));
 sky130_fd_sc_hd__a21oi_2 _32730_ (.A1(_10749_),
    .A2(_10741_),
    .B1(_11092_),
    .Y(_11093_));
 sky130_vsdinv _32731_ (.A(_11093_),
    .Y(_11094_));
 sky130_fd_sc_hd__o21bai_2 _32732_ (.A1(_11089_),
    .A2(_11091_),
    .B1_N(_11094_),
    .Y(_11095_));
 sky130_fd_sc_hd__nand3b_2 _32733_ (.A_N(_11089_),
    .B(_11094_),
    .C(_11090_),
    .Y(_11096_));
 sky130_fd_sc_hd__nand2_2 _32734_ (.A(_11095_),
    .B(_11096_),
    .Y(_11097_));
 sky130_fd_sc_hd__buf_1 _32735_ (.A(_11097_),
    .X(_11098_));
 sky130_fd_sc_hd__a21boi_2 _32736_ (.A1(_11059_),
    .A2(_11063_),
    .B1_N(_11098_),
    .Y(_11099_));
 sky130_fd_sc_hd__a21oi_2 _32737_ (.A1(_11060_),
    .A2(_11061_),
    .B1(_11058_),
    .Y(_11100_));
 sky130_fd_sc_hd__nor3b_2 _32738_ (.A(_11098_),
    .B(_11100_),
    .C_N(_11063_),
    .Y(_11101_));
 sky130_fd_sc_hd__o21ai_2 _32739_ (.A1(_10765_),
    .A2(_10766_),
    .B1(_10730_),
    .Y(_11102_));
 sky130_fd_sc_hd__o21bai_2 _32740_ (.A1(_11099_),
    .A2(_11101_),
    .B1_N(_11102_),
    .Y(_11103_));
 sky130_fd_sc_hd__nand2_2 _32741_ (.A(_11059_),
    .B(_11062_),
    .Y(_11104_));
 sky130_fd_sc_hd__nand2_2 _32742_ (.A(_11104_),
    .B(_11098_),
    .Y(_11105_));
 sky130_fd_sc_hd__nand3b_2 _32743_ (.A_N(_11097_),
    .B(_11059_),
    .C(_11063_),
    .Y(_11106_));
 sky130_fd_sc_hd__nand3_2 _32744_ (.A(_11105_),
    .B(_11106_),
    .C(_11102_),
    .Y(_11107_));
 sky130_fd_sc_hd__buf_1 _32745_ (.A(_07472_),
    .X(_11108_));
 sky130_fd_sc_hd__nand2_2 _32746_ (.A(_11108_),
    .B(_06735_),
    .Y(_11109_));
 sky130_fd_sc_hd__buf_1 _32747_ (.A(_07118_),
    .X(_11110_));
 sky130_fd_sc_hd__nand2_2 _32748_ (.A(_10774_),
    .B(_11110_),
    .Y(_11111_));
 sky130_fd_sc_hd__nand2_2 _32749_ (.A(_11109_),
    .B(_11111_),
    .Y(_11112_));
 sky130_fd_sc_hd__nand3b_2 _32750_ (.A_N(_11109_),
    .B(_18787_),
    .C(_11110_),
    .Y(_11113_));
 sky130_fd_sc_hd__o2bb2ai_2 _32751_ (.A1_N(_11112_),
    .A2_N(_11113_),
    .B1(_18793_),
    .B2(_19209_),
    .Y(_11114_));
 sky130_fd_sc_hd__and2_2 _32752_ (.A(_06667_),
    .B(_10379_),
    .X(_11115_));
 sky130_fd_sc_hd__nand3_2 _32753_ (.A(_11113_),
    .B(_11115_),
    .C(_11112_),
    .Y(_11116_));
 sky130_fd_sc_hd__nand2_2 _32754_ (.A(_10746_),
    .B(_10747_),
    .Y(_11117_));
 sky130_fd_sc_hd__nor2_2 _32755_ (.A(_10746_),
    .B(_10747_),
    .Y(_11118_));
 sky130_fd_sc_hd__a21oi_2 _32756_ (.A1(_11117_),
    .A2(_10744_),
    .B1(_11118_),
    .Y(_11119_));
 sky130_vsdinv _32757_ (.A(_11119_),
    .Y(_11120_));
 sky130_fd_sc_hd__a21oi_2 _32758_ (.A1(_11114_),
    .A2(_11116_),
    .B1(_11120_),
    .Y(_11121_));
 sky130_fd_sc_hd__nand3_2 _32759_ (.A(_11114_),
    .B(_11120_),
    .C(_11116_),
    .Y(_11122_));
 sky130_vsdinv _32760_ (.A(_11122_),
    .Y(_11123_));
 sky130_fd_sc_hd__a21boi_2 _32761_ (.A1(_10776_),
    .A2(_10782_),
    .B1_N(_10779_),
    .Y(_11124_));
 sky130_vsdinv _32762_ (.A(_11124_),
    .Y(_11125_));
 sky130_fd_sc_hd__o21bai_2 _32763_ (.A1(_11121_),
    .A2(_11123_),
    .B1_N(_11125_),
    .Y(_11126_));
 sky130_fd_sc_hd__nand3b_2 _32764_ (.A_N(_11121_),
    .B(_11125_),
    .C(_11122_),
    .Y(_11127_));
 sky130_fd_sc_hd__nand2_2 _32765_ (.A(_10792_),
    .B(_10788_),
    .Y(_11128_));
 sky130_fd_sc_hd__a21o_2 _32766_ (.A1(_11126_),
    .A2(_11127_),
    .B1(_11128_),
    .X(_11129_));
 sky130_fd_sc_hd__nand3_2 _32767_ (.A(_11128_),
    .B(_11126_),
    .C(_11127_),
    .Y(_11130_));
 sky130_fd_sc_hd__nand2_2 _32768_ (.A(_08169_),
    .B(_07966_),
    .Y(_11131_));
 sky130_fd_sc_hd__nand2_2 _32769_ (.A(_18802_),
    .B(_07591_),
    .Y(_11132_));
 sky130_fd_sc_hd__nand2_2 _32770_ (.A(_11131_),
    .B(_11132_),
    .Y(_11133_));
 sky130_fd_sc_hd__nand3b_2 _32771_ (.A_N(_11131_),
    .B(_06538_),
    .C(_08314_),
    .Y(_11134_));
 sky130_fd_sc_hd__o2bb2ai_2 _32772_ (.A1_N(_11133_),
    .A2_N(_11134_),
    .B1(_06692_),
    .B2(_19193_),
    .Y(_11135_));
 sky130_fd_sc_hd__buf_1 _32773_ (.A(_08569_),
    .X(_11136_));
 sky130_fd_sc_hd__and2_2 _32774_ (.A(_06550_),
    .B(_11136_),
    .X(_11137_));
 sky130_fd_sc_hd__nand3_2 _32775_ (.A(_11134_),
    .B(_11137_),
    .C(_11133_),
    .Y(_11138_));
 sky130_fd_sc_hd__nor2_2 _32776_ (.A(_10797_),
    .B(_10798_),
    .Y(_11139_));
 sky130_fd_sc_hd__a21oi_2 _32777_ (.A1(_10799_),
    .A2(_10802_),
    .B1(_11139_),
    .Y(_11140_));
 sky130_vsdinv _32778_ (.A(_11140_),
    .Y(_11141_));
 sky130_fd_sc_hd__a21oi_2 _32779_ (.A1(_11135_),
    .A2(_11138_),
    .B1(_11141_),
    .Y(_11142_));
 sky130_fd_sc_hd__nand3_2 _32780_ (.A(_11135_),
    .B(_11141_),
    .C(_11138_),
    .Y(_11143_));
 sky130_vsdinv _32781_ (.A(_11143_),
    .Y(_11144_));
 sky130_fd_sc_hd__and2_2 _32782_ (.A(_06136_),
    .B(_19171_),
    .X(_11145_));
 sky130_fd_sc_hd__buf_1 _32783_ (.A(_11145_),
    .X(_11146_));
 sky130_fd_sc_hd__nand2_2 _32784_ (.A(_06147_),
    .B(_08565_),
    .Y(_11147_));
 sky130_fd_sc_hd__nand2_2 _32785_ (.A(_06141_),
    .B(_19180_),
    .Y(_11148_));
 sky130_fd_sc_hd__xnor2_2 _32786_ (.A(_11147_),
    .B(_11148_),
    .Y(_11149_));
 sky130_fd_sc_hd__xor2_2 _32787_ (.A(_11146_),
    .B(_11149_),
    .X(_11150_));
 sky130_fd_sc_hd__o21ai_2 _32788_ (.A1(_11142_),
    .A2(_11144_),
    .B1(_11150_),
    .Y(_11151_));
 sky130_fd_sc_hd__xnor2_2 _32789_ (.A(_11146_),
    .B(_11149_),
    .Y(_11152_));
 sky130_fd_sc_hd__nand3b_2 _32790_ (.A_N(_11142_),
    .B(_11152_),
    .C(_11143_),
    .Y(_11153_));
 sky130_fd_sc_hd__nand2_2 _32791_ (.A(_11151_),
    .B(_11153_),
    .Y(_11154_));
 sky130_vsdinv _32792_ (.A(_11154_),
    .Y(_11155_));
 sky130_fd_sc_hd__a21oi_2 _32793_ (.A1(_11129_),
    .A2(_11130_),
    .B1(_11155_),
    .Y(_11156_));
 sky130_fd_sc_hd__nand3_2 _32794_ (.A(_11129_),
    .B(_11155_),
    .C(_11130_),
    .Y(_11157_));
 sky130_vsdinv _32795_ (.A(_11157_),
    .Y(_11158_));
 sky130_fd_sc_hd__a21boi_2 _32796_ (.A1(_10754_),
    .A2(_10758_),
    .B1_N(_10756_),
    .Y(_11159_));
 sky130_fd_sc_hd__o21ai_2 _32797_ (.A1(_11156_),
    .A2(_11158_),
    .B1(_11159_),
    .Y(_11160_));
 sky130_fd_sc_hd__nand2_2 _32798_ (.A(_10760_),
    .B(_10756_),
    .Y(_11161_));
 sky130_fd_sc_hd__a21o_2 _32799_ (.A1(_11129_),
    .A2(_11130_),
    .B1(_11155_),
    .X(_11162_));
 sky130_fd_sc_hd__nand3_2 _32800_ (.A(_11161_),
    .B(_11162_),
    .C(_11157_),
    .Y(_11163_));
 sky130_fd_sc_hd__buf_1 _32801_ (.A(_11163_),
    .X(_11164_));
 sky130_vsdinv _32802_ (.A(_10794_),
    .Y(_11165_));
 sky130_fd_sc_hd__a21oi_2 _32803_ (.A1(_10818_),
    .A2(_10796_),
    .B1(_11165_),
    .Y(_11166_));
 sky130_fd_sc_hd__buf_1 _32804_ (.A(_11166_),
    .X(_11167_));
 sky130_fd_sc_hd__a21boi_2 _32805_ (.A1(_11160_),
    .A2(_11164_),
    .B1_N(_11167_),
    .Y(_11168_));
 sky130_fd_sc_hd__a21oi_2 _32806_ (.A1(_11162_),
    .A2(_11157_),
    .B1(_11161_),
    .Y(_11169_));
 sky130_fd_sc_hd__nor3b_2 _32807_ (.A(_11167_),
    .B(_11169_),
    .C_N(_11164_),
    .Y(_11170_));
 sky130_fd_sc_hd__nor2_2 _32808_ (.A(_11168_),
    .B(_11170_),
    .Y(_11171_));
 sky130_fd_sc_hd__a21oi_2 _32809_ (.A1(_11103_),
    .A2(_11107_),
    .B1(_11171_),
    .Y(_11172_));
 sky130_fd_sc_hd__a21bo_2 _32810_ (.A1(_11160_),
    .A2(_11163_),
    .B1_N(_11167_),
    .X(_11173_));
 sky130_fd_sc_hd__nand3b_2 _32811_ (.A_N(_11166_),
    .B(_11160_),
    .C(_11164_),
    .Y(_11174_));
 sky130_fd_sc_hd__nand2_2 _32812_ (.A(_11173_),
    .B(_11174_),
    .Y(_11175_));
 sky130_fd_sc_hd__a21oi_2 _32813_ (.A1(_11105_),
    .A2(_11106_),
    .B1(_11102_),
    .Y(_11176_));
 sky130_vsdinv _32814_ (.A(_11107_),
    .Y(_11177_));
 sky130_fd_sc_hd__nor3_2 _32815_ (.A(_11175_),
    .B(_11176_),
    .C(_11177_),
    .Y(_11178_));
 sky130_fd_sc_hd__o21ai_2 _32816_ (.A1(_10833_),
    .A2(_10834_),
    .B1(_10773_),
    .Y(_11179_));
 sky130_fd_sc_hd__o21bai_2 _32817_ (.A1(_11172_),
    .A2(_11178_),
    .B1_N(_11179_),
    .Y(_11180_));
 sky130_fd_sc_hd__o22ai_2 _32818_ (.A1(_11170_),
    .A2(_11168_),
    .B1(_11176_),
    .B2(_11177_),
    .Y(_11181_));
 sky130_fd_sc_hd__nand3_2 _32819_ (.A(_11103_),
    .B(_11171_),
    .C(_11107_),
    .Y(_11182_));
 sky130_fd_sc_hd__nand3_2 _32820_ (.A(_11181_),
    .B(_11179_),
    .C(_11182_),
    .Y(_11183_));
 sky130_fd_sc_hd__buf_1 _32821_ (.A(_11183_),
    .X(_11184_));
 sky130_fd_sc_hd__nand2_2 _32822_ (.A(_07595_),
    .B(_10877_),
    .Y(_11185_));
 sky130_fd_sc_hd__nand2_2 _32823_ (.A(_05732_),
    .B(_10894_),
    .Y(_11186_));
 sky130_fd_sc_hd__nor2_2 _32824_ (.A(_11185_),
    .B(_11186_),
    .Y(_11187_));
 sky130_fd_sc_hd__buf_1 _32825_ (.A(_10882_),
    .X(_11188_));
 sky130_fd_sc_hd__nand2_2 _32826_ (.A(_11185_),
    .B(_11186_),
    .Y(_11189_));
 sky130_fd_sc_hd__nand3b_2 _32827_ (.A_N(_11187_),
    .B(_11188_),
    .C(_11189_),
    .Y(_11190_));
 sky130_vsdinv _32828_ (.A(_11187_),
    .Y(_11191_));
 sky130_fd_sc_hd__o2bb2ai_2 _32829_ (.A1_N(_11189_),
    .A2_N(_11191_),
    .B1(_16963_),
    .B2(_18881_),
    .Y(_11192_));
 sky130_fd_sc_hd__nor2_2 _32830_ (.A(_10876_),
    .B(_10878_),
    .Y(_11193_));
 sky130_fd_sc_hd__o21bai_2 _32831_ (.A1(_10888_),
    .A2(_10886_),
    .B1_N(_11193_),
    .Y(_11194_));
 sky130_fd_sc_hd__a21oi_2 _32832_ (.A1(_11190_),
    .A2(_11192_),
    .B1(_11194_),
    .Y(_11195_));
 sky130_fd_sc_hd__nand3_2 _32833_ (.A(_11194_),
    .B(_11190_),
    .C(_11192_),
    .Y(_11196_));
 sky130_vsdinv _32834_ (.A(_11196_),
    .Y(_11197_));
 sky130_fd_sc_hd__buf_1 _32835_ (.A(_19138_),
    .X(_11198_));
 sky130_fd_sc_hd__buf_1 _32836_ (.A(_11198_),
    .X(_11199_));
 sky130_fd_sc_hd__and2_2 _32837_ (.A(_05439_),
    .B(_11199_),
    .X(_11200_));
 sky130_fd_sc_hd__buf_1 _32838_ (.A(_10899_),
    .X(_11201_));
 sky130_fd_sc_hd__nand2_2 _32839_ (.A(_05422_),
    .B(_11201_),
    .Y(_11202_));
 sky130_fd_sc_hd__buf_1 _32840_ (.A(_16960_),
    .X(_11203_));
 sky130_fd_sc_hd__buf_1 _32841_ (.A(_11203_),
    .X(_11204_));
 sky130_fd_sc_hd__nand2_2 _32842_ (.A(_11204_),
    .B(_06363_),
    .Y(_11205_));
 sky130_fd_sc_hd__xnor2_2 _32843_ (.A(_11202_),
    .B(_11205_),
    .Y(_11206_));
 sky130_fd_sc_hd__xor2_2 _32844_ (.A(_11200_),
    .B(_11206_),
    .X(_11207_));
 sky130_fd_sc_hd__o21a_2 _32845_ (.A1(_11195_),
    .A2(_11197_),
    .B1(_11207_),
    .X(_11208_));
 sky130_fd_sc_hd__nor3b_2 _32846_ (.A(_11207_),
    .B(_11195_),
    .C_N(_11196_),
    .Y(_11209_));
 sky130_vsdinv _32847_ (.A(_11209_),
    .Y(_11210_));
 sky130_fd_sc_hd__a21boi_2 _32848_ (.A1(_10892_),
    .A2(_10903_),
    .B1_N(_10893_),
    .Y(_11211_));
 sky130_vsdinv _32849_ (.A(_11211_),
    .Y(_11212_));
 sky130_fd_sc_hd__nand3b_2 _32850_ (.A_N(_11208_),
    .B(_11210_),
    .C(_11212_),
    .Y(_11213_));
 sky130_fd_sc_hd__nor3_2 _32851_ (.A(_18859_),
    .B(_19147_),
    .C(_10902_),
    .Y(_11214_));
 sky130_fd_sc_hd__a41oi_2 _32852_ (.A1(_18869_),
    .A2(_05408_),
    .A3(_19137_),
    .A4(_10916_),
    .B1(_11214_),
    .Y(_11215_));
 sky130_vsdinv _32853_ (.A(_11215_),
    .Y(_11216_));
 sky130_fd_sc_hd__o21ai_2 _32854_ (.A1(_11209_),
    .A2(_11208_),
    .B1(_11211_),
    .Y(_11217_));
 sky130_fd_sc_hd__nand3_2 _32855_ (.A(_11213_),
    .B(_11216_),
    .C(_11217_),
    .Y(_11218_));
 sky130_vsdinv _32856_ (.A(_11218_),
    .Y(_11219_));
 sky130_fd_sc_hd__a21oi_2 _32857_ (.A1(_11213_),
    .A2(_11217_),
    .B1(_11216_),
    .Y(_11220_));
 sky130_fd_sc_hd__buf_1 _32858_ (.A(_09224_),
    .X(_11221_));
 sky130_fd_sc_hd__a22o_2 _32859_ (.A1(_06105_),
    .A2(_09786_),
    .B1(_05768_),
    .B2(_11221_),
    .X(_11222_));
 sky130_fd_sc_hd__nand2_2 _32860_ (.A(_18833_),
    .B(_09808_),
    .Y(_11223_));
 sky130_fd_sc_hd__buf_1 _32861_ (.A(_09086_),
    .X(_11224_));
 sky130_fd_sc_hd__nand3b_2 _32862_ (.A_N(_11223_),
    .B(_06225_),
    .C(_11224_),
    .Y(_11225_));
 sky130_fd_sc_hd__o2bb2ai_2 _32863_ (.A1_N(_11222_),
    .A2_N(_11225_),
    .B1(_18840_),
    .B2(_19157_),
    .Y(_11226_));
 sky130_fd_sc_hd__and2_2 _32864_ (.A(_06771_),
    .B(_09802_),
    .X(_11227_));
 sky130_fd_sc_hd__nand3_2 _32865_ (.A(_11225_),
    .B(_11222_),
    .C(_11227_),
    .Y(_11228_));
 sky130_fd_sc_hd__nand2_2 _32866_ (.A(_10809_),
    .B(_10810_),
    .Y(_11229_));
 sky130_fd_sc_hd__nor2_2 _32867_ (.A(_10809_),
    .B(_10810_),
    .Y(_11230_));
 sky130_fd_sc_hd__a21oi_2 _32868_ (.A1(_11229_),
    .A2(_10808_),
    .B1(_11230_),
    .Y(_11231_));
 sky130_vsdinv _32869_ (.A(_11231_),
    .Y(_11232_));
 sky130_fd_sc_hd__a21o_2 _32870_ (.A1(_11226_),
    .A2(_11228_),
    .B1(_11232_),
    .X(_11233_));
 sky130_fd_sc_hd__nand3_2 _32871_ (.A(_11226_),
    .B(_11232_),
    .C(_11228_),
    .Y(_11234_));
 sky130_fd_sc_hd__a21boi_2 _32872_ (.A1(_10845_),
    .A2(_10850_),
    .B1_N(_10847_),
    .Y(_11235_));
 sky130_fd_sc_hd__a21bo_2 _32873_ (.A1(_11233_),
    .A2(_11234_),
    .B1_N(_11235_),
    .X(_11236_));
 sky130_fd_sc_hd__nand3b_2 _32874_ (.A_N(_11235_),
    .B(_11233_),
    .C(_11234_),
    .Y(_11237_));
 sky130_fd_sc_hd__o21ai_2 _32875_ (.A1(_10807_),
    .A2(_10812_),
    .B1(_10813_),
    .Y(_11238_));
 sky130_fd_sc_hd__a21oi_2 _32876_ (.A1(_11236_),
    .A2(_11237_),
    .B1(_11238_),
    .Y(_11239_));
 sky130_fd_sc_hd__nand3_2 _32877_ (.A(_11236_),
    .B(_11238_),
    .C(_11237_),
    .Y(_11240_));
 sky130_vsdinv _32878_ (.A(_11240_),
    .Y(_11241_));
 sky130_vsdinv _32879_ (.A(_10857_),
    .Y(_11242_));
 sky130_fd_sc_hd__a21oi_2 _32880_ (.A1(_10856_),
    .A2(_10859_),
    .B1(_11242_),
    .Y(_11243_));
 sky130_vsdinv _32881_ (.A(_11243_),
    .Y(_11244_));
 sky130_fd_sc_hd__o21bai_2 _32882_ (.A1(_11239_),
    .A2(_11241_),
    .B1_N(_11244_),
    .Y(_11245_));
 sky130_fd_sc_hd__nand3b_2 _32883_ (.A_N(_11239_),
    .B(_11244_),
    .C(_11240_),
    .Y(_11246_));
 sky130_fd_sc_hd__nand2_2 _32884_ (.A(_10870_),
    .B(_10866_),
    .Y(_11247_));
 sky130_fd_sc_hd__a21oi_2 _32885_ (.A1(_11245_),
    .A2(_11246_),
    .B1(_11247_),
    .Y(_11248_));
 sky130_fd_sc_hd__nand3_2 _32886_ (.A(_11245_),
    .B(_11247_),
    .C(_11246_),
    .Y(_11249_));
 sky130_vsdinv _32887_ (.A(_11249_),
    .Y(_11250_));
 sky130_fd_sc_hd__o22ai_2 _32888_ (.A1(_11219_),
    .A2(_11220_),
    .B1(_11248_),
    .B2(_11250_),
    .Y(_11251_));
 sky130_fd_sc_hd__nor2_2 _32889_ (.A(_11220_),
    .B(_11219_),
    .Y(_11252_));
 sky130_fd_sc_hd__a21o_2 _32890_ (.A1(_11245_),
    .A2(_11246_),
    .B1(_11247_),
    .X(_11253_));
 sky130_fd_sc_hd__nand3_2 _32891_ (.A(_11252_),
    .B(_11249_),
    .C(_11253_),
    .Y(_11254_));
 sky130_fd_sc_hd__nand2_2 _32892_ (.A(_11251_),
    .B(_11254_),
    .Y(_11255_));
 sky130_fd_sc_hd__o21ai_2 _32893_ (.A1(_10824_),
    .A2(_10827_),
    .B1(_10823_),
    .Y(_11256_));
 sky130_vsdinv _32894_ (.A(_11256_),
    .Y(_11257_));
 sky130_fd_sc_hd__nand2_2 _32895_ (.A(_11255_),
    .B(_11257_),
    .Y(_11258_));
 sky130_fd_sc_hd__nand3_2 _32896_ (.A(_11251_),
    .B(_11256_),
    .C(_11254_),
    .Y(_11259_));
 sky130_fd_sc_hd__nand2_2 _32897_ (.A(_11258_),
    .B(_11259_),
    .Y(_11260_));
 sky130_fd_sc_hd__o21a_2 _32898_ (.A1(_10922_),
    .A2(_10924_),
    .B1(_10874_),
    .X(_11261_));
 sky130_fd_sc_hd__nand2_2 _32899_ (.A(_11260_),
    .B(_11261_),
    .Y(_11262_));
 sky130_fd_sc_hd__nand3b_2 _32900_ (.A_N(_11261_),
    .B(_11258_),
    .C(_11259_),
    .Y(_11263_));
 sky130_fd_sc_hd__nand2_2 _32901_ (.A(_11262_),
    .B(_11263_),
    .Y(_11264_));
 sky130_fd_sc_hd__buf_1 _32902_ (.A(_11264_),
    .X(_11265_));
 sky130_fd_sc_hd__a21boi_2 _32903_ (.A1(_11180_),
    .A2(_11184_),
    .B1_N(_11265_),
    .Y(_11266_));
 sky130_fd_sc_hd__a21oi_2 _32904_ (.A1(_11181_),
    .A2(_11182_),
    .B1(_11179_),
    .Y(_11267_));
 sky130_fd_sc_hd__nor3b_2 _32905_ (.A(_11265_),
    .B(_11267_),
    .C_N(_11184_),
    .Y(_11268_));
 sky130_fd_sc_hd__o21ai_2 _32906_ (.A1(_10941_),
    .A2(_10942_),
    .B1(_10842_),
    .Y(_11269_));
 sky130_fd_sc_hd__o21bai_2 _32907_ (.A1(_11266_),
    .A2(_11268_),
    .B1_N(_11269_),
    .Y(_11270_));
 sky130_fd_sc_hd__nand2_2 _32908_ (.A(_11180_),
    .B(_11183_),
    .Y(_11271_));
 sky130_fd_sc_hd__nand2_2 _32909_ (.A(_11271_),
    .B(_11265_),
    .Y(_11272_));
 sky130_fd_sc_hd__nand3b_2 _32910_ (.A_N(_11264_),
    .B(_11184_),
    .C(_11180_),
    .Y(_11273_));
 sky130_fd_sc_hd__nand3_2 _32911_ (.A(_11272_),
    .B(_11273_),
    .C(_11269_),
    .Y(_11274_));
 sky130_fd_sc_hd__nand2_2 _32912_ (.A(_11270_),
    .B(_11274_),
    .Y(_11275_));
 sky130_fd_sc_hd__and2_2 _32913_ (.A(_10920_),
    .B(_10909_),
    .X(_11276_));
 sky130_fd_sc_hd__o21a_2 _32914_ (.A1(_10933_),
    .A2(_10935_),
    .B1(_10931_),
    .X(_11277_));
 sky130_fd_sc_hd__xor2_2 _32915_ (.A(_11276_),
    .B(_11277_),
    .X(_11278_));
 sky130_vsdinv _32916_ (.A(_11278_),
    .Y(_11279_));
 sky130_fd_sc_hd__nand2_2 _32917_ (.A(_11275_),
    .B(_11279_),
    .Y(_11280_));
 sky130_fd_sc_hd__nand3_2 _32918_ (.A(_11270_),
    .B(_11278_),
    .C(_11274_),
    .Y(_11281_));
 sky130_fd_sc_hd__nor3_2 _32919_ (.A(_10945_),
    .B(_10938_),
    .C(_10944_),
    .Y(_11282_));
 sky130_fd_sc_hd__a21o_2 _32920_ (.A1(_10948_),
    .A2(_10957_),
    .B1(_11282_),
    .X(_11283_));
 sky130_fd_sc_hd__a21oi_2 _32921_ (.A1(_11280_),
    .A2(_11281_),
    .B1(_11283_),
    .Y(_11284_));
 sky130_fd_sc_hd__a21oi_2 _32922_ (.A1(_10948_),
    .A2(_10957_),
    .B1(_11282_),
    .Y(_11285_));
 sky130_fd_sc_hd__a21oi_2 _32923_ (.A1(_11270_),
    .A2(_11274_),
    .B1(_11278_),
    .Y(_11286_));
 sky130_vsdinv _32924_ (.A(_11281_),
    .Y(_11287_));
 sky130_fd_sc_hd__nor3_2 _32925_ (.A(_11285_),
    .B(_11286_),
    .C(_11287_),
    .Y(_11288_));
 sky130_fd_sc_hd__buf_1 _32926_ (.A(_10672_),
    .X(_11289_));
 sky130_fd_sc_hd__buf_1 _32927_ (.A(_11289_),
    .X(_11290_));
 sky130_fd_sc_hd__buf_1 _32928_ (.A(_11290_),
    .X(_11291_));
 sky130_fd_sc_hd__a21boi_2 _32929_ (.A1(_11291_),
    .A2(_10954_),
    .B1_N(_10953_),
    .Y(_11292_));
 sky130_vsdinv _32930_ (.A(_11292_),
    .Y(_11293_));
 sky130_fd_sc_hd__o21bai_2 _32931_ (.A1(_11284_),
    .A2(_11288_),
    .B1_N(_11293_),
    .Y(_11294_));
 sky130_fd_sc_hd__o21ai_2 _32932_ (.A1(_11286_),
    .A2(_11287_),
    .B1(_11285_),
    .Y(_11295_));
 sky130_fd_sc_hd__nand3_2 _32933_ (.A(_11283_),
    .B(_11280_),
    .C(_11281_),
    .Y(_11296_));
 sky130_fd_sc_hd__nand3_2 _32934_ (.A(_11295_),
    .B(_11293_),
    .C(_11296_),
    .Y(_11297_));
 sky130_vsdinv _32935_ (.A(_10965_),
    .Y(_11298_));
 sky130_fd_sc_hd__a21oi_2 _32936_ (.A1(_10963_),
    .A2(_10959_),
    .B1(_10961_),
    .Y(_11299_));
 sky130_fd_sc_hd__o21ai_2 _32937_ (.A1(_11298_),
    .A2(_11299_),
    .B1(_10964_),
    .Y(_11300_));
 sky130_fd_sc_hd__a21o_2 _32938_ (.A1(_11294_),
    .A2(_11297_),
    .B1(_11300_),
    .X(_11301_));
 sky130_fd_sc_hd__nand3_2 _32939_ (.A(_11294_),
    .B(_11300_),
    .C(_11297_),
    .Y(_11302_));
 sky130_fd_sc_hd__nand2_2 _32940_ (.A(_11301_),
    .B(_11302_),
    .Y(_11303_));
 sky130_fd_sc_hd__a21boi_2 _32941_ (.A1(_10993_),
    .A2(_10969_),
    .B1_N(_10970_),
    .Y(_11304_));
 sky130_fd_sc_hd__xor2_2 _32942_ (.A(_11303_),
    .B(_11304_),
    .X(_02652_));
 sky130_fd_sc_hd__nand2_2 _32943_ (.A(_18727_),
    .B(_07375_),
    .Y(_11305_));
 sky130_fd_sc_hd__nand2_2 _32944_ (.A(_09589_),
    .B(_07216_),
    .Y(_11306_));
 sky130_fd_sc_hd__xor2_2 _32945_ (.A(_11305_),
    .B(_11306_),
    .X(_11307_));
 sky130_fd_sc_hd__and2_2 _32946_ (.A(_08457_),
    .B(_05935_),
    .X(_11308_));
 sky130_fd_sc_hd__nand2_2 _32947_ (.A(_11307_),
    .B(_11308_),
    .Y(_11309_));
 sky130_fd_sc_hd__xnor2_2 _32948_ (.A(_11305_),
    .B(_11306_),
    .Y(_11310_));
 sky130_fd_sc_hd__o21ai_2 _32949_ (.A1(_09011_),
    .A2(_19253_),
    .B1(_11310_),
    .Y(_11311_));
 sky130_fd_sc_hd__nand2_2 _32950_ (.A(_11309_),
    .B(_11311_),
    .Y(_11312_));
 sky130_fd_sc_hd__a21oi_2 _32951_ (.A1(_11017_),
    .A2(_11013_),
    .B1(_11012_),
    .Y(_11313_));
 sky130_fd_sc_hd__nand2_2 _32952_ (.A(_11312_),
    .B(_11313_),
    .Y(_11314_));
 sky130_fd_sc_hd__nor2_2 _32953_ (.A(_11031_),
    .B(_11032_),
    .Y(_11315_));
 sky130_fd_sc_hd__a21oi_2 _32954_ (.A1(_11033_),
    .A2(_11034_),
    .B1(_11315_),
    .Y(_11316_));
 sky130_vsdinv _32955_ (.A(_11316_),
    .Y(_11317_));
 sky130_fd_sc_hd__nand3b_2 _32956_ (.A_N(_11313_),
    .B(_11309_),
    .C(_11311_),
    .Y(_11318_));
 sky130_fd_sc_hd__nand3_2 _32957_ (.A(_11314_),
    .B(_11317_),
    .C(_11318_),
    .Y(_11319_));
 sky130_fd_sc_hd__a21o_2 _32958_ (.A1(_11314_),
    .A2(_11318_),
    .B1(_11317_),
    .X(_11320_));
 sky130_fd_sc_hd__nand2_2 _32959_ (.A(_10994_),
    .B(_07171_),
    .Y(_11321_));
 sky130_fd_sc_hd__buf_1 _32960_ (.A(_10671_),
    .X(_11322_));
 sky130_fd_sc_hd__nand3b_2 _32961_ (.A_N(_11321_),
    .B(_11322_),
    .C(_19294_),
    .Y(_11323_));
 sky130_fd_sc_hd__buf_1 _32962_ (.A(_16968_),
    .X(_11324_));
 sky130_fd_sc_hd__o21ai_2 _32963_ (.A1(_07013_),
    .A2(_11324_),
    .B1(_11321_),
    .Y(_11325_));
 sky130_fd_sc_hd__buf_1 _32964_ (.A(_10266_),
    .X(_11326_));
 sky130_fd_sc_hd__and2_2 _32965_ (.A(_11326_),
    .B(_07794_),
    .X(_11327_));
 sky130_fd_sc_hd__a21oi_2 _32966_ (.A1(_11323_),
    .A2(_11325_),
    .B1(_11327_),
    .Y(_11328_));
 sky130_fd_sc_hd__nand3_2 _32967_ (.A(_11323_),
    .B(_11327_),
    .C(_11325_),
    .Y(_11329_));
 sky130_vsdinv _32968_ (.A(_11329_),
    .Y(_11330_));
 sky130_fd_sc_hd__buf_1 _32969_ (.A(_16967_),
    .X(_11331_));
 sky130_fd_sc_hd__buf_1 _32970_ (.A(_11331_),
    .X(_11332_));
 sky130_fd_sc_hd__nor3_2 _32971_ (.A(_06144_),
    .B(_11332_),
    .C(_10995_),
    .Y(_11333_));
 sky130_fd_sc_hd__a21o_2 _32972_ (.A1(_10999_),
    .A2(_11000_),
    .B1(_11333_),
    .X(_11334_));
 sky130_fd_sc_hd__o21bai_2 _32973_ (.A1(_11328_),
    .A2(_11330_),
    .B1_N(_11334_),
    .Y(_11335_));
 sky130_fd_sc_hd__a21o_2 _32974_ (.A1(_11323_),
    .A2(_11325_),
    .B1(_11327_),
    .X(_11336_));
 sky130_fd_sc_hd__nand3_2 _32975_ (.A(_11336_),
    .B(_11334_),
    .C(_11329_),
    .Y(_11337_));
 sky130_fd_sc_hd__buf_1 _32976_ (.A(_09957_),
    .X(_11338_));
 sky130_fd_sc_hd__a22oi_2 _32977_ (.A1(_11338_),
    .A2(_06820_),
    .B1(_09603_),
    .B2(_06041_),
    .Y(_11339_));
 sky130_fd_sc_hd__buf_1 _32978_ (.A(_18716_),
    .X(_11340_));
 sky130_fd_sc_hd__and4_2 _32979_ (.A(_10683_),
    .B(_11340_),
    .C(_05931_),
    .D(_05927_),
    .X(_11341_));
 sky130_fd_sc_hd__and2_2 _32980_ (.A(_10474_),
    .B(_08007_),
    .X(_11342_));
 sky130_fd_sc_hd__o21bai_2 _32981_ (.A1(_11339_),
    .A2(_11341_),
    .B1_N(_11342_),
    .Y(_11343_));
 sky130_fd_sc_hd__nand2_2 _32982_ (.A(_11338_),
    .B(_06991_),
    .Y(_11344_));
 sky130_fd_sc_hd__nand3b_2 _32983_ (.A_N(_11344_),
    .B(_10263_),
    .C(_19273_),
    .Y(_11345_));
 sky130_fd_sc_hd__nand3b_2 _32984_ (.A_N(_11339_),
    .B(_11345_),
    .C(_11342_),
    .Y(_11346_));
 sky130_fd_sc_hd__nand2_2 _32985_ (.A(_11343_),
    .B(_11346_),
    .Y(_11347_));
 sky130_vsdinv _32986_ (.A(_11347_),
    .Y(_11348_));
 sky130_fd_sc_hd__a21oi_2 _32987_ (.A1(_11335_),
    .A2(_11337_),
    .B1(_11348_),
    .Y(_11349_));
 sky130_fd_sc_hd__nand3_2 _32988_ (.A(_11335_),
    .B(_11348_),
    .C(_11337_),
    .Y(_11350_));
 sky130_vsdinv _32989_ (.A(_11350_),
    .Y(_11351_));
 sky130_fd_sc_hd__a21oi_2 _32990_ (.A1(_11009_),
    .A2(_11002_),
    .B1(_11007_),
    .Y(_11352_));
 sky130_fd_sc_hd__o21ai_2 _32991_ (.A1(_11020_),
    .A2(_11352_),
    .B1(_11010_),
    .Y(_11353_));
 sky130_fd_sc_hd__o21bai_2 _32992_ (.A1(_11349_),
    .A2(_11351_),
    .B1_N(_11353_),
    .Y(_11354_));
 sky130_fd_sc_hd__a21o_2 _32993_ (.A1(_11335_),
    .A2(_11337_),
    .B1(_11348_),
    .X(_11355_));
 sky130_fd_sc_hd__nand3_2 _32994_ (.A(_11355_),
    .B(_11350_),
    .C(_11353_),
    .Y(_11356_));
 sky130_fd_sc_hd__a22oi_2 _32995_ (.A1(_11319_),
    .A2(_11320_),
    .B1(_11354_),
    .B2(_11356_),
    .Y(_11357_));
 sky130_fd_sc_hd__nand2_2 _32996_ (.A(_11320_),
    .B(_11319_),
    .Y(_11358_));
 sky130_fd_sc_hd__nand2_2 _32997_ (.A(_11354_),
    .B(_11356_),
    .Y(_11359_));
 sky130_fd_sc_hd__nor2_2 _32998_ (.A(_11358_),
    .B(_11359_),
    .Y(_11360_));
 sky130_fd_sc_hd__o21ai_2 _32999_ (.A1(_11054_),
    .A2(_11055_),
    .B1(_11028_),
    .Y(_11361_));
 sky130_fd_sc_hd__o21bai_2 _33000_ (.A1(_11357_),
    .A2(_11360_),
    .B1_N(_11361_),
    .Y(_11362_));
 sky130_fd_sc_hd__nand2_2 _33001_ (.A(_11359_),
    .B(_11358_),
    .Y(_11363_));
 sky130_fd_sc_hd__nand3b_2 _33002_ (.A_N(_11358_),
    .B(_11356_),
    .C(_11354_),
    .Y(_11364_));
 sky130_fd_sc_hd__nand3_2 _33003_ (.A(_11363_),
    .B(_11361_),
    .C(_11364_),
    .Y(_11365_));
 sky130_fd_sc_hd__nand2_2 _33004_ (.A(_08729_),
    .B(_07515_),
    .Y(_11366_));
 sky130_fd_sc_hd__nand2_2 _33005_ (.A(_09266_),
    .B(_06728_),
    .Y(_11367_));
 sky130_fd_sc_hd__nand2_2 _33006_ (.A(_11366_),
    .B(_11367_),
    .Y(_11368_));
 sky130_fd_sc_hd__nand3b_2 _33007_ (.A_N(_11366_),
    .B(_11074_),
    .C(_06464_),
    .Y(_11369_));
 sky130_fd_sc_hd__o2bb2ai_2 _33008_ (.A1_N(_11368_),
    .A2_N(_11369_),
    .B1(_18760_),
    .B2(_19238_),
    .Y(_11370_));
 sky130_fd_sc_hd__and2_2 _33009_ (.A(_08235_),
    .B(_06466_),
    .X(_11371_));
 sky130_fd_sc_hd__nand3_2 _33010_ (.A(_11369_),
    .B(_11371_),
    .C(_11368_),
    .Y(_11372_));
 sky130_fd_sc_hd__nor2_2 _33011_ (.A(_11071_),
    .B(_11072_),
    .Y(_11373_));
 sky130_fd_sc_hd__a21oi_2 _33012_ (.A1(_11073_),
    .A2(_11081_),
    .B1(_11373_),
    .Y(_11374_));
 sky130_vsdinv _33013_ (.A(_11374_),
    .Y(_11375_));
 sky130_fd_sc_hd__a21o_2 _33014_ (.A1(_11370_),
    .A2(_11372_),
    .B1(_11375_),
    .X(_11376_));
 sky130_fd_sc_hd__nand3_2 _33015_ (.A(_11370_),
    .B(_11375_),
    .C(_11372_),
    .Y(_11377_));
 sky130_fd_sc_hd__and2_2 _33016_ (.A(_11064_),
    .B(_10150_),
    .X(_11378_));
 sky130_fd_sc_hd__nand2_2 _33017_ (.A(_08218_),
    .B(_07102_),
    .Y(_11379_));
 sky130_fd_sc_hd__nand2_2 _33018_ (.A(_11067_),
    .B(_08256_),
    .Y(_11380_));
 sky130_fd_sc_hd__xnor2_2 _33019_ (.A(_11379_),
    .B(_11380_),
    .Y(_11381_));
 sky130_fd_sc_hd__xnor2_2 _33020_ (.A(_11378_),
    .B(_11381_),
    .Y(_11382_));
 sky130_fd_sc_hd__a21oi_2 _33021_ (.A1(_11376_),
    .A2(_11377_),
    .B1(_11382_),
    .Y(_11383_));
 sky130_fd_sc_hd__nand3_2 _33022_ (.A(_11382_),
    .B(_11376_),
    .C(_11377_),
    .Y(_11384_));
 sky130_vsdinv _33023_ (.A(_11384_),
    .Y(_11385_));
 sky130_fd_sc_hd__o21ai_2 _33024_ (.A1(_11044_),
    .A2(_11051_),
    .B1(_11041_),
    .Y(_11386_));
 sky130_fd_sc_hd__o21bai_2 _33025_ (.A1(_11383_),
    .A2(_11385_),
    .B1_N(_11386_),
    .Y(_11387_));
 sky130_fd_sc_hd__a21o_2 _33026_ (.A1(_11376_),
    .A2(_11377_),
    .B1(_11382_),
    .X(_11388_));
 sky130_fd_sc_hd__nand3_2 _33027_ (.A(_11388_),
    .B(_11386_),
    .C(_11384_),
    .Y(_11389_));
 sky130_fd_sc_hd__buf_1 _33028_ (.A(_11389_),
    .X(_11390_));
 sky130_fd_sc_hd__o21a_2 _33029_ (.A1(_11070_),
    .A2(_11086_),
    .B1(_11083_),
    .X(_11391_));
 sky130_vsdinv _33030_ (.A(_11391_),
    .Y(_11392_));
 sky130_fd_sc_hd__a21oi_2 _33031_ (.A1(_11387_),
    .A2(_11390_),
    .B1(_11392_),
    .Y(_11393_));
 sky130_fd_sc_hd__a21oi_2 _33032_ (.A1(_11388_),
    .A2(_11384_),
    .B1(_11386_),
    .Y(_11394_));
 sky130_fd_sc_hd__nor3b_2 _33033_ (.A(_11391_),
    .B(_11394_),
    .C_N(_11390_),
    .Y(_11395_));
 sky130_fd_sc_hd__nor2_2 _33034_ (.A(_11393_),
    .B(_11395_),
    .Y(_11396_));
 sky130_fd_sc_hd__a21oi_2 _33035_ (.A1(_11362_),
    .A2(_11365_),
    .B1(_11396_),
    .Y(_11397_));
 sky130_fd_sc_hd__nand3_2 _33036_ (.A(_11362_),
    .B(_11396_),
    .C(_11365_),
    .Y(_11398_));
 sky130_vsdinv _33037_ (.A(_11398_),
    .Y(_11399_));
 sky130_fd_sc_hd__o21ai_2 _33038_ (.A1(_11098_),
    .A2(_11100_),
    .B1(_11063_),
    .Y(_11400_));
 sky130_fd_sc_hd__o21bai_2 _33039_ (.A1(_11397_),
    .A2(_11399_),
    .B1_N(_11400_),
    .Y(_11401_));
 sky130_fd_sc_hd__a21oi_2 _33040_ (.A1(_11363_),
    .A2(_11364_),
    .B1(_11361_),
    .Y(_11402_));
 sky130_vsdinv _33041_ (.A(_11365_),
    .Y(_11403_));
 sky130_fd_sc_hd__o21bai_2 _33042_ (.A1(_11402_),
    .A2(_11403_),
    .B1_N(_11396_),
    .Y(_11404_));
 sky130_fd_sc_hd__nand3_2 _33043_ (.A(_11404_),
    .B(_11400_),
    .C(_11398_),
    .Y(_11405_));
 sky130_fd_sc_hd__nand2_2 _33044_ (.A(_10356_),
    .B(_07737_),
    .Y(_11406_));
 sky130_fd_sc_hd__nand2_2 _33045_ (.A(_07395_),
    .B(_07944_),
    .Y(_11407_));
 sky130_fd_sc_hd__xor2_2 _33046_ (.A(_11406_),
    .B(_11407_),
    .X(_11408_));
 sky130_fd_sc_hd__buf_1 _33047_ (.A(_06666_),
    .X(_11409_));
 sky130_fd_sc_hd__and2_2 _33048_ (.A(_11409_),
    .B(_07967_),
    .X(_11410_));
 sky130_fd_sc_hd__nand2_2 _33049_ (.A(_11408_),
    .B(_11410_),
    .Y(_11411_));
 sky130_fd_sc_hd__xnor2_2 _33050_ (.A(_11406_),
    .B(_11407_),
    .Y(_11412_));
 sky130_fd_sc_hd__o21ai_2 _33051_ (.A1(_07400_),
    .A2(_19205_),
    .B1(_11412_),
    .Y(_11413_));
 sky130_fd_sc_hd__nand2_2 _33052_ (.A(_11066_),
    .B(_11068_),
    .Y(_11414_));
 sky130_fd_sc_hd__nor2_2 _33053_ (.A(_11066_),
    .B(_11068_),
    .Y(_11415_));
 sky130_fd_sc_hd__a21oi_2 _33054_ (.A1(_11414_),
    .A2(_11065_),
    .B1(_11415_),
    .Y(_11416_));
 sky130_vsdinv _33055_ (.A(_11416_),
    .Y(_11417_));
 sky130_fd_sc_hd__a21oi_2 _33056_ (.A1(_11411_),
    .A2(_11413_),
    .B1(_11417_),
    .Y(_11418_));
 sky130_fd_sc_hd__nand3_2 _33057_ (.A(_11411_),
    .B(_11413_),
    .C(_11417_),
    .Y(_11419_));
 sky130_vsdinv _33058_ (.A(_11419_),
    .Y(_11420_));
 sky130_fd_sc_hd__a21boi_2 _33059_ (.A1(_11115_),
    .A2(_11112_),
    .B1_N(_11113_),
    .Y(_11421_));
 sky130_vsdinv _33060_ (.A(_11421_),
    .Y(_11422_));
 sky130_fd_sc_hd__o21bai_2 _33061_ (.A1(_11418_),
    .A2(_11420_),
    .B1_N(_11422_),
    .Y(_11423_));
 sky130_fd_sc_hd__a21o_2 _33062_ (.A1(_11411_),
    .A2(_11413_),
    .B1(_11417_),
    .X(_11424_));
 sky130_fd_sc_hd__nand3_2 _33063_ (.A(_11424_),
    .B(_11422_),
    .C(_11419_),
    .Y(_11425_));
 sky130_fd_sc_hd__o21ai_2 _33064_ (.A1(_11124_),
    .A2(_11121_),
    .B1(_11122_),
    .Y(_11426_));
 sky130_fd_sc_hd__a21oi_2 _33065_ (.A1(_11423_),
    .A2(_11425_),
    .B1(_11426_),
    .Y(_11427_));
 sky130_fd_sc_hd__nand3_2 _33066_ (.A(_11423_),
    .B(_11426_),
    .C(_11425_),
    .Y(_11428_));
 sky130_vsdinv _33067_ (.A(_11428_),
    .Y(_11429_));
 sky130_fd_sc_hd__and2_2 _33068_ (.A(_06816_),
    .B(_11224_),
    .X(_11430_));
 sky130_fd_sc_hd__a22oi_2 _33069_ (.A1(_10393_),
    .A2(_08830_),
    .B1(_06674_),
    .B2(_08833_),
    .Y(_11431_));
 sky130_fd_sc_hd__buf_1 _33070_ (.A(_07377_),
    .X(_11432_));
 sky130_fd_sc_hd__buf_1 _33071_ (.A(_08556_),
    .X(_11433_));
 sky130_fd_sc_hd__buf_1 _33072_ (.A(_08829_),
    .X(_11434_));
 sky130_fd_sc_hd__and4_2 _33073_ (.A(_10393_),
    .B(_11432_),
    .C(_11433_),
    .D(_11434_),
    .X(_11435_));
 sky130_fd_sc_hd__nor2_2 _33074_ (.A(_11431_),
    .B(_11435_),
    .Y(_11436_));
 sky130_fd_sc_hd__xnor2_2 _33075_ (.A(_11430_),
    .B(_11436_),
    .Y(_11437_));
 sky130_fd_sc_hd__nand2_2 _33076_ (.A(_08169_),
    .B(_08812_),
    .Y(_11438_));
 sky130_fd_sc_hd__nand2_2 _33077_ (.A(_09870_),
    .B(_11136_),
    .Y(_11439_));
 sky130_fd_sc_hd__nand2_2 _33078_ (.A(_11438_),
    .B(_11439_),
    .Y(_11440_));
 sky130_fd_sc_hd__buf_1 _33079_ (.A(_08570_),
    .X(_11441_));
 sky130_fd_sc_hd__nand3b_2 _33080_ (.A_N(_11438_),
    .B(_08043_),
    .C(_11441_),
    .Y(_11442_));
 sky130_fd_sc_hd__o2bb2ai_2 _33081_ (.A1_N(_11440_),
    .A2_N(_11442_),
    .B1(_18810_),
    .B2(_19187_),
    .Y(_11443_));
 sky130_fd_sc_hd__and2_2 _33082_ (.A(_08039_),
    .B(_09216_),
    .X(_11444_));
 sky130_fd_sc_hd__nand3_2 _33083_ (.A(_11442_),
    .B(_11444_),
    .C(_11440_),
    .Y(_11445_));
 sky130_fd_sc_hd__nor2_2 _33084_ (.A(_11131_),
    .B(_11132_),
    .Y(_11446_));
 sky130_fd_sc_hd__a21oi_2 _33085_ (.A1(_11133_),
    .A2(_11137_),
    .B1(_11446_),
    .Y(_11447_));
 sky130_vsdinv _33086_ (.A(_11447_),
    .Y(_11448_));
 sky130_fd_sc_hd__a21o_2 _33087_ (.A1(_11443_),
    .A2(_11445_),
    .B1(_11448_),
    .X(_11449_));
 sky130_fd_sc_hd__nand3_2 _33088_ (.A(_11443_),
    .B(_11448_),
    .C(_11445_),
    .Y(_11450_));
 sky130_fd_sc_hd__nand2_2 _33089_ (.A(_11449_),
    .B(_11450_),
    .Y(_11451_));
 sky130_fd_sc_hd__xor2_2 _33090_ (.A(_11437_),
    .B(_11451_),
    .X(_11452_));
 sky130_fd_sc_hd__o21bai_2 _33091_ (.A1(_11427_),
    .A2(_11429_),
    .B1_N(_11452_),
    .Y(_11453_));
 sky130_fd_sc_hd__a21o_2 _33092_ (.A1(_11423_),
    .A2(_11425_),
    .B1(_11426_),
    .X(_11454_));
 sky130_fd_sc_hd__nand3_2 _33093_ (.A(_11454_),
    .B(_11452_),
    .C(_11428_),
    .Y(_11455_));
 sky130_fd_sc_hd__o21ai_2 _33094_ (.A1(_11093_),
    .A2(_11089_),
    .B1(_11090_),
    .Y(_11456_));
 sky130_fd_sc_hd__a21o_2 _33095_ (.A1(_11453_),
    .A2(_11455_),
    .B1(_11456_),
    .X(_11457_));
 sky130_fd_sc_hd__nand3_2 _33096_ (.A(_11453_),
    .B(_11456_),
    .C(_11455_),
    .Y(_11458_));
 sky130_vsdinv _33097_ (.A(_11130_),
    .Y(_11459_));
 sky130_fd_sc_hd__a21oi_2 _33098_ (.A1(_11129_),
    .A2(_11155_),
    .B1(_11459_),
    .Y(_11460_));
 sky130_vsdinv _33099_ (.A(_11460_),
    .Y(_11461_));
 sky130_fd_sc_hd__a21oi_2 _33100_ (.A1(_11457_),
    .A2(_11458_),
    .B1(_11461_),
    .Y(_11462_));
 sky130_fd_sc_hd__nand3_2 _33101_ (.A(_11457_),
    .B(_11461_),
    .C(_11458_),
    .Y(_11463_));
 sky130_vsdinv _33102_ (.A(_11463_),
    .Y(_11464_));
 sky130_fd_sc_hd__nor2_2 _33103_ (.A(_11462_),
    .B(_11464_),
    .Y(_11465_));
 sky130_fd_sc_hd__a21oi_2 _33104_ (.A1(_11401_),
    .A2(_11405_),
    .B1(_11465_),
    .Y(_11466_));
 sky130_fd_sc_hd__a21oi_2 _33105_ (.A1(_11453_),
    .A2(_11455_),
    .B1(_11456_),
    .Y(_11467_));
 sky130_vsdinv _33106_ (.A(_11458_),
    .Y(_11468_));
 sky130_fd_sc_hd__o21bai_2 _33107_ (.A1(_11467_),
    .A2(_11468_),
    .B1_N(_11461_),
    .Y(_11469_));
 sky130_fd_sc_hd__nand2_2 _33108_ (.A(_11469_),
    .B(_11463_),
    .Y(_11470_));
 sky130_fd_sc_hd__a21oi_2 _33109_ (.A1(_11404_),
    .A2(_11398_),
    .B1(_11400_),
    .Y(_11471_));
 sky130_vsdinv _33110_ (.A(_11405_),
    .Y(_11472_));
 sky130_fd_sc_hd__nor3_2 _33111_ (.A(_11470_),
    .B(_11471_),
    .C(_11472_),
    .Y(_11473_));
 sky130_fd_sc_hd__o21ai_2 _33112_ (.A1(_11175_),
    .A2(_11176_),
    .B1(_11107_),
    .Y(_11474_));
 sky130_fd_sc_hd__o21bai_2 _33113_ (.A1(_11466_),
    .A2(_11473_),
    .B1_N(_11474_),
    .Y(_11475_));
 sky130_fd_sc_hd__o22ai_2 _33114_ (.A1(_11464_),
    .A2(_11462_),
    .B1(_11471_),
    .B2(_11472_),
    .Y(_11476_));
 sky130_fd_sc_hd__nand3_2 _33115_ (.A(_11465_),
    .B(_11401_),
    .C(_11405_),
    .Y(_11477_));
 sky130_fd_sc_hd__nand3_2 _33116_ (.A(_11476_),
    .B(_11474_),
    .C(_11477_),
    .Y(_11478_));
 sky130_fd_sc_hd__buf_1 _33117_ (.A(_11478_),
    .X(_11479_));
 sky130_fd_sc_hd__nand2_2 _33118_ (.A(_05926_),
    .B(_10555_),
    .Y(_11480_));
 sky130_fd_sc_hd__nand2_2 _33119_ (.A(_05816_),
    .B(_10912_),
    .Y(_11481_));
 sky130_fd_sc_hd__nor2_2 _33120_ (.A(_11480_),
    .B(_11481_),
    .Y(_11482_));
 sky130_fd_sc_hd__nand2_2 _33121_ (.A(_11480_),
    .B(_11481_),
    .Y(_11483_));
 sky130_fd_sc_hd__nor3b_2 _33122_ (.A(_11482_),
    .B(_10887_),
    .C_N(_11483_),
    .Y(_11484_));
 sky130_vsdinv _33123_ (.A(_11484_),
    .Y(_11485_));
 sky130_vsdinv _33124_ (.A(_11482_),
    .Y(_11486_));
 sky130_fd_sc_hd__buf_1 _33125_ (.A(_16962_),
    .X(_11487_));
 sky130_fd_sc_hd__o2bb2ai_2 _33126_ (.A1_N(_11483_),
    .A2_N(_11486_),
    .B1(_11487_),
    .B2(_18880_),
    .Y(_11488_));
 sky130_fd_sc_hd__a21oi_2 _33127_ (.A1(_11189_),
    .A2(_10883_),
    .B1(_11187_),
    .Y(_11489_));
 sky130_vsdinv _33128_ (.A(_11489_),
    .Y(_11490_));
 sky130_fd_sc_hd__a21oi_2 _33129_ (.A1(_11485_),
    .A2(_11488_),
    .B1(_11490_),
    .Y(_11491_));
 sky130_fd_sc_hd__nand3b_2 _33130_ (.A_N(_11484_),
    .B(_11488_),
    .C(_11490_),
    .Y(_11492_));
 sky130_vsdinv _33131_ (.A(_11492_),
    .Y(_11493_));
 sky130_fd_sc_hd__and2_2 _33132_ (.A(_05438_),
    .B(_11201_),
    .X(_11494_));
 sky130_fd_sc_hd__o21a_2 _33133_ (.A1(_05549_),
    .A2(_07323_),
    .B1(_16961_),
    .X(_11495_));
 sky130_fd_sc_hd__buf_1 _33134_ (.A(_11495_),
    .X(_11496_));
 sky130_fd_sc_hd__nand3_2 _33135_ (.A(_11203_),
    .B(_18866_),
    .C(_05526_),
    .Y(_11497_));
 sky130_fd_sc_hd__nand2_2 _33136_ (.A(_11496_),
    .B(_11497_),
    .Y(_11498_));
 sky130_fd_sc_hd__xnor2_2 _33137_ (.A(_11494_),
    .B(_11498_),
    .Y(_11499_));
 sky130_fd_sc_hd__o21bai_2 _33138_ (.A1(_11491_),
    .A2(_11493_),
    .B1_N(_11499_),
    .Y(_11500_));
 sky130_fd_sc_hd__nand3b_2 _33139_ (.A_N(_11491_),
    .B(_11499_),
    .C(_11492_),
    .Y(_11501_));
 sky130_fd_sc_hd__o21ai_2 _33140_ (.A1(_11207_),
    .A2(_11195_),
    .B1(_11196_),
    .Y(_11502_));
 sky130_fd_sc_hd__a21o_2 _33141_ (.A1(_11500_),
    .A2(_11501_),
    .B1(_11502_),
    .X(_11503_));
 sky130_vsdinv _33142_ (.A(_11200_),
    .Y(_11504_));
 sky130_fd_sc_hd__nor2_2 _33143_ (.A(_11202_),
    .B(_11205_),
    .Y(_11505_));
 sky130_fd_sc_hd__o21ba_2 _33144_ (.A1(_11504_),
    .A2(_11206_),
    .B1_N(_11505_),
    .X(_11506_));
 sky130_vsdinv _33145_ (.A(_11506_),
    .Y(_11507_));
 sky130_fd_sc_hd__nand3_2 _33146_ (.A(_11500_),
    .B(_11501_),
    .C(_11502_),
    .Y(_11508_));
 sky130_fd_sc_hd__nand3_2 _33147_ (.A(_11503_),
    .B(_11507_),
    .C(_11508_),
    .Y(_11509_));
 sky130_fd_sc_hd__a21o_2 _33148_ (.A1(_11503_),
    .A2(_11508_),
    .B1(_11507_),
    .X(_11510_));
 sky130_fd_sc_hd__a22o_2 _33149_ (.A1(_18829_),
    .A2(_11221_),
    .B1(_05873_),
    .B2(_10875_),
    .X(_11511_));
 sky130_fd_sc_hd__nand2_2 _33150_ (.A(_07556_),
    .B(_19156_),
    .Y(_11512_));
 sky130_fd_sc_hd__nand3b_2 _33151_ (.A_N(_11512_),
    .B(_06225_),
    .C(_19162_),
    .Y(_11513_));
 sky130_fd_sc_hd__o2bb2ai_2 _33152_ (.A1_N(_11511_),
    .A2_N(_11513_),
    .B1(_18840_),
    .B2(_19151_),
    .Y(_11514_));
 sky130_fd_sc_hd__buf_1 _33153_ (.A(_09804_),
    .X(_11515_));
 sky130_fd_sc_hd__and2_2 _33154_ (.A(_06101_),
    .B(_11515_),
    .X(_11516_));
 sky130_fd_sc_hd__nand3_2 _33155_ (.A(_11513_),
    .B(_11511_),
    .C(_11516_),
    .Y(_11517_));
 sky130_fd_sc_hd__nand2_2 _33156_ (.A(_11147_),
    .B(_11148_),
    .Y(_11518_));
 sky130_fd_sc_hd__nor2_2 _33157_ (.A(_11147_),
    .B(_11148_),
    .Y(_11519_));
 sky130_fd_sc_hd__a21oi_2 _33158_ (.A1(_11518_),
    .A2(_11146_),
    .B1(_11519_),
    .Y(_11520_));
 sky130_vsdinv _33159_ (.A(_11520_),
    .Y(_11521_));
 sky130_fd_sc_hd__a21o_2 _33160_ (.A1(_11514_),
    .A2(_11517_),
    .B1(_11521_),
    .X(_11522_));
 sky130_fd_sc_hd__nand3_2 _33161_ (.A(_11514_),
    .B(_11521_),
    .C(_11517_),
    .Y(_11523_));
 sky130_fd_sc_hd__a21boi_2 _33162_ (.A1(_11222_),
    .A2(_11227_),
    .B1_N(_11225_),
    .Y(_11524_));
 sky130_vsdinv _33163_ (.A(_11524_),
    .Y(_11525_));
 sky130_fd_sc_hd__a21oi_2 _33164_ (.A1(_11522_),
    .A2(_11523_),
    .B1(_11525_),
    .Y(_11526_));
 sky130_fd_sc_hd__nand3_2 _33165_ (.A(_11522_),
    .B(_11525_),
    .C(_11523_),
    .Y(_11527_));
 sky130_vsdinv _33166_ (.A(_11527_),
    .Y(_11528_));
 sky130_fd_sc_hd__o21ai_2 _33167_ (.A1(_11142_),
    .A2(_11150_),
    .B1(_11143_),
    .Y(_11529_));
 sky130_fd_sc_hd__o21bai_2 _33168_ (.A1(_11526_),
    .A2(_11528_),
    .B1_N(_11529_),
    .Y(_11530_));
 sky130_fd_sc_hd__nand3b_2 _33169_ (.A_N(_11526_),
    .B(_11529_),
    .C(_11527_),
    .Y(_11531_));
 sky130_fd_sc_hd__buf_1 _33170_ (.A(_11531_),
    .X(_11532_));
 sky130_fd_sc_hd__and2_2 _33171_ (.A(_11237_),
    .B(_11234_),
    .X(_11533_));
 sky130_vsdinv _33172_ (.A(_11533_),
    .Y(_11534_));
 sky130_fd_sc_hd__a21oi_2 _33173_ (.A1(_11530_),
    .A2(_11532_),
    .B1(_11534_),
    .Y(_11535_));
 sky130_fd_sc_hd__nand2_2 _33174_ (.A(_11530_),
    .B(_11532_),
    .Y(_11536_));
 sky130_fd_sc_hd__nor2_2 _33175_ (.A(_11533_),
    .B(_11536_),
    .Y(_11537_));
 sky130_fd_sc_hd__o21ai_2 _33176_ (.A1(_11243_),
    .A2(_11239_),
    .B1(_11240_),
    .Y(_11538_));
 sky130_fd_sc_hd__o21bai_2 _33177_ (.A1(_11535_),
    .A2(_11537_),
    .B1_N(_11538_),
    .Y(_11539_));
 sky130_fd_sc_hd__nand2_2 _33178_ (.A(_11536_),
    .B(_11533_),
    .Y(_11540_));
 sky130_fd_sc_hd__nand3b_2 _33179_ (.A_N(_11533_),
    .B(_11530_),
    .C(_11531_),
    .Y(_11541_));
 sky130_fd_sc_hd__nand3_2 _33180_ (.A(_11540_),
    .B(_11538_),
    .C(_11541_),
    .Y(_11542_));
 sky130_fd_sc_hd__a22oi_2 _33181_ (.A1(_11509_),
    .A2(_11510_),
    .B1(_11539_),
    .B2(_11542_),
    .Y(_11543_));
 sky130_fd_sc_hd__nand2_2 _33182_ (.A(_11510_),
    .B(_11509_),
    .Y(_11544_));
 sky130_fd_sc_hd__nand2_2 _33183_ (.A(_11539_),
    .B(_11542_),
    .Y(_11545_));
 sky130_fd_sc_hd__nor2_2 _33184_ (.A(_11544_),
    .B(_11545_),
    .Y(_11546_));
 sky130_fd_sc_hd__o21ai_2 _33185_ (.A1(_11167_),
    .A2(_11169_),
    .B1(_11164_),
    .Y(_11547_));
 sky130_fd_sc_hd__o21bai_2 _33186_ (.A1(_11543_),
    .A2(_11546_),
    .B1_N(_11547_),
    .Y(_11548_));
 sky130_fd_sc_hd__nand2_2 _33187_ (.A(_11545_),
    .B(_11544_),
    .Y(_11549_));
 sky130_fd_sc_hd__a21oi_2 _33188_ (.A1(_11503_),
    .A2(_11508_),
    .B1(_11507_),
    .Y(_11550_));
 sky130_vsdinv _33189_ (.A(_11509_),
    .Y(_11551_));
 sky130_fd_sc_hd__nor2_2 _33190_ (.A(_11550_),
    .B(_11551_),
    .Y(_11552_));
 sky130_fd_sc_hd__nand3_2 _33191_ (.A(_11552_),
    .B(_11542_),
    .C(_11539_),
    .Y(_11553_));
 sky130_fd_sc_hd__nand3_2 _33192_ (.A(_11549_),
    .B(_11547_),
    .C(_11553_),
    .Y(_11554_));
 sky130_fd_sc_hd__buf_1 _33193_ (.A(_11554_),
    .X(_11555_));
 sky130_fd_sc_hd__a21oi_2 _33194_ (.A1(_11252_),
    .A2(_11253_),
    .B1(_11250_),
    .Y(_11556_));
 sky130_fd_sc_hd__a21boi_2 _33195_ (.A1(_11548_),
    .A2(_11555_),
    .B1_N(_11556_),
    .Y(_11557_));
 sky130_fd_sc_hd__buf_1 _33196_ (.A(_11556_),
    .X(_11558_));
 sky130_fd_sc_hd__a21oi_2 _33197_ (.A1(_11549_),
    .A2(_11553_),
    .B1(_11547_),
    .Y(_11559_));
 sky130_fd_sc_hd__nor3b_2 _33198_ (.A(_11558_),
    .B(_11559_),
    .C_N(_11554_),
    .Y(_11560_));
 sky130_fd_sc_hd__nor2_2 _33199_ (.A(_11557_),
    .B(_11560_),
    .Y(_11561_));
 sky130_fd_sc_hd__a21oi_2 _33200_ (.A1(_11475_),
    .A2(_11479_),
    .B1(_11561_),
    .Y(_11562_));
 sky130_fd_sc_hd__nand3_2 _33201_ (.A(_11475_),
    .B(_11561_),
    .C(_11479_),
    .Y(_11563_));
 sky130_vsdinv _33202_ (.A(_11563_),
    .Y(_11564_));
 sky130_fd_sc_hd__o21ai_2 _33203_ (.A1(_11265_),
    .A2(_11267_),
    .B1(_11184_),
    .Y(_11565_));
 sky130_fd_sc_hd__o21bai_2 _33204_ (.A1(_11562_),
    .A2(_11564_),
    .B1_N(_11565_),
    .Y(_11566_));
 sky130_fd_sc_hd__nand2_2 _33205_ (.A(_11475_),
    .B(_11478_),
    .Y(_11567_));
 sky130_fd_sc_hd__a21bo_2 _33206_ (.A1(_11548_),
    .A2(_11555_),
    .B1_N(_11558_),
    .X(_11568_));
 sky130_fd_sc_hd__nand3b_2 _33207_ (.A_N(_11558_),
    .B(_11548_),
    .C(_11555_),
    .Y(_11569_));
 sky130_fd_sc_hd__nand2_2 _33208_ (.A(_11568_),
    .B(_11569_),
    .Y(_11570_));
 sky130_fd_sc_hd__nand2_2 _33209_ (.A(_11567_),
    .B(_11570_),
    .Y(_11571_));
 sky130_fd_sc_hd__nand3_2 _33210_ (.A(_11571_),
    .B(_11565_),
    .C(_11563_),
    .Y(_11572_));
 sky130_fd_sc_hd__buf_1 _33211_ (.A(_11572_),
    .X(_11573_));
 sky130_fd_sc_hd__nand2_2 _33212_ (.A(_11218_),
    .B(_11213_),
    .Y(_11574_));
 sky130_fd_sc_hd__nand2_2 _33213_ (.A(_11263_),
    .B(_11259_),
    .Y(_11575_));
 sky130_fd_sc_hd__xor2_2 _33214_ (.A(_11574_),
    .B(_11575_),
    .X(_11576_));
 sky130_fd_sc_hd__a21o_2 _33215_ (.A1(_11566_),
    .A2(_11573_),
    .B1(_11576_),
    .X(_11577_));
 sky130_fd_sc_hd__nand3_2 _33216_ (.A(_11566_),
    .B(_11576_),
    .C(_11573_),
    .Y(_11578_));
 sky130_fd_sc_hd__a21oi_2 _33217_ (.A1(_11272_),
    .A2(_11273_),
    .B1(_11269_),
    .Y(_11579_));
 sky130_fd_sc_hd__o21ai_2 _33218_ (.A1(_11279_),
    .A2(_11579_),
    .B1(_11274_),
    .Y(_11580_));
 sky130_fd_sc_hd__nand3_2 _33219_ (.A(_11577_),
    .B(_11578_),
    .C(_11580_),
    .Y(_11581_));
 sky130_fd_sc_hd__a21oi_2 _33220_ (.A1(_11566_),
    .A2(_11573_),
    .B1(_11576_),
    .Y(_11582_));
 sky130_vsdinv _33221_ (.A(_11576_),
    .Y(_11583_));
 sky130_fd_sc_hd__a21oi_2 _33222_ (.A1(_11571_),
    .A2(_11563_),
    .B1(_11565_),
    .Y(_11584_));
 sky130_fd_sc_hd__nor3b_2 _33223_ (.A(_11583_),
    .B(_11584_),
    .C_N(_11572_),
    .Y(_11585_));
 sky130_fd_sc_hd__o21bai_2 _33224_ (.A1(_11582_),
    .A2(_11585_),
    .B1_N(_11580_),
    .Y(_11586_));
 sky130_fd_sc_hd__o2bb2ai_2 _33225_ (.A1_N(_11581_),
    .A2_N(_11586_),
    .B1(_11277_),
    .B2(_11276_),
    .Y(_11587_));
 sky130_fd_sc_hd__a21oi_2 _33226_ (.A1(_10940_),
    .A2(_10931_),
    .B1(_11276_),
    .Y(_11588_));
 sky130_fd_sc_hd__nand3_2 _33227_ (.A(_11586_),
    .B(_11588_),
    .C(_11581_),
    .Y(_11589_));
 sky130_fd_sc_hd__o21ai_2 _33228_ (.A1(_11292_),
    .A2(_11284_),
    .B1(_11296_),
    .Y(_11590_));
 sky130_fd_sc_hd__a21oi_2 _33229_ (.A1(_11587_),
    .A2(_11589_),
    .B1(_11590_),
    .Y(_11591_));
 sky130_fd_sc_hd__nand3_2 _33230_ (.A(_11587_),
    .B(_11589_),
    .C(_11590_),
    .Y(_11592_));
 sky130_vsdinv _33231_ (.A(_11592_),
    .Y(_11593_));
 sky130_fd_sc_hd__nor2_2 _33232_ (.A(_11591_),
    .B(_11593_),
    .Y(_11594_));
 sky130_fd_sc_hd__nor2_2 _33233_ (.A(_11303_),
    .B(_10971_),
    .Y(_11595_));
 sky130_fd_sc_hd__a21oi_2 _33234_ (.A1(_11294_),
    .A2(_11297_),
    .B1(_11300_),
    .Y(_11596_));
 sky130_fd_sc_hd__a21oi_2 _33235_ (.A1(_10970_),
    .A2(_11302_),
    .B1(_11596_),
    .Y(_11597_));
 sky130_fd_sc_hd__a21oi_2 _33236_ (.A1(_10993_),
    .A2(_11595_),
    .B1(_11597_),
    .Y(_11598_));
 sky130_fd_sc_hd__xnor2_2 _33237_ (.A(_11594_),
    .B(_11598_),
    .Y(_02653_));
 sky130_fd_sc_hd__buf_1 _33238_ (.A(_10671_),
    .X(_11599_));
 sky130_fd_sc_hd__a22oi_2 _33239_ (.A1(_10481_),
    .A2(_05555_),
    .B1(_19288_),
    .B2(_11599_),
    .Y(_11600_));
 sky130_fd_sc_hd__nand2_2 _33240_ (.A(_18694_),
    .B(_05469_),
    .Y(_11601_));
 sky130_fd_sc_hd__nor3_2 _33241_ (.A(_05987_),
    .B(_11331_),
    .C(_11601_),
    .Y(_11602_));
 sky130_fd_sc_hd__and2_2 _33242_ (.A(_18703_),
    .B(_05528_),
    .X(_11603_));
 sky130_fd_sc_hd__o21bai_2 _33243_ (.A1(_11600_),
    .A2(_11602_),
    .B1_N(_11603_),
    .Y(_11604_));
 sky130_fd_sc_hd__nand3b_2 _33244_ (.A_N(_11601_),
    .B(_10997_),
    .C(_19289_),
    .Y(_11605_));
 sky130_fd_sc_hd__o21ai_2 _33245_ (.A1(_06827_),
    .A2(_16969_),
    .B1(_11601_),
    .Y(_11606_));
 sky130_fd_sc_hd__nand3_2 _33246_ (.A(_11605_),
    .B(_11603_),
    .C(_11606_),
    .Y(_11607_));
 sky130_fd_sc_hd__nor3_2 _33247_ (.A(_05874_),
    .B(_10675_),
    .C(_11321_),
    .Y(_11608_));
 sky130_fd_sc_hd__a21o_2 _33248_ (.A1(_11325_),
    .A2(_11327_),
    .B1(_11608_),
    .X(_11609_));
 sky130_fd_sc_hd__a21o_2 _33249_ (.A1(_11604_),
    .A2(_11607_),
    .B1(_11609_),
    .X(_11610_));
 sky130_fd_sc_hd__nand3_2 _33250_ (.A(_11609_),
    .B(_11604_),
    .C(_11607_),
    .Y(_11611_));
 sky130_fd_sc_hd__buf_1 _33251_ (.A(\pcpi_mul.rs2[28] ),
    .X(_11612_));
 sky130_fd_sc_hd__a22oi_2 _33252_ (.A1(_11014_),
    .A2(_07365_),
    .B1(_11612_),
    .B2(_05837_),
    .Y(_11613_));
 sky130_fd_sc_hd__and4_2 _33253_ (.A(_11011_),
    .B(_11015_),
    .C(_05649_),
    .D(_05739_),
    .X(_11614_));
 sky130_fd_sc_hd__and2_2 _33254_ (.A(_09319_),
    .B(_06074_),
    .X(_11615_));
 sky130_fd_sc_hd__o21bai_2 _33255_ (.A1(_11613_),
    .A2(_11614_),
    .B1_N(_11615_),
    .Y(_11616_));
 sky130_fd_sc_hd__nand2_2 _33256_ (.A(_11612_),
    .B(_07208_),
    .Y(_11617_));
 sky130_fd_sc_hd__buf_1 _33257_ (.A(_18710_),
    .X(_11618_));
 sky130_fd_sc_hd__nand3b_2 _33258_ (.A_N(_11617_),
    .B(_11618_),
    .C(_05931_),
    .Y(_11619_));
 sky130_fd_sc_hd__nand3b_2 _33259_ (.A_N(_11613_),
    .B(_11619_),
    .C(_11615_),
    .Y(_11620_));
 sky130_fd_sc_hd__nand2_2 _33260_ (.A(_11616_),
    .B(_11620_),
    .Y(_11621_));
 sky130_vsdinv _33261_ (.A(_11621_),
    .Y(_11622_));
 sky130_fd_sc_hd__a21oi_2 _33262_ (.A1(_11610_),
    .A2(_11611_),
    .B1(_11622_),
    .Y(_11623_));
 sky130_fd_sc_hd__nand3_2 _33263_ (.A(_11610_),
    .B(_11622_),
    .C(_11611_),
    .Y(_11624_));
 sky130_vsdinv _33264_ (.A(_11624_),
    .Y(_11625_));
 sky130_fd_sc_hd__a21oi_2 _33265_ (.A1(_11336_),
    .A2(_11329_),
    .B1(_11334_),
    .Y(_11626_));
 sky130_fd_sc_hd__o21ai_2 _33266_ (.A1(_11347_),
    .A2(_11626_),
    .B1(_11337_),
    .Y(_11627_));
 sky130_fd_sc_hd__o21bai_2 _33267_ (.A1(_11623_),
    .A2(_11625_),
    .B1_N(_11627_),
    .Y(_11628_));
 sky130_fd_sc_hd__a21oi_2 _33268_ (.A1(_11604_),
    .A2(_11607_),
    .B1(_11609_),
    .Y(_11629_));
 sky130_vsdinv _33269_ (.A(_11611_),
    .Y(_11630_));
 sky130_fd_sc_hd__o21bai_2 _33270_ (.A1(_11629_),
    .A2(_11630_),
    .B1_N(_11622_),
    .Y(_11631_));
 sky130_fd_sc_hd__nand3_2 _33271_ (.A(_11631_),
    .B(_11627_),
    .C(_11624_),
    .Y(_11632_));
 sky130_fd_sc_hd__a22o_2 _33272_ (.A1(_18728_),
    .A2(_05822_),
    .B1(_10453_),
    .B2(_06199_),
    .X(_11633_));
 sky130_fd_sc_hd__buf_1 _33273_ (.A(_09005_),
    .X(_11634_));
 sky130_fd_sc_hd__nand2_2 _33274_ (.A(_11634_),
    .B(_05958_),
    .Y(_11635_));
 sky130_fd_sc_hd__buf_1 _33275_ (.A(_09305_),
    .X(_11636_));
 sky130_fd_sc_hd__nand3b_2 _33276_ (.A_N(_11635_),
    .B(_11636_),
    .C(_06069_),
    .Y(_11637_));
 sky130_fd_sc_hd__o2bb2ai_2 _33277_ (.A1_N(_11633_),
    .A2_N(_11637_),
    .B1(_09011_),
    .B2(_19249_),
    .Y(_11638_));
 sky130_fd_sc_hd__and2_2 _33278_ (.A(_08457_),
    .B(_06360_),
    .X(_11639_));
 sky130_fd_sc_hd__nand3_2 _33279_ (.A(_11637_),
    .B(_11633_),
    .C(_11639_),
    .Y(_11640_));
 sky130_fd_sc_hd__o31ai_2 _33280_ (.A1(_18725_),
    .A2(_19268_),
    .A3(_11339_),
    .B1(_11345_),
    .Y(_11641_));
 sky130_fd_sc_hd__a21o_2 _33281_ (.A1(_11638_),
    .A2(_11640_),
    .B1(_11641_),
    .X(_11642_));
 sky130_fd_sc_hd__nand3_2 _33282_ (.A(_11641_),
    .B(_11638_),
    .C(_11640_),
    .Y(_11643_));
 sky130_fd_sc_hd__buf_1 _33283_ (.A(_11643_),
    .X(_11644_));
 sky130_fd_sc_hd__nand3b_2 _33284_ (.A_N(_11305_),
    .B(_11042_),
    .C(_06344_),
    .Y(_11645_));
 sky130_fd_sc_hd__a21boi_2 _33285_ (.A1(_11307_),
    .A2(_11308_),
    .B1_N(_11645_),
    .Y(_11646_));
 sky130_vsdinv _33286_ (.A(_11646_),
    .Y(_11647_));
 sky130_fd_sc_hd__a21oi_2 _33287_ (.A1(_11642_),
    .A2(_11644_),
    .B1(_11647_),
    .Y(_11648_));
 sky130_fd_sc_hd__a21oi_2 _33288_ (.A1(_11638_),
    .A2(_11640_),
    .B1(_11641_),
    .Y(_11649_));
 sky130_fd_sc_hd__nor3b_2 _33289_ (.A(_11646_),
    .B(_11649_),
    .C_N(_11643_),
    .Y(_11650_));
 sky130_fd_sc_hd__nor2_2 _33290_ (.A(_11648_),
    .B(_11650_),
    .Y(_11651_));
 sky130_fd_sc_hd__a21oi_2 _33291_ (.A1(_11628_),
    .A2(_11632_),
    .B1(_11651_),
    .Y(_11652_));
 sky130_fd_sc_hd__nand3_2 _33292_ (.A(_11628_),
    .B(_11651_),
    .C(_11632_),
    .Y(_11653_));
 sky130_vsdinv _33293_ (.A(_11653_),
    .Y(_11654_));
 sky130_fd_sc_hd__a21oi_2 _33294_ (.A1(_11355_),
    .A2(_11350_),
    .B1(_11353_),
    .Y(_11655_));
 sky130_fd_sc_hd__o21ai_2 _33295_ (.A1(_11358_),
    .A2(_11655_),
    .B1(_11356_),
    .Y(_11656_));
 sky130_fd_sc_hd__o21bai_2 _33296_ (.A1(_11652_),
    .A2(_11654_),
    .B1_N(_11656_),
    .Y(_11657_));
 sky130_fd_sc_hd__a21oi_2 _33297_ (.A1(_11631_),
    .A2(_11624_),
    .B1(_11627_),
    .Y(_11658_));
 sky130_vsdinv _33298_ (.A(_11632_),
    .Y(_11659_));
 sky130_fd_sc_hd__o21bai_2 _33299_ (.A1(_11658_),
    .A2(_11659_),
    .B1_N(_11651_),
    .Y(_11660_));
 sky130_fd_sc_hd__nand3_2 _33300_ (.A(_11660_),
    .B(_11656_),
    .C(_11653_),
    .Y(_11661_));
 sky130_fd_sc_hd__buf_1 _33301_ (.A(_11661_),
    .X(_11662_));
 sky130_fd_sc_hd__nand2_2 _33302_ (.A(_08471_),
    .B(_06364_),
    .Y(_11663_));
 sky130_fd_sc_hd__nand2_2 _33303_ (.A(_08971_),
    .B(_07099_),
    .Y(_11664_));
 sky130_fd_sc_hd__xnor2_2 _33304_ (.A(_11663_),
    .B(_11664_),
    .Y(_11665_));
 sky130_fd_sc_hd__o21ai_2 _33305_ (.A1(_18759_),
    .A2(_19233_),
    .B1(_11665_),
    .Y(_11666_));
 sky130_fd_sc_hd__nor2_2 _33306_ (.A(_11663_),
    .B(_11664_),
    .Y(_11667_));
 sky130_fd_sc_hd__and2_2 _33307_ (.A(_08235_),
    .B(_08186_),
    .X(_11668_));
 sky130_fd_sc_hd__nand2_2 _33308_ (.A(_11663_),
    .B(_11664_),
    .Y(_11669_));
 sky130_fd_sc_hd__nand3b_2 _33309_ (.A_N(_11667_),
    .B(_11668_),
    .C(_11669_),
    .Y(_11670_));
 sky130_fd_sc_hd__nand2_2 _33310_ (.A(_11666_),
    .B(_11670_),
    .Y(_11671_));
 sky130_fd_sc_hd__nor2_2 _33311_ (.A(_11366_),
    .B(_11367_),
    .Y(_11672_));
 sky130_fd_sc_hd__a21oi_2 _33312_ (.A1(_11368_),
    .A2(_11371_),
    .B1(_11672_),
    .Y(_11673_));
 sky130_fd_sc_hd__nand2_2 _33313_ (.A(_11671_),
    .B(_11673_),
    .Y(_11674_));
 sky130_fd_sc_hd__nand3b_2 _33314_ (.A_N(_11673_),
    .B(_11666_),
    .C(_11670_),
    .Y(_11675_));
 sky130_fd_sc_hd__nand2_2 _33315_ (.A(_11674_),
    .B(_11675_),
    .Y(_11676_));
 sky130_fd_sc_hd__and2_2 _33316_ (.A(_07421_),
    .B(_06937_),
    .X(_11677_));
 sky130_fd_sc_hd__and4_2 _33317_ (.A(_07850_),
    .B(_08214_),
    .C(_19215_),
    .D(_08261_),
    .X(_11678_));
 sky130_vsdinv _33318_ (.A(_11678_),
    .Y(_11679_));
 sky130_fd_sc_hd__a22oi_2 _33319_ (.A1(_07537_),
    .A2(_19225_),
    .B1(_07535_),
    .B2(_07328_),
    .Y(_11680_));
 sky130_vsdinv _33320_ (.A(_11680_),
    .Y(_11681_));
 sky130_fd_sc_hd__nand2_2 _33321_ (.A(_11679_),
    .B(_11681_),
    .Y(_11682_));
 sky130_fd_sc_hd__xor2_2 _33322_ (.A(_11677_),
    .B(_11682_),
    .X(_11683_));
 sky130_fd_sc_hd__nand2_2 _33323_ (.A(_11676_),
    .B(_11683_),
    .Y(_11684_));
 sky130_fd_sc_hd__xnor2_2 _33324_ (.A(_11677_),
    .B(_11682_),
    .Y(_11685_));
 sky130_fd_sc_hd__nand3_2 _33325_ (.A(_11685_),
    .B(_11674_),
    .C(_11675_),
    .Y(_11686_));
 sky130_fd_sc_hd__nand2_2 _33326_ (.A(_11684_),
    .B(_11686_),
    .Y(_11687_));
 sky130_fd_sc_hd__nand3_2 _33327_ (.A(_11687_),
    .B(_11318_),
    .C(_11319_),
    .Y(_11688_));
 sky130_fd_sc_hd__nand2_2 _33328_ (.A(_11319_),
    .B(_11318_),
    .Y(_11689_));
 sky130_fd_sc_hd__nand3_2 _33329_ (.A(_11689_),
    .B(_11684_),
    .C(_11686_),
    .Y(_11690_));
 sky130_fd_sc_hd__nand2_2 _33330_ (.A(_11688_),
    .B(_11690_),
    .Y(_11691_));
 sky130_vsdinv _33331_ (.A(_11377_),
    .Y(_11692_));
 sky130_fd_sc_hd__a21oi_2 _33332_ (.A1(_11382_),
    .A2(_11376_),
    .B1(_11692_),
    .Y(_11693_));
 sky130_fd_sc_hd__nand2_2 _33333_ (.A(_11691_),
    .B(_11693_),
    .Y(_11694_));
 sky130_vsdinv _33334_ (.A(_11693_),
    .Y(_11695_));
 sky130_fd_sc_hd__nand3_2 _33335_ (.A(_11688_),
    .B(_11695_),
    .C(_11690_),
    .Y(_11696_));
 sky130_fd_sc_hd__nand2_2 _33336_ (.A(_11694_),
    .B(_11696_),
    .Y(_11697_));
 sky130_fd_sc_hd__buf_1 _33337_ (.A(_11697_),
    .X(_11698_));
 sky130_fd_sc_hd__a21boi_2 _33338_ (.A1(_11657_),
    .A2(_11662_),
    .B1_N(_11698_),
    .Y(_11699_));
 sky130_fd_sc_hd__a21oi_2 _33339_ (.A1(_11660_),
    .A2(_11653_),
    .B1(_11656_),
    .Y(_11700_));
 sky130_fd_sc_hd__nor3b_2 _33340_ (.A(_11698_),
    .B(_11700_),
    .C_N(_11662_),
    .Y(_11701_));
 sky130_fd_sc_hd__a21o_2 _33341_ (.A1(_11387_),
    .A2(_11390_),
    .B1(_11392_),
    .X(_11702_));
 sky130_fd_sc_hd__nand3_2 _33342_ (.A(_11392_),
    .B(_11387_),
    .C(_11390_),
    .Y(_11703_));
 sky130_fd_sc_hd__nand2_2 _33343_ (.A(_11702_),
    .B(_11703_),
    .Y(_11704_));
 sky130_fd_sc_hd__o21ai_2 _33344_ (.A1(_11704_),
    .A2(_11402_),
    .B1(_11365_),
    .Y(_11705_));
 sky130_fd_sc_hd__o21bai_2 _33345_ (.A1(_11699_),
    .A2(_11701_),
    .B1_N(_11705_),
    .Y(_11706_));
 sky130_fd_sc_hd__nand2_2 _33346_ (.A(_11657_),
    .B(_11661_),
    .Y(_11707_));
 sky130_fd_sc_hd__nand2_2 _33347_ (.A(_11707_),
    .B(_11698_),
    .Y(_11708_));
 sky130_fd_sc_hd__nand3b_2 _33348_ (.A_N(_11697_),
    .B(_11657_),
    .C(_11662_),
    .Y(_11709_));
 sky130_fd_sc_hd__nand3_2 _33349_ (.A(_11708_),
    .B(_11705_),
    .C(_11709_),
    .Y(_11710_));
 sky130_fd_sc_hd__buf_1 _33350_ (.A(_11710_),
    .X(_11711_));
 sky130_fd_sc_hd__a22o_2 _33351_ (.A1(_11108_),
    .A2(_07942_),
    .B1(_08142_),
    .B2(_08303_),
    .X(_11712_));
 sky130_fd_sc_hd__nand2_2 _33352_ (.A(_10120_),
    .B(_09364_),
    .Y(_11713_));
 sky130_fd_sc_hd__buf_1 _33353_ (.A(_08551_),
    .X(_11714_));
 sky130_fd_sc_hd__nand3b_2 _33354_ (.A_N(_11713_),
    .B(_18786_),
    .C(_11714_),
    .Y(_11715_));
 sky130_fd_sc_hd__buf_1 _33355_ (.A(_18792_),
    .X(_11716_));
 sky130_fd_sc_hd__o2bb2ai_2 _33356_ (.A1_N(_11712_),
    .A2_N(_11715_),
    .B1(_11716_),
    .B2(_19198_),
    .Y(_11717_));
 sky130_fd_sc_hd__and2_2 _33357_ (.A(_07402_),
    .B(_10162_),
    .X(_11718_));
 sky130_fd_sc_hd__nand3_2 _33358_ (.A(_11715_),
    .B(_11712_),
    .C(_11718_),
    .Y(_11719_));
 sky130_fd_sc_hd__nand2_2 _33359_ (.A(_11379_),
    .B(_11380_),
    .Y(_11720_));
 sky130_fd_sc_hd__nor2_2 _33360_ (.A(_11379_),
    .B(_11380_),
    .Y(_11721_));
 sky130_fd_sc_hd__a21oi_2 _33361_ (.A1(_11720_),
    .A2(_11378_),
    .B1(_11721_),
    .Y(_11722_));
 sky130_vsdinv _33362_ (.A(_11722_),
    .Y(_11723_));
 sky130_fd_sc_hd__a21oi_2 _33363_ (.A1(_11717_),
    .A2(_11719_),
    .B1(_11723_),
    .Y(_11724_));
 sky130_fd_sc_hd__nand3_2 _33364_ (.A(_11717_),
    .B(_11723_),
    .C(_11719_),
    .Y(_11725_));
 sky130_vsdinv _33365_ (.A(_11725_),
    .Y(_11726_));
 sky130_fd_sc_hd__nand3b_2 _33366_ (.A_N(_11406_),
    .B(_18787_),
    .C(_08301_),
    .Y(_11727_));
 sky130_fd_sc_hd__a21boi_2 _33367_ (.A1(_11408_),
    .A2(_11410_),
    .B1_N(_11727_),
    .Y(_11728_));
 sky130_fd_sc_hd__o21ai_2 _33368_ (.A1(_11724_),
    .A2(_11726_),
    .B1(_11728_),
    .Y(_11729_));
 sky130_vsdinv _33369_ (.A(_11728_),
    .Y(_11730_));
 sky130_fd_sc_hd__nand3b_2 _33370_ (.A_N(_11724_),
    .B(_11730_),
    .C(_11725_),
    .Y(_11731_));
 sky130_fd_sc_hd__o21ai_2 _33371_ (.A1(_11421_),
    .A2(_11418_),
    .B1(_11419_),
    .Y(_11732_));
 sky130_fd_sc_hd__a21o_2 _33372_ (.A1(_11729_),
    .A2(_11731_),
    .B1(_11732_),
    .X(_11733_));
 sky130_fd_sc_hd__nand3_2 _33373_ (.A(_11732_),
    .B(_11729_),
    .C(_11731_),
    .Y(_11734_));
 sky130_fd_sc_hd__and2_2 _33374_ (.A(_06138_),
    .B(_10538_),
    .X(_11735_));
 sky130_fd_sc_hd__buf_1 _33375_ (.A(_19166_),
    .X(_11736_));
 sky130_fd_sc_hd__a22oi_2 _33376_ (.A1(_06671_),
    .A2(_08833_),
    .B1(_06142_),
    .B2(_11736_),
    .Y(_11737_));
 sky130_fd_sc_hd__and4_2 _33377_ (.A(_06811_),
    .B(_11432_),
    .C(_09786_),
    .D(_11433_),
    .X(_11738_));
 sky130_fd_sc_hd__nor2_2 _33378_ (.A(_11737_),
    .B(_11738_),
    .Y(_11739_));
 sky130_fd_sc_hd__xnor2_2 _33379_ (.A(_11735_),
    .B(_11739_),
    .Y(_11740_));
 sky130_fd_sc_hd__nand2_2 _33380_ (.A(_08414_),
    .B(_09456_),
    .Y(_11741_));
 sky130_fd_sc_hd__nand2_2 _33381_ (.A(_06540_),
    .B(_07951_),
    .Y(_11742_));
 sky130_fd_sc_hd__nand2_2 _33382_ (.A(_11741_),
    .B(_11742_),
    .Y(_11743_));
 sky130_fd_sc_hd__nand3b_2 _33383_ (.A_N(_11741_),
    .B(_06538_),
    .C(_08827_),
    .Y(_11744_));
 sky130_fd_sc_hd__buf_1 _33384_ (.A(_18809_),
    .X(_11745_));
 sky130_fd_sc_hd__o2bb2ai_2 _33385_ (.A1_N(_11743_),
    .A2_N(_11744_),
    .B1(_11745_),
    .B2(_09092_),
    .Y(_11746_));
 sky130_fd_sc_hd__and2_2 _33386_ (.A(_06550_),
    .B(_19180_),
    .X(_11747_));
 sky130_fd_sc_hd__nand3_2 _33387_ (.A(_11744_),
    .B(_11747_),
    .C(_11743_),
    .Y(_11748_));
 sky130_fd_sc_hd__nor2_2 _33388_ (.A(_11438_),
    .B(_11439_),
    .Y(_11749_));
 sky130_fd_sc_hd__a21oi_2 _33389_ (.A1(_11440_),
    .A2(_11444_),
    .B1(_11749_),
    .Y(_11750_));
 sky130_vsdinv _33390_ (.A(_11750_),
    .Y(_11751_));
 sky130_fd_sc_hd__a21oi_2 _33391_ (.A1(_11746_),
    .A2(_11748_),
    .B1(_11751_),
    .Y(_11752_));
 sky130_vsdinv _33392_ (.A(_11752_),
    .Y(_11753_));
 sky130_fd_sc_hd__nand3_2 _33393_ (.A(_11746_),
    .B(_11751_),
    .C(_11748_),
    .Y(_11754_));
 sky130_fd_sc_hd__nand3b_2 _33394_ (.A_N(_11740_),
    .B(_11753_),
    .C(_11754_),
    .Y(_11755_));
 sky130_vsdinv _33395_ (.A(_11754_),
    .Y(_11756_));
 sky130_fd_sc_hd__o21ai_2 _33396_ (.A1(_11752_),
    .A2(_11756_),
    .B1(_11740_),
    .Y(_11757_));
 sky130_fd_sc_hd__nand2_2 _33397_ (.A(_11755_),
    .B(_11757_),
    .Y(_11758_));
 sky130_vsdinv _33398_ (.A(_11758_),
    .Y(_11759_));
 sky130_fd_sc_hd__a21o_2 _33399_ (.A1(_11733_),
    .A2(_11734_),
    .B1(_11759_),
    .X(_11760_));
 sky130_fd_sc_hd__nand3_2 _33400_ (.A(_11733_),
    .B(_11759_),
    .C(_11734_),
    .Y(_11761_));
 sky130_fd_sc_hd__o21ai_2 _33401_ (.A1(_11391_),
    .A2(_11394_),
    .B1(_11389_),
    .Y(_11762_));
 sky130_fd_sc_hd__a21o_2 _33402_ (.A1(_11760_),
    .A2(_11761_),
    .B1(_11762_),
    .X(_11763_));
 sky130_fd_sc_hd__nand3_2 _33403_ (.A(_11760_),
    .B(_11762_),
    .C(_11761_),
    .Y(_11764_));
 sky130_fd_sc_hd__a21oi_2 _33404_ (.A1(_11454_),
    .A2(_11452_),
    .B1(_11429_),
    .Y(_11765_));
 sky130_vsdinv _33405_ (.A(_11765_),
    .Y(_11766_));
 sky130_fd_sc_hd__a21oi_2 _33406_ (.A1(_11763_),
    .A2(_11764_),
    .B1(_11766_),
    .Y(_11767_));
 sky130_fd_sc_hd__a21oi_2 _33407_ (.A1(_11760_),
    .A2(_11761_),
    .B1(_11762_),
    .Y(_11768_));
 sky130_vsdinv _33408_ (.A(_11764_),
    .Y(_11769_));
 sky130_fd_sc_hd__nor3_2 _33409_ (.A(_11765_),
    .B(_11768_),
    .C(_11769_),
    .Y(_11770_));
 sky130_fd_sc_hd__nor2_2 _33410_ (.A(_11767_),
    .B(_11770_),
    .Y(_11771_));
 sky130_fd_sc_hd__a21oi_2 _33411_ (.A1(_11706_),
    .A2(_11711_),
    .B1(_11771_),
    .Y(_11772_));
 sky130_fd_sc_hd__o21bai_2 _33412_ (.A1(_11768_),
    .A2(_11769_),
    .B1_N(_11766_),
    .Y(_11773_));
 sky130_fd_sc_hd__nand3_2 _33413_ (.A(_11763_),
    .B(_11766_),
    .C(_11764_),
    .Y(_11774_));
 sky130_fd_sc_hd__nand2_2 _33414_ (.A(_11773_),
    .B(_11774_),
    .Y(_11775_));
 sky130_fd_sc_hd__a21oi_2 _33415_ (.A1(_11708_),
    .A2(_11709_),
    .B1(_11705_),
    .Y(_11776_));
 sky130_vsdinv _33416_ (.A(_11711_),
    .Y(_11777_));
 sky130_fd_sc_hd__nor3_2 _33417_ (.A(_11775_),
    .B(_11776_),
    .C(_11777_),
    .Y(_11778_));
 sky130_fd_sc_hd__o21ai_2 _33418_ (.A1(_11470_),
    .A2(_11471_),
    .B1(_11405_),
    .Y(_11779_));
 sky130_fd_sc_hd__o21bai_2 _33419_ (.A1(_11772_),
    .A2(_11778_),
    .B1_N(_11779_),
    .Y(_11780_));
 sky130_fd_sc_hd__nand2_2 _33420_ (.A(_11706_),
    .B(_11710_),
    .Y(_11781_));
 sky130_fd_sc_hd__nand2_2 _33421_ (.A(_11781_),
    .B(_11775_),
    .Y(_11782_));
 sky130_fd_sc_hd__nand3_2 _33422_ (.A(_11771_),
    .B(_11706_),
    .C(_11711_),
    .Y(_11783_));
 sky130_fd_sc_hd__nand3_2 _33423_ (.A(_11782_),
    .B(_11779_),
    .C(_11783_),
    .Y(_11784_));
 sky130_fd_sc_hd__buf_1 _33424_ (.A(_11784_),
    .X(_11785_));
 sky130_fd_sc_hd__a22o_2 _33425_ (.A1(_18829_),
    .A2(_10875_),
    .B1(_06230_),
    .B2(_11515_),
    .X(_11786_));
 sky130_fd_sc_hd__nand2_2 _33426_ (.A(_07697_),
    .B(_09500_),
    .Y(_11787_));
 sky130_fd_sc_hd__buf_1 _33427_ (.A(_10532_),
    .X(_11788_));
 sky130_fd_sc_hd__nand3b_2 _33428_ (.A_N(_11787_),
    .B(_05983_),
    .C(_11788_),
    .Y(_11789_));
 sky130_fd_sc_hd__o2bb2ai_2 _33429_ (.A1_N(_11786_),
    .A2_N(_11789_),
    .B1(_07920_),
    .B2(_19145_),
    .Y(_11790_));
 sky130_fd_sc_hd__buf_1 _33430_ (.A(_10554_),
    .X(_11791_));
 sky130_fd_sc_hd__and2_2 _33431_ (.A(_06101_),
    .B(_11791_),
    .X(_11792_));
 sky130_fd_sc_hd__nand3_2 _33432_ (.A(_11789_),
    .B(_11786_),
    .C(_11792_),
    .Y(_11793_));
 sky130_fd_sc_hd__nand2_2 _33433_ (.A(_11790_),
    .B(_11793_),
    .Y(_11794_));
 sky130_vsdinv _33434_ (.A(_11431_),
    .Y(_11795_));
 sky130_fd_sc_hd__a21oi_2 _33435_ (.A1(_11795_),
    .A2(_11430_),
    .B1(_11435_),
    .Y(_11796_));
 sky130_fd_sc_hd__nand2_2 _33436_ (.A(_11794_),
    .B(_11796_),
    .Y(_11797_));
 sky130_fd_sc_hd__a21o_2 _33437_ (.A1(_11795_),
    .A2(_11430_),
    .B1(_11435_),
    .X(_11798_));
 sky130_fd_sc_hd__nand3_2 _33438_ (.A(_11798_),
    .B(_11790_),
    .C(_11793_),
    .Y(_11799_));
 sky130_fd_sc_hd__a21boi_2 _33439_ (.A1(_11511_),
    .A2(_11516_),
    .B1_N(_11513_),
    .Y(_11800_));
 sky130_vsdinv _33440_ (.A(_11800_),
    .Y(_11801_));
 sky130_fd_sc_hd__a21oi_2 _33441_ (.A1(_11797_),
    .A2(_11799_),
    .B1(_11801_),
    .Y(_11802_));
 sky130_vsdinv _33442_ (.A(_11450_),
    .Y(_11803_));
 sky130_fd_sc_hd__o21bai_2 _33443_ (.A1(_11437_),
    .A2(_11451_),
    .B1_N(_11803_),
    .Y(_11804_));
 sky130_fd_sc_hd__nand3_2 _33444_ (.A(_11797_),
    .B(_11799_),
    .C(_11801_),
    .Y(_11805_));
 sky130_fd_sc_hd__nand3b_2 _33445_ (.A_N(_11802_),
    .B(_11804_),
    .C(_11805_),
    .Y(_11806_));
 sky130_vsdinv _33446_ (.A(_11805_),
    .Y(_11807_));
 sky130_vsdinv _33447_ (.A(_11437_),
    .Y(_11808_));
 sky130_fd_sc_hd__a21oi_2 _33448_ (.A1(_11808_),
    .A2(_11449_),
    .B1(_11803_),
    .Y(_11809_));
 sky130_fd_sc_hd__o21ai_2 _33449_ (.A1(_11802_),
    .A2(_11807_),
    .B1(_11809_),
    .Y(_11810_));
 sky130_fd_sc_hd__a21boi_2 _33450_ (.A1(_11522_),
    .A2(_11525_),
    .B1_N(_11523_),
    .Y(_11811_));
 sky130_vsdinv _33451_ (.A(_11811_),
    .Y(_11812_));
 sky130_fd_sc_hd__a21oi_2 _33452_ (.A1(_11806_),
    .A2(_11810_),
    .B1(_11812_),
    .Y(_11813_));
 sky130_fd_sc_hd__nand3_2 _33453_ (.A(_11806_),
    .B(_11810_),
    .C(_11812_),
    .Y(_11814_));
 sky130_vsdinv _33454_ (.A(_11814_),
    .Y(_11815_));
 sky130_fd_sc_hd__a21boi_2 _33455_ (.A1(_11534_),
    .A2(_11530_),
    .B1_N(_11532_),
    .Y(_11816_));
 sky130_fd_sc_hd__o21ai_2 _33456_ (.A1(_11813_),
    .A2(_11815_),
    .B1(_11816_),
    .Y(_11817_));
 sky130_fd_sc_hd__nand2_2 _33457_ (.A(_11541_),
    .B(_11532_),
    .Y(_11818_));
 sky130_fd_sc_hd__nand3b_2 _33458_ (.A_N(_11813_),
    .B(_11814_),
    .C(_11818_),
    .Y(_11819_));
 sky130_fd_sc_hd__nand2_2 _33459_ (.A(_06040_),
    .B(_10912_),
    .Y(_11820_));
 sky130_fd_sc_hd__nand2_2 _33460_ (.A(_08291_),
    .B(_10899_),
    .Y(_11821_));
 sky130_fd_sc_hd__nand2_2 _33461_ (.A(_11820_),
    .B(_11821_),
    .Y(_11822_));
 sky130_fd_sc_hd__nand3b_2 _33462_ (.A_N(_11820_),
    .B(_05826_),
    .C(_19133_),
    .Y(_11823_));
 sky130_fd_sc_hd__o2bb2ai_2 _33463_ (.A1_N(_11822_),
    .A2_N(_11823_),
    .B1(_16962_),
    .B2(_06346_),
    .Y(_11824_));
 sky130_fd_sc_hd__nand3_2 _33464_ (.A(_11823_),
    .B(_10883_),
    .C(_11822_),
    .Y(_11825_));
 sky130_fd_sc_hd__a21oi_2 _33465_ (.A1(_11483_),
    .A2(_10882_),
    .B1(_11482_),
    .Y(_11826_));
 sky130_vsdinv _33466_ (.A(_11826_),
    .Y(_11827_));
 sky130_fd_sc_hd__a21o_2 _33467_ (.A1(_11824_),
    .A2(_11825_),
    .B1(_11827_),
    .X(_11828_));
 sky130_fd_sc_hd__nand3b_2 _33468_ (.A_N(_11826_),
    .B(_11824_),
    .C(_11825_),
    .Y(_11829_));
 sky130_fd_sc_hd__buf_1 _33469_ (.A(_16960_),
    .X(_11830_));
 sky130_fd_sc_hd__and2_2 _33470_ (.A(_11830_),
    .B(_05437_),
    .X(_11831_));
 sky130_fd_sc_hd__a21oi_2 _33471_ (.A1(_11496_),
    .A2(_11497_),
    .B1(_11831_),
    .Y(_11832_));
 sky130_fd_sc_hd__and3_2 _33472_ (.A(_11495_),
    .B(_11831_),
    .C(_11497_),
    .X(_11833_));
 sky130_fd_sc_hd__nor2_2 _33473_ (.A(_11832_),
    .B(_11833_),
    .Y(_11834_));
 sky130_fd_sc_hd__buf_1 _33474_ (.A(_11834_),
    .X(_11835_));
 sky130_fd_sc_hd__a21oi_2 _33475_ (.A1(_11828_),
    .A2(_11829_),
    .B1(_11835_),
    .Y(_11836_));
 sky130_fd_sc_hd__and3_2 _33476_ (.A(_11828_),
    .B(_11834_),
    .C(_11829_),
    .X(_11837_));
 sky130_vsdinv _33477_ (.A(_11837_),
    .Y(_11838_));
 sky130_vsdinv _33478_ (.A(_11499_),
    .Y(_11839_));
 sky130_fd_sc_hd__o21ai_2 _33479_ (.A1(_11839_),
    .A2(_11491_),
    .B1(_11492_),
    .Y(_11840_));
 sky130_fd_sc_hd__nand3b_2 _33480_ (.A_N(_11836_),
    .B(_11838_),
    .C(_11840_),
    .Y(_11841_));
 sky130_fd_sc_hd__o21bai_2 _33481_ (.A1(_11836_),
    .A2(_11837_),
    .B1_N(_11840_),
    .Y(_11842_));
 sky130_vsdinv _33482_ (.A(_11497_),
    .Y(_11843_));
 sky130_fd_sc_hd__a21oi_2 _33483_ (.A1(_11496_),
    .A2(_11494_),
    .B1(_11843_),
    .Y(_11844_));
 sky130_fd_sc_hd__a21bo_2 _33484_ (.A1(_11841_),
    .A2(_11842_),
    .B1_N(_11844_),
    .X(_11845_));
 sky130_fd_sc_hd__nand3b_2 _33485_ (.A_N(_11844_),
    .B(_11841_),
    .C(_11842_),
    .Y(_11846_));
 sky130_fd_sc_hd__nand2_2 _33486_ (.A(_11845_),
    .B(_11846_),
    .Y(_11847_));
 sky130_fd_sc_hd__buf_1 _33487_ (.A(_11847_),
    .X(_11848_));
 sky130_fd_sc_hd__a21boi_2 _33488_ (.A1(_11817_),
    .A2(_11819_),
    .B1_N(_11848_),
    .Y(_11849_));
 sky130_fd_sc_hd__nand2_2 _33489_ (.A(_11817_),
    .B(_11819_),
    .Y(_11850_));
 sky130_fd_sc_hd__nor2_2 _33490_ (.A(_11848_),
    .B(_11850_),
    .Y(_11851_));
 sky130_fd_sc_hd__o21ai_2 _33491_ (.A1(_11460_),
    .A2(_11467_),
    .B1(_11458_),
    .Y(_11852_));
 sky130_fd_sc_hd__o21bai_2 _33492_ (.A1(_11849_),
    .A2(_11851_),
    .B1_N(_11852_),
    .Y(_11853_));
 sky130_fd_sc_hd__nand2_2 _33493_ (.A(_11850_),
    .B(_11848_),
    .Y(_11854_));
 sky130_fd_sc_hd__nand3b_2 _33494_ (.A_N(_11847_),
    .B(_11819_),
    .C(_11817_),
    .Y(_11855_));
 sky130_fd_sc_hd__nand3_2 _33495_ (.A(_11854_),
    .B(_11855_),
    .C(_11852_),
    .Y(_11856_));
 sky130_fd_sc_hd__nand2_2 _33496_ (.A(_11853_),
    .B(_11856_),
    .Y(_11857_));
 sky130_fd_sc_hd__a21boi_2 _33497_ (.A1(_11552_),
    .A2(_11539_),
    .B1_N(_11542_),
    .Y(_11858_));
 sky130_fd_sc_hd__nand2_2 _33498_ (.A(_11857_),
    .B(_11858_),
    .Y(_11859_));
 sky130_fd_sc_hd__nand3b_2 _33499_ (.A_N(_11858_),
    .B(_11853_),
    .C(_11856_),
    .Y(_11860_));
 sky130_fd_sc_hd__nand2_2 _33500_ (.A(_11859_),
    .B(_11860_),
    .Y(_11861_));
 sky130_fd_sc_hd__buf_1 _33501_ (.A(_11861_),
    .X(_11862_));
 sky130_fd_sc_hd__a21boi_2 _33502_ (.A1(_11780_),
    .A2(_11785_),
    .B1_N(_11862_),
    .Y(_11863_));
 sky130_fd_sc_hd__a21oi_2 _33503_ (.A1(_11782_),
    .A2(_11783_),
    .B1(_11779_),
    .Y(_11864_));
 sky130_fd_sc_hd__nor3b_2 _33504_ (.A(_11862_),
    .B(_11864_),
    .C_N(_11785_),
    .Y(_11865_));
 sky130_fd_sc_hd__a21oi_2 _33505_ (.A1(_11476_),
    .A2(_11477_),
    .B1(_11474_),
    .Y(_11866_));
 sky130_fd_sc_hd__o21ai_2 _33506_ (.A1(_11570_),
    .A2(_11866_),
    .B1(_11479_),
    .Y(_11867_));
 sky130_fd_sc_hd__o21bai_2 _33507_ (.A1(_11863_),
    .A2(_11865_),
    .B1_N(_11867_),
    .Y(_11868_));
 sky130_fd_sc_hd__nand2_2 _33508_ (.A(_11780_),
    .B(_11785_),
    .Y(_11869_));
 sky130_fd_sc_hd__nand2_2 _33509_ (.A(_11869_),
    .B(_11862_),
    .Y(_11870_));
 sky130_fd_sc_hd__nand3b_2 _33510_ (.A_N(_11862_),
    .B(_11780_),
    .C(_11785_),
    .Y(_11871_));
 sky130_fd_sc_hd__nand3_2 _33511_ (.A(_11870_),
    .B(_11867_),
    .C(_11871_),
    .Y(_11872_));
 sky130_vsdinv _33512_ (.A(_11508_),
    .Y(_11873_));
 sky130_fd_sc_hd__a21oi_2 _33513_ (.A1(_11503_),
    .A2(_11507_),
    .B1(_11873_),
    .Y(_11874_));
 sky130_fd_sc_hd__o21ai_2 _33514_ (.A1(_11558_),
    .A2(_11559_),
    .B1(_11555_),
    .Y(_11875_));
 sky130_fd_sc_hd__xnor2_2 _33515_ (.A(_11874_),
    .B(_11875_),
    .Y(_11876_));
 sky130_fd_sc_hd__a21oi_2 _33516_ (.A1(_11868_),
    .A2(_11872_),
    .B1(_11876_),
    .Y(_11877_));
 sky130_vsdinv _33517_ (.A(_11876_),
    .Y(_11878_));
 sky130_fd_sc_hd__a21oi_2 _33518_ (.A1(_11870_),
    .A2(_11871_),
    .B1(_11867_),
    .Y(_11879_));
 sky130_fd_sc_hd__a21boi_2 _33519_ (.A1(_11475_),
    .A2(_11561_),
    .B1_N(_11479_),
    .Y(_11880_));
 sky130_fd_sc_hd__nor3_2 _33520_ (.A(_11863_),
    .B(_11880_),
    .C(_11865_),
    .Y(_11881_));
 sky130_fd_sc_hd__nor3_2 _33521_ (.A(_11878_),
    .B(_11879_),
    .C(_11881_),
    .Y(_11882_));
 sky130_fd_sc_hd__o21ai_2 _33522_ (.A1(_11583_),
    .A2(_11584_),
    .B1(_11573_),
    .Y(_11883_));
 sky130_fd_sc_hd__o21bai_2 _33523_ (.A1(_11877_),
    .A2(_11882_),
    .B1_N(_11883_),
    .Y(_11884_));
 sky130_fd_sc_hd__o21bai_2 _33524_ (.A1(_11879_),
    .A2(_11881_),
    .B1_N(_11876_),
    .Y(_11885_));
 sky130_fd_sc_hd__nand3_2 _33525_ (.A(_11868_),
    .B(_11876_),
    .C(_11872_),
    .Y(_11886_));
 sky130_fd_sc_hd__nand3_2 _33526_ (.A(_11885_),
    .B(_11883_),
    .C(_11886_),
    .Y(_11887_));
 sky130_fd_sc_hd__a21boi_2 _33527_ (.A1(_11263_),
    .A2(_11259_),
    .B1_N(_11574_),
    .Y(_11888_));
 sky130_fd_sc_hd__a21o_2 _33528_ (.A1(_11884_),
    .A2(_11887_),
    .B1(_11888_),
    .X(_11889_));
 sky130_fd_sc_hd__nand3_2 _33529_ (.A(_11884_),
    .B(_11888_),
    .C(_11887_),
    .Y(_11890_));
 sky130_fd_sc_hd__nand2_2 _33530_ (.A(_11589_),
    .B(_11581_),
    .Y(_11891_));
 sky130_fd_sc_hd__a21oi_2 _33531_ (.A1(_11889_),
    .A2(_11890_),
    .B1(_11891_),
    .Y(_11892_));
 sky130_fd_sc_hd__a21oi_2 _33532_ (.A1(_11884_),
    .A2(_11887_),
    .B1(_11888_),
    .Y(_11893_));
 sky130_fd_sc_hd__a21boi_2 _33533_ (.A1(_11586_),
    .A2(_11588_),
    .B1_N(_11581_),
    .Y(_11894_));
 sky130_vsdinv _33534_ (.A(_11890_),
    .Y(_11895_));
 sky130_fd_sc_hd__nor3_2 _33535_ (.A(_11893_),
    .B(_11894_),
    .C(_11895_),
    .Y(_11896_));
 sky130_fd_sc_hd__nor2_2 _33536_ (.A(_11892_),
    .B(_11896_),
    .Y(_11897_));
 sky130_fd_sc_hd__o21bai_2 _33537_ (.A1(_11591_),
    .A2(_11598_),
    .B1_N(_11593_),
    .Y(_11898_));
 sky130_fd_sc_hd__xor2_2 _33538_ (.A(_11897_),
    .B(_11898_),
    .X(_02654_));
 sky130_fd_sc_hd__nand2_2 _33539_ (.A(_10480_),
    .B(_05527_),
    .Y(_11899_));
 sky130_fd_sc_hd__nand3b_2 _33540_ (.A_N(_11899_),
    .B(_10996_),
    .C(_19282_),
    .Y(_11900_));
 sky130_fd_sc_hd__o21ai_2 _33541_ (.A1(_07794_),
    .A2(_16968_),
    .B1(_11899_),
    .Y(_11901_));
 sky130_fd_sc_hd__and2_2 _33542_ (.A(_18703_),
    .B(_05665_),
    .X(_11902_));
 sky130_fd_sc_hd__a21oi_2 _33543_ (.A1(_11900_),
    .A2(_11901_),
    .B1(_11902_),
    .Y(_11903_));
 sky130_fd_sc_hd__nand3_2 _33544_ (.A(_11900_),
    .B(_11902_),
    .C(_11901_),
    .Y(_11904_));
 sky130_vsdinv _33545_ (.A(_11904_),
    .Y(_11905_));
 sky130_fd_sc_hd__a21oi_2 _33546_ (.A1(_11606_),
    .A2(_11603_),
    .B1(_11602_),
    .Y(_11906_));
 sky130_fd_sc_hd__o21ai_2 _33547_ (.A1(_11903_),
    .A2(_11905_),
    .B1(_11906_),
    .Y(_11907_));
 sky130_fd_sc_hd__a21o_2 _33548_ (.A1(_11606_),
    .A2(_11603_),
    .B1(_11602_),
    .X(_11908_));
 sky130_fd_sc_hd__a22oi_2 _33549_ (.A1(_10487_),
    .A2(_05927_),
    .B1(_19282_),
    .B2(_10672_),
    .Y(_11909_));
 sky130_fd_sc_hd__nor3_2 _33550_ (.A(_07790_),
    .B(_11324_),
    .C(_11899_),
    .Y(_11910_));
 sky130_fd_sc_hd__o21bai_2 _33551_ (.A1(_11909_),
    .A2(_11910_),
    .B1_N(_11902_),
    .Y(_11911_));
 sky130_fd_sc_hd__nand3_2 _33552_ (.A(_11908_),
    .B(_11911_),
    .C(_11904_),
    .Y(_11912_));
 sky130_fd_sc_hd__nand2_2 _33553_ (.A(_10259_),
    .B(_05836_),
    .Y(_11913_));
 sky130_fd_sc_hd__nand2_2 _33554_ (.A(_10252_),
    .B(_05845_),
    .Y(_11914_));
 sky130_fd_sc_hd__nor2_2 _33555_ (.A(_11913_),
    .B(_11914_),
    .Y(_11915_));
 sky130_fd_sc_hd__nand2_2 _33556_ (.A(_11913_),
    .B(_11914_),
    .Y(_11916_));
 sky130_vsdinv _33557_ (.A(_11916_),
    .Y(_11917_));
 sky130_fd_sc_hd__and2_2 _33558_ (.A(_18722_),
    .B(_05949_),
    .X(_11918_));
 sky130_fd_sc_hd__o21bai_2 _33559_ (.A1(_11915_),
    .A2(_11917_),
    .B1_N(_11918_),
    .Y(_11919_));
 sky130_fd_sc_hd__nand3b_2 _33560_ (.A_N(_11915_),
    .B(_11918_),
    .C(_11916_),
    .Y(_11920_));
 sky130_fd_sc_hd__nand2_2 _33561_ (.A(_11919_),
    .B(_11920_),
    .Y(_11921_));
 sky130_vsdinv _33562_ (.A(_11921_),
    .Y(_11922_));
 sky130_fd_sc_hd__a21oi_2 _33563_ (.A1(_11907_),
    .A2(_11912_),
    .B1(_11922_),
    .Y(_11923_));
 sky130_fd_sc_hd__a21oi_2 _33564_ (.A1(_11911_),
    .A2(_11904_),
    .B1(_11908_),
    .Y(_11924_));
 sky130_fd_sc_hd__nor3_2 _33565_ (.A(_11906_),
    .B(_11903_),
    .C(_11905_),
    .Y(_11925_));
 sky130_fd_sc_hd__nor3_2 _33566_ (.A(_11921_),
    .B(_11924_),
    .C(_11925_),
    .Y(_11926_));
 sky130_fd_sc_hd__o21ai_2 _33567_ (.A1(_11621_),
    .A2(_11629_),
    .B1(_11611_),
    .Y(_11927_));
 sky130_fd_sc_hd__o21bai_2 _33568_ (.A1(_11923_),
    .A2(_11926_),
    .B1_N(_11927_),
    .Y(_11928_));
 sky130_fd_sc_hd__o21bai_2 _33569_ (.A1(_11924_),
    .A2(_11925_),
    .B1_N(_11922_),
    .Y(_11929_));
 sky130_fd_sc_hd__nand3_2 _33570_ (.A(_11907_),
    .B(_11922_),
    .C(_11912_),
    .Y(_11930_));
 sky130_fd_sc_hd__nand3_2 _33571_ (.A(_11929_),
    .B(_11930_),
    .C(_11927_),
    .Y(_11931_));
 sky130_fd_sc_hd__a22o_2 _33572_ (.A1(_11634_),
    .A2(_06357_),
    .B1(_10231_),
    .B2(_06886_),
    .X(_11932_));
 sky130_fd_sc_hd__nand2_2 _33573_ (.A(_09006_),
    .B(_07382_),
    .Y(_11933_));
 sky130_fd_sc_hd__nand3b_2 _33574_ (.A_N(_11933_),
    .B(_11636_),
    .C(_06203_),
    .Y(_11934_));
 sky130_fd_sc_hd__o2bb2ai_2 _33575_ (.A1_N(_11932_),
    .A2_N(_11934_),
    .B1(_09011_),
    .B2(_19243_),
    .Y(_11935_));
 sky130_fd_sc_hd__and2_2 _33576_ (.A(_08457_),
    .B(_06187_),
    .X(_11936_));
 sky130_fd_sc_hd__nand3_2 _33577_ (.A(_11934_),
    .B(_11932_),
    .C(_11936_),
    .Y(_11937_));
 sky130_fd_sc_hd__o31ai_2 _33578_ (.A1(_18724_),
    .A2(_19262_),
    .A3(_11613_),
    .B1(_11619_),
    .Y(_11938_));
 sky130_fd_sc_hd__a21oi_2 _33579_ (.A1(_11935_),
    .A2(_11937_),
    .B1(_11938_),
    .Y(_11939_));
 sky130_fd_sc_hd__nand3_2 _33580_ (.A(_11938_),
    .B(_11935_),
    .C(_11937_),
    .Y(_11940_));
 sky130_vsdinv _33581_ (.A(_11940_),
    .Y(_11941_));
 sky130_fd_sc_hd__a21boi_2 _33582_ (.A1(_11639_),
    .A2(_11633_),
    .B1_N(_11637_),
    .Y(_11942_));
 sky130_vsdinv _33583_ (.A(_11942_),
    .Y(_11943_));
 sky130_fd_sc_hd__o21bai_2 _33584_ (.A1(_11939_),
    .A2(_11941_),
    .B1_N(_11943_),
    .Y(_11944_));
 sky130_fd_sc_hd__nand3b_2 _33585_ (.A_N(_11939_),
    .B(_11943_),
    .C(_11940_),
    .Y(_11945_));
 sky130_fd_sc_hd__nand2_2 _33586_ (.A(_11944_),
    .B(_11945_),
    .Y(_11946_));
 sky130_fd_sc_hd__buf_1 _33587_ (.A(_11946_),
    .X(_11947_));
 sky130_fd_sc_hd__a21boi_2 _33588_ (.A1(_11928_),
    .A2(_11931_),
    .B1_N(_11947_),
    .Y(_11948_));
 sky130_fd_sc_hd__a21oi_2 _33589_ (.A1(_11929_),
    .A2(_11930_),
    .B1(_11927_),
    .Y(_11949_));
 sky130_vsdinv _33590_ (.A(_11931_),
    .Y(_11950_));
 sky130_fd_sc_hd__nor3_2 _33591_ (.A(_11947_),
    .B(_11949_),
    .C(_11950_),
    .Y(_11951_));
 sky130_fd_sc_hd__a21o_2 _33592_ (.A1(_11642_),
    .A2(_11644_),
    .B1(_11647_),
    .X(_11952_));
 sky130_fd_sc_hd__nand3_2 _33593_ (.A(_11647_),
    .B(_11642_),
    .C(_11644_),
    .Y(_11953_));
 sky130_fd_sc_hd__nand2_2 _33594_ (.A(_11952_),
    .B(_11953_),
    .Y(_11954_));
 sky130_fd_sc_hd__o21ai_2 _33595_ (.A1(_11954_),
    .A2(_11658_),
    .B1(_11632_),
    .Y(_11955_));
 sky130_fd_sc_hd__o21bai_2 _33596_ (.A1(_11948_),
    .A2(_11951_),
    .B1_N(_11955_),
    .Y(_11956_));
 sky130_fd_sc_hd__o21ai_2 _33597_ (.A1(_11949_),
    .A2(_11950_),
    .B1(_11947_),
    .Y(_11957_));
 sky130_fd_sc_hd__nand3b_2 _33598_ (.A_N(_11946_),
    .B(_11928_),
    .C(_11931_),
    .Y(_11958_));
 sky130_fd_sc_hd__nand3_2 _33599_ (.A(_11957_),
    .B(_11955_),
    .C(_11958_),
    .Y(_11959_));
 sky130_fd_sc_hd__buf_1 _33600_ (.A(_11959_),
    .X(_11960_));
 sky130_fd_sc_hd__a21oi_2 _33601_ (.A1(_11669_),
    .A2(_11668_),
    .B1(_11667_),
    .Y(_11961_));
 sky130_fd_sc_hd__nand2_2 _33602_ (.A(_18748_),
    .B(_06466_),
    .Y(_11962_));
 sky130_fd_sc_hd__nand2_2 _33603_ (.A(_09548_),
    .B(_07304_),
    .Y(_11963_));
 sky130_fd_sc_hd__nor2_2 _33604_ (.A(_11962_),
    .B(_11963_),
    .Y(_11964_));
 sky130_fd_sc_hd__and2_2 _33605_ (.A(_11080_),
    .B(_08262_),
    .X(_11965_));
 sky130_fd_sc_hd__nand2_2 _33606_ (.A(_11962_),
    .B(_11963_),
    .Y(_11966_));
 sky130_fd_sc_hd__nand3b_2 _33607_ (.A_N(_11964_),
    .B(_11965_),
    .C(_11966_),
    .Y(_11967_));
 sky130_fd_sc_hd__buf_1 _33608_ (.A(_09263_),
    .X(_11968_));
 sky130_fd_sc_hd__a22oi_2 _33609_ (.A1(_10417_),
    .A2(_06351_),
    .B1(_11968_),
    .B2(_07314_),
    .Y(_11969_));
 sky130_fd_sc_hd__o21bai_2 _33610_ (.A1(_11969_),
    .A2(_11964_),
    .B1_N(_11965_),
    .Y(_11970_));
 sky130_fd_sc_hd__nand3b_2 _33611_ (.A_N(_11961_),
    .B(_11967_),
    .C(_11970_),
    .Y(_11971_));
 sky130_fd_sc_hd__a21bo_2 _33612_ (.A1(_11967_),
    .A2(_11970_),
    .B1_N(_11961_),
    .X(_11972_));
 sky130_fd_sc_hd__and2_2 _33613_ (.A(_10436_),
    .B(_10376_),
    .X(_11973_));
 sky130_fd_sc_hd__nand2_2 _33614_ (.A(_08074_),
    .B(_08510_),
    .Y(_11974_));
 sky130_fd_sc_hd__nand2_2 _33615_ (.A(_07853_),
    .B(_07947_),
    .Y(_11975_));
 sky130_fd_sc_hd__xnor2_2 _33616_ (.A(_11974_),
    .B(_11975_),
    .Y(_11976_));
 sky130_fd_sc_hd__xnor2_2 _33617_ (.A(_11973_),
    .B(_11976_),
    .Y(_11977_));
 sky130_fd_sc_hd__a21o_2 _33618_ (.A1(_11971_),
    .A2(_11972_),
    .B1(_11977_),
    .X(_11978_));
 sky130_fd_sc_hd__nand3_2 _33619_ (.A(_11977_),
    .B(_11971_),
    .C(_11972_),
    .Y(_11979_));
 sky130_fd_sc_hd__o21ai_2 _33620_ (.A1(_11646_),
    .A2(_11649_),
    .B1(_11644_),
    .Y(_11980_));
 sky130_fd_sc_hd__a21oi_2 _33621_ (.A1(_11978_),
    .A2(_11979_),
    .B1(_11980_),
    .Y(_11981_));
 sky130_fd_sc_hd__nand3_2 _33622_ (.A(_11978_),
    .B(_11980_),
    .C(_11979_),
    .Y(_11982_));
 sky130_vsdinv _33623_ (.A(_11982_),
    .Y(_11983_));
 sky130_fd_sc_hd__nand2_2 _33624_ (.A(_11686_),
    .B(_11675_),
    .Y(_11984_));
 sky130_fd_sc_hd__o21bai_2 _33625_ (.A1(_11981_),
    .A2(_11983_),
    .B1_N(_11984_),
    .Y(_11985_));
 sky130_fd_sc_hd__nand3b_2 _33626_ (.A_N(_11981_),
    .B(_11984_),
    .C(_11982_),
    .Y(_11986_));
 sky130_fd_sc_hd__nand2_2 _33627_ (.A(_11985_),
    .B(_11986_),
    .Y(_11987_));
 sky130_fd_sc_hd__buf_1 _33628_ (.A(_11987_),
    .X(_11988_));
 sky130_fd_sc_hd__a21boi_2 _33629_ (.A1(_11956_),
    .A2(_11960_),
    .B1_N(_11988_),
    .Y(_11989_));
 sky130_fd_sc_hd__a21oi_2 _33630_ (.A1(_11957_),
    .A2(_11958_),
    .B1(_11955_),
    .Y(_11990_));
 sky130_fd_sc_hd__nor3b_2 _33631_ (.A(_11988_),
    .B(_11990_),
    .C_N(_11960_),
    .Y(_11991_));
 sky130_fd_sc_hd__o21ai_2 _33632_ (.A1(_11698_),
    .A2(_11700_),
    .B1(_11662_),
    .Y(_11992_));
 sky130_fd_sc_hd__o21bai_2 _33633_ (.A1(_11989_),
    .A2(_11991_),
    .B1_N(_11992_),
    .Y(_11993_));
 sky130_fd_sc_hd__nand2_2 _33634_ (.A(_11956_),
    .B(_11959_),
    .Y(_11994_));
 sky130_fd_sc_hd__nand2_2 _33635_ (.A(_11994_),
    .B(_11988_),
    .Y(_11995_));
 sky130_fd_sc_hd__nand3b_2 _33636_ (.A_N(_11987_),
    .B(_11956_),
    .C(_11960_),
    .Y(_11996_));
 sky130_fd_sc_hd__nand3_2 _33637_ (.A(_11995_),
    .B(_11992_),
    .C(_11996_),
    .Y(_11997_));
 sky130_fd_sc_hd__buf_1 _33638_ (.A(_11997_),
    .X(_11998_));
 sky130_fd_sc_hd__nand2_2 _33639_ (.A(_07006_),
    .B(_19203_),
    .Y(_11999_));
 sky130_fd_sc_hd__nand2_2 _33640_ (.A(_18785_),
    .B(_19196_),
    .Y(_12000_));
 sky130_fd_sc_hd__nor2_2 _33641_ (.A(_11999_),
    .B(_12000_),
    .Y(_12001_));
 sky130_vsdinv _33642_ (.A(_12001_),
    .Y(_12002_));
 sky130_fd_sc_hd__nand2_2 _33643_ (.A(_11999_),
    .B(_12000_),
    .Y(_12003_));
 sky130_fd_sc_hd__buf_1 _33644_ (.A(_19190_),
    .X(_12004_));
 sky130_fd_sc_hd__and2_2 _33645_ (.A(_06666_),
    .B(_12004_),
    .X(_12005_));
 sky130_fd_sc_hd__a21oi_2 _33646_ (.A1(_12002_),
    .A2(_12003_),
    .B1(_12005_),
    .Y(_12006_));
 sky130_fd_sc_hd__nand3b_2 _33647_ (.A_N(_12001_),
    .B(_12003_),
    .C(_12005_),
    .Y(_12007_));
 sky130_vsdinv _33648_ (.A(_12007_),
    .Y(_12008_));
 sky130_fd_sc_hd__o31ai_2 _33649_ (.A1(_18776_),
    .A2(_08524_),
    .A3(_11680_),
    .B1(_11679_),
    .Y(_12009_));
 sky130_fd_sc_hd__o21bai_2 _33650_ (.A1(_12006_),
    .A2(_12008_),
    .B1_N(_12009_),
    .Y(_12010_));
 sky130_fd_sc_hd__o2bb2ai_2 _33651_ (.A1_N(_12003_),
    .A2_N(_12002_),
    .B1(_08918_),
    .B2(_19192_),
    .Y(_12011_));
 sky130_fd_sc_hd__nand3_2 _33652_ (.A(_12011_),
    .B(_12009_),
    .C(_12007_),
    .Y(_12012_));
 sky130_fd_sc_hd__a21boi_2 _33653_ (.A1(_11718_),
    .A2(_11712_),
    .B1_N(_11715_),
    .Y(_12013_));
 sky130_vsdinv _33654_ (.A(_12013_),
    .Y(_12014_));
 sky130_fd_sc_hd__a21oi_2 _33655_ (.A1(_12010_),
    .A2(_12012_),
    .B1(_12014_),
    .Y(_12015_));
 sky130_fd_sc_hd__nand3_2 _33656_ (.A(_12010_),
    .B(_12014_),
    .C(_12012_),
    .Y(_12016_));
 sky130_vsdinv _33657_ (.A(_12016_),
    .Y(_12017_));
 sky130_fd_sc_hd__o21ai_2 _33658_ (.A1(_11728_),
    .A2(_11724_),
    .B1(_11725_),
    .Y(_12018_));
 sky130_fd_sc_hd__o21bai_2 _33659_ (.A1(_12015_),
    .A2(_12017_),
    .B1_N(_12018_),
    .Y(_12019_));
 sky130_fd_sc_hd__nand3b_2 _33660_ (.A_N(_12015_),
    .B(_12016_),
    .C(_12018_),
    .Y(_12020_));
 sky130_fd_sc_hd__nand2_2 _33661_ (.A(_12019_),
    .B(_12020_),
    .Y(_12021_));
 sky130_fd_sc_hd__a22o_2 _33662_ (.A1(_18798_),
    .A2(_08826_),
    .B1(_07824_),
    .B2(_11434_),
    .X(_12022_));
 sky130_fd_sc_hd__nand2_2 _33663_ (.A(_08032_),
    .B(_19185_),
    .Y(_12023_));
 sky130_fd_sc_hd__nand3b_2 _33664_ (.A_N(_12023_),
    .B(_06541_),
    .C(_09089_),
    .Y(_12024_));
 sky130_fd_sc_hd__o2bb2ai_2 _33665_ (.A1_N(_12022_),
    .A2_N(_12024_),
    .B1(_18809_),
    .B2(_19174_),
    .Y(_12025_));
 sky130_fd_sc_hd__and2_2 _33666_ (.A(_06275_),
    .B(_09497_),
    .X(_12026_));
 sky130_fd_sc_hd__nand3_2 _33667_ (.A(_12024_),
    .B(_12022_),
    .C(_12026_),
    .Y(_12027_));
 sky130_fd_sc_hd__nor2_2 _33668_ (.A(_11741_),
    .B(_11742_),
    .Y(_12028_));
 sky130_fd_sc_hd__a21oi_2 _33669_ (.A1(_11743_),
    .A2(_11747_),
    .B1(_12028_),
    .Y(_12029_));
 sky130_vsdinv _33670_ (.A(_12029_),
    .Y(_12030_));
 sky130_fd_sc_hd__a21oi_2 _33671_ (.A1(_12025_),
    .A2(_12027_),
    .B1(_12030_),
    .Y(_12031_));
 sky130_vsdinv _33672_ (.A(_12031_),
    .Y(_12032_));
 sky130_fd_sc_hd__nand3_2 _33673_ (.A(_12025_),
    .B(_12030_),
    .C(_12027_),
    .Y(_12033_));
 sky130_fd_sc_hd__nand2_2 _33674_ (.A(_12032_),
    .B(_12033_),
    .Y(_12034_));
 sky130_fd_sc_hd__buf_1 _33675_ (.A(_10532_),
    .X(_12035_));
 sky130_fd_sc_hd__and2_2 _33676_ (.A(_06816_),
    .B(_12035_),
    .X(_12036_));
 sky130_fd_sc_hd__nand2_2 _33677_ (.A(_18814_),
    .B(_09511_),
    .Y(_12037_));
 sky130_fd_sc_hd__nand2_2 _33678_ (.A(_11432_),
    .B(_11221_),
    .Y(_12038_));
 sky130_fd_sc_hd__xnor2_2 _33679_ (.A(_12037_),
    .B(_12038_),
    .Y(_12039_));
 sky130_fd_sc_hd__xor2_2 _33680_ (.A(_12036_),
    .B(_12039_),
    .X(_12040_));
 sky130_fd_sc_hd__nand2_2 _33681_ (.A(_12034_),
    .B(_12040_),
    .Y(_12041_));
 sky130_fd_sc_hd__nand3b_2 _33682_ (.A_N(_12040_),
    .B(_12032_),
    .C(_12033_),
    .Y(_12042_));
 sky130_fd_sc_hd__nand2_2 _33683_ (.A(_12041_),
    .B(_12042_),
    .Y(_12043_));
 sky130_fd_sc_hd__nand2_2 _33684_ (.A(_12021_),
    .B(_12043_),
    .Y(_12044_));
 sky130_fd_sc_hd__nand3b_2 _33685_ (.A_N(_12043_),
    .B(_12020_),
    .C(_12019_),
    .Y(_12045_));
 sky130_fd_sc_hd__nand2_2 _33686_ (.A(_12044_),
    .B(_12045_),
    .Y(_12046_));
 sky130_fd_sc_hd__a21boi_2 _33687_ (.A1(_11688_),
    .A2(_11695_),
    .B1_N(_11690_),
    .Y(_12047_));
 sky130_fd_sc_hd__nand2_2 _33688_ (.A(_12046_),
    .B(_12047_),
    .Y(_12048_));
 sky130_fd_sc_hd__nand2_2 _33689_ (.A(_11696_),
    .B(_11690_),
    .Y(_12049_));
 sky130_fd_sc_hd__nand3_2 _33690_ (.A(_12049_),
    .B(_12045_),
    .C(_12044_),
    .Y(_12050_));
 sky130_fd_sc_hd__nand2_2 _33691_ (.A(_12048_),
    .B(_12050_),
    .Y(_12051_));
 sky130_fd_sc_hd__a21boi_2 _33692_ (.A1(_11733_),
    .A2(_11759_),
    .B1_N(_11734_),
    .Y(_12052_));
 sky130_fd_sc_hd__nand2_2 _33693_ (.A(_12051_),
    .B(_12052_),
    .Y(_12053_));
 sky130_fd_sc_hd__nand3b_2 _33694_ (.A_N(_12052_),
    .B(_12048_),
    .C(_12050_),
    .Y(_12054_));
 sky130_fd_sc_hd__nand2_2 _33695_ (.A(_12053_),
    .B(_12054_),
    .Y(_12055_));
 sky130_fd_sc_hd__buf_1 _33696_ (.A(_12055_),
    .X(_12056_));
 sky130_fd_sc_hd__a21boi_2 _33697_ (.A1(_11993_),
    .A2(_11998_),
    .B1_N(_12056_),
    .Y(_12057_));
 sky130_fd_sc_hd__a21oi_2 _33698_ (.A1(_11995_),
    .A2(_11996_),
    .B1(_11992_),
    .Y(_12058_));
 sky130_fd_sc_hd__nor3b_2 _33699_ (.A(_12056_),
    .B(_12058_),
    .C_N(_11998_),
    .Y(_12059_));
 sky130_fd_sc_hd__o21ai_2 _33700_ (.A1(_11775_),
    .A2(_11776_),
    .B1(_11711_),
    .Y(_12060_));
 sky130_fd_sc_hd__o21bai_2 _33701_ (.A1(_12057_),
    .A2(_12059_),
    .B1_N(_12060_),
    .Y(_12061_));
 sky130_fd_sc_hd__nand2_2 _33702_ (.A(_11993_),
    .B(_11997_),
    .Y(_12062_));
 sky130_fd_sc_hd__nand2_2 _33703_ (.A(_12062_),
    .B(_12056_),
    .Y(_12063_));
 sky130_fd_sc_hd__nand3b_2 _33704_ (.A_N(_12055_),
    .B(_11998_),
    .C(_11993_),
    .Y(_12064_));
 sky130_fd_sc_hd__nand3_2 _33705_ (.A(_12063_),
    .B(_12060_),
    .C(_12064_),
    .Y(_12065_));
 sky130_fd_sc_hd__buf_1 _33706_ (.A(_12065_),
    .X(_12066_));
 sky130_fd_sc_hd__a22o_2 _33707_ (.A1(_05870_),
    .A2(_11515_),
    .B1(_06230_),
    .B2(_10894_),
    .X(_12067_));
 sky130_fd_sc_hd__nand2_2 _33708_ (.A(_05772_),
    .B(_09500_),
    .Y(_12068_));
 sky130_fd_sc_hd__buf_1 _33709_ (.A(_19143_),
    .X(_12069_));
 sky130_fd_sc_hd__nand3b_2 _33710_ (.A_N(_12068_),
    .B(_06227_),
    .C(_12069_),
    .Y(_12070_));
 sky130_fd_sc_hd__o2bb2ai_2 _33711_ (.A1_N(_12067_),
    .A2_N(_12070_),
    .B1(_07920_),
    .B2(_19140_),
    .Y(_12071_));
 sky130_fd_sc_hd__and2_2 _33712_ (.A(_06101_),
    .B(_11198_),
    .X(_12072_));
 sky130_fd_sc_hd__nand3_2 _33713_ (.A(_12070_),
    .B(_12067_),
    .C(_12072_),
    .Y(_12073_));
 sky130_fd_sc_hd__nand2_2 _33714_ (.A(_12071_),
    .B(_12073_),
    .Y(_12074_));
 sky130_vsdinv _33715_ (.A(_11737_),
    .Y(_12075_));
 sky130_fd_sc_hd__a21oi_2 _33716_ (.A1(_12075_),
    .A2(_11735_),
    .B1(_11738_),
    .Y(_12076_));
 sky130_fd_sc_hd__nand2_2 _33717_ (.A(_12074_),
    .B(_12076_),
    .Y(_12077_));
 sky130_fd_sc_hd__a21o_2 _33718_ (.A1(_12075_),
    .A2(_11735_),
    .B1(_11738_),
    .X(_12078_));
 sky130_fd_sc_hd__nand3_2 _33719_ (.A(_12078_),
    .B(_12071_),
    .C(_12073_),
    .Y(_12079_));
 sky130_fd_sc_hd__a21boi_2 _33720_ (.A1(_11786_),
    .A2(_11792_),
    .B1_N(_11789_),
    .Y(_12080_));
 sky130_vsdinv _33721_ (.A(_12080_),
    .Y(_12081_));
 sky130_fd_sc_hd__a21o_2 _33722_ (.A1(_12077_),
    .A2(_12079_),
    .B1(_12081_),
    .X(_12082_));
 sky130_fd_sc_hd__nand3_2 _33723_ (.A(_12077_),
    .B(_12079_),
    .C(_12081_),
    .Y(_12083_));
 sky130_fd_sc_hd__o21ai_2 _33724_ (.A1(_11752_),
    .A2(_11740_),
    .B1(_11754_),
    .Y(_12084_));
 sky130_fd_sc_hd__a21oi_2 _33725_ (.A1(_12082_),
    .A2(_12083_),
    .B1(_12084_),
    .Y(_12085_));
 sky130_fd_sc_hd__nand3_2 _33726_ (.A(_12082_),
    .B(_12084_),
    .C(_12083_),
    .Y(_12086_));
 sky130_vsdinv _33727_ (.A(_12086_),
    .Y(_12087_));
 sky130_fd_sc_hd__a21boi_2 _33728_ (.A1(_11797_),
    .A2(_11801_),
    .B1_N(_11799_),
    .Y(_12088_));
 sky130_vsdinv _33729_ (.A(_12088_),
    .Y(_12089_));
 sky130_fd_sc_hd__o21bai_2 _33730_ (.A1(_12085_),
    .A2(_12087_),
    .B1_N(_12089_),
    .Y(_12090_));
 sky130_fd_sc_hd__nand3b_2 _33731_ (.A_N(_12085_),
    .B(_12089_),
    .C(_12086_),
    .Y(_12091_));
 sky130_fd_sc_hd__nand2_2 _33732_ (.A(_12090_),
    .B(_12091_),
    .Y(_12092_));
 sky130_fd_sc_hd__a21boi_2 _33733_ (.A1(_11810_),
    .A2(_11812_),
    .B1_N(_11806_),
    .Y(_12093_));
 sky130_fd_sc_hd__nand2_2 _33734_ (.A(_12092_),
    .B(_12093_),
    .Y(_12094_));
 sky130_fd_sc_hd__nand2_2 _33735_ (.A(_11814_),
    .B(_11806_),
    .Y(_12095_));
 sky130_fd_sc_hd__nand3_2 _33736_ (.A(_12095_),
    .B(_12091_),
    .C(_12090_),
    .Y(_12096_));
 sky130_fd_sc_hd__buf_1 _33737_ (.A(\pcpi_mul.rs1[31] ),
    .X(_12097_));
 sky130_fd_sc_hd__nand2_2 _33738_ (.A(_18844_),
    .B(_12097_),
    .Y(_12098_));
 sky130_fd_sc_hd__buf_1 _33739_ (.A(_10881_),
    .X(_12099_));
 sky130_fd_sc_hd__nand2_2 _33740_ (.A(_12099_),
    .B(_05638_),
    .Y(_12100_));
 sky130_fd_sc_hd__xor2_2 _33741_ (.A(_12098_),
    .B(_12100_),
    .X(_12101_));
 sky130_fd_sc_hd__nand2_2 _33742_ (.A(_12101_),
    .B(_11188_),
    .Y(_12102_));
 sky130_fd_sc_hd__xnor2_2 _33743_ (.A(_12098_),
    .B(_12100_),
    .Y(_12103_));
 sky130_fd_sc_hd__nand2_2 _33744_ (.A(_12103_),
    .B(_10888_),
    .Y(_12104_));
 sky130_fd_sc_hd__nor2_2 _33745_ (.A(_11820_),
    .B(_11821_),
    .Y(_12105_));
 sky130_fd_sc_hd__a21oi_2 _33746_ (.A1(_11822_),
    .A2(_11188_),
    .B1(_12105_),
    .Y(_12106_));
 sky130_vsdinv _33747_ (.A(_12106_),
    .Y(_12107_));
 sky130_fd_sc_hd__a21o_2 _33748_ (.A1(_12102_),
    .A2(_12104_),
    .B1(_12107_),
    .X(_12108_));
 sky130_fd_sc_hd__nand3_2 _33749_ (.A(_12102_),
    .B(_12104_),
    .C(_12107_),
    .Y(_12109_));
 sky130_fd_sc_hd__buf_1 _33750_ (.A(_11834_),
    .X(_12110_));
 sky130_fd_sc_hd__a21o_2 _33751_ (.A1(_12108_),
    .A2(_12109_),
    .B1(_12110_),
    .X(_12111_));
 sky130_fd_sc_hd__nand3_2 _33752_ (.A(_12108_),
    .B(_12110_),
    .C(_12109_),
    .Y(_12112_));
 sky130_fd_sc_hd__a21boi_2 _33753_ (.A1(_11828_),
    .A2(_12110_),
    .B1_N(_11829_),
    .Y(_12113_));
 sky130_fd_sc_hd__a21bo_2 _33754_ (.A1(_12111_),
    .A2(_12112_),
    .B1_N(_12113_),
    .X(_12114_));
 sky130_fd_sc_hd__nand3b_2 _33755_ (.A_N(_12113_),
    .B(_12111_),
    .C(_12112_),
    .Y(_12115_));
 sky130_fd_sc_hd__a21oi_2 _33756_ (.A1(_11496_),
    .A2(_11831_),
    .B1(_11843_),
    .Y(_12116_));
 sky130_vsdinv _33757_ (.A(_12116_),
    .Y(_12117_));
 sky130_fd_sc_hd__buf_1 _33758_ (.A(_12117_),
    .X(_12118_));
 sky130_fd_sc_hd__a21oi_2 _33759_ (.A1(_12114_),
    .A2(_12115_),
    .B1(_12118_),
    .Y(_12119_));
 sky130_fd_sc_hd__nand3_2 _33760_ (.A(_12114_),
    .B(_12117_),
    .C(_12115_),
    .Y(_12120_));
 sky130_vsdinv _33761_ (.A(_12120_),
    .Y(_12121_));
 sky130_fd_sc_hd__nor2_2 _33762_ (.A(_12119_),
    .B(_12121_),
    .Y(_12122_));
 sky130_fd_sc_hd__a21oi_2 _33763_ (.A1(_12094_),
    .A2(_12096_),
    .B1(_12122_),
    .Y(_12123_));
 sky130_fd_sc_hd__or2b_2 _33764_ (.A(_12119_),
    .B_N(_12120_),
    .X(_12124_));
 sky130_fd_sc_hd__nand2_2 _33765_ (.A(_12094_),
    .B(_12096_),
    .Y(_12125_));
 sky130_fd_sc_hd__nor2_2 _33766_ (.A(_12124_),
    .B(_12125_),
    .Y(_12126_));
 sky130_fd_sc_hd__o21ai_2 _33767_ (.A1(_11765_),
    .A2(_11768_),
    .B1(_11764_),
    .Y(_12127_));
 sky130_fd_sc_hd__o21bai_2 _33768_ (.A1(_12123_),
    .A2(_12126_),
    .B1_N(_12127_),
    .Y(_12128_));
 sky130_fd_sc_hd__nand3_2 _33769_ (.A(_12122_),
    .B(_12094_),
    .C(_12096_),
    .Y(_12129_));
 sky130_fd_sc_hd__nand3b_2 _33770_ (.A_N(_12123_),
    .B(_12127_),
    .C(_12129_),
    .Y(_12130_));
 sky130_fd_sc_hd__buf_1 _33771_ (.A(_12130_),
    .X(_12131_));
 sky130_fd_sc_hd__o21a_2 _33772_ (.A1(_11848_),
    .A2(_11850_),
    .B1(_11819_),
    .X(_12132_));
 sky130_fd_sc_hd__a21boi_2 _33773_ (.A1(_12128_),
    .A2(_12131_),
    .B1_N(_12132_),
    .Y(_12133_));
 sky130_fd_sc_hd__nand2_2 _33774_ (.A(_12128_),
    .B(_12130_),
    .Y(_12134_));
 sky130_fd_sc_hd__nor2_2 _33775_ (.A(_12132_),
    .B(_12134_),
    .Y(_12135_));
 sky130_fd_sc_hd__nor2_2 _33776_ (.A(_12133_),
    .B(_12135_),
    .Y(_12136_));
 sky130_fd_sc_hd__a21oi_2 _33777_ (.A1(_12061_),
    .A2(_12066_),
    .B1(_12136_),
    .Y(_12137_));
 sky130_fd_sc_hd__nand2_2 _33778_ (.A(_12134_),
    .B(_12132_),
    .Y(_12138_));
 sky130_fd_sc_hd__nand3b_2 _33779_ (.A_N(_12132_),
    .B(_12128_),
    .C(_12131_),
    .Y(_12139_));
 sky130_fd_sc_hd__nand2_2 _33780_ (.A(_12138_),
    .B(_12139_),
    .Y(_12140_));
 sky130_fd_sc_hd__a21oi_2 _33781_ (.A1(_12063_),
    .A2(_12064_),
    .B1(_12060_),
    .Y(_12141_));
 sky130_fd_sc_hd__nor3b_2 _33782_ (.A(_12140_),
    .B(_12141_),
    .C_N(_12066_),
    .Y(_12142_));
 sky130_fd_sc_hd__o21ai_2 _33783_ (.A1(_11861_),
    .A2(_11864_),
    .B1(_11784_),
    .Y(_12143_));
 sky130_fd_sc_hd__o21bai_2 _33784_ (.A1(_12137_),
    .A2(_12142_),
    .B1_N(_12143_),
    .Y(_12144_));
 sky130_fd_sc_hd__nand2_2 _33785_ (.A(_12061_),
    .B(_12065_),
    .Y(_12145_));
 sky130_fd_sc_hd__nand2_2 _33786_ (.A(_12145_),
    .B(_12140_),
    .Y(_12146_));
 sky130_fd_sc_hd__nand3_2 _33787_ (.A(_12136_),
    .B(_12061_),
    .C(_12066_),
    .Y(_12147_));
 sky130_fd_sc_hd__nand3_2 _33788_ (.A(_12146_),
    .B(_12143_),
    .C(_12147_),
    .Y(_12148_));
 sky130_fd_sc_hd__buf_1 _33789_ (.A(_12148_),
    .X(_12149_));
 sky130_fd_sc_hd__and2_2 _33790_ (.A(_11846_),
    .B(_11841_),
    .X(_12150_));
 sky130_fd_sc_hd__nand2_2 _33791_ (.A(_11860_),
    .B(_11856_),
    .Y(_12151_));
 sky130_fd_sc_hd__xnor2_2 _33792_ (.A(_12150_),
    .B(_12151_),
    .Y(_12152_));
 sky130_fd_sc_hd__a21oi_2 _33793_ (.A1(_12144_),
    .A2(_12149_),
    .B1(_12152_),
    .Y(_12153_));
 sky130_vsdinv _33794_ (.A(_12152_),
    .Y(_12154_));
 sky130_fd_sc_hd__a21oi_2 _33795_ (.A1(_12146_),
    .A2(_12147_),
    .B1(_12143_),
    .Y(_12155_));
 sky130_fd_sc_hd__nor3b_2 _33796_ (.A(_12154_),
    .B(_12155_),
    .C_N(_12149_),
    .Y(_12156_));
 sky130_fd_sc_hd__o21ai_2 _33797_ (.A1(_11878_),
    .A2(_11879_),
    .B1(_11872_),
    .Y(_12157_));
 sky130_fd_sc_hd__o21bai_2 _33798_ (.A1(_12153_),
    .A2(_12156_),
    .B1_N(_12157_),
    .Y(_12158_));
 sky130_fd_sc_hd__nand2_2 _33799_ (.A(_12144_),
    .B(_12148_),
    .Y(_12159_));
 sky130_fd_sc_hd__nand2_2 _33800_ (.A(_12159_),
    .B(_12154_),
    .Y(_12160_));
 sky130_fd_sc_hd__nand3_2 _33801_ (.A(_12144_),
    .B(_12152_),
    .C(_12149_),
    .Y(_12161_));
 sky130_fd_sc_hd__nand3_2 _33802_ (.A(_12160_),
    .B(_12157_),
    .C(_12161_),
    .Y(_12162_));
 sky130_fd_sc_hd__o21a_2 _33803_ (.A1(_11873_),
    .A2(_11551_),
    .B1(_11875_),
    .X(_12163_));
 sky130_fd_sc_hd__a21oi_2 _33804_ (.A1(_12158_),
    .A2(_12162_),
    .B1(_12163_),
    .Y(_12164_));
 sky130_vsdinv _33805_ (.A(_12163_),
    .Y(_12165_));
 sky130_fd_sc_hd__a21oi_2 _33806_ (.A1(_12160_),
    .A2(_12161_),
    .B1(_12157_),
    .Y(_12166_));
 sky130_vsdinv _33807_ (.A(_12162_),
    .Y(_12167_));
 sky130_fd_sc_hd__nor3_2 _33808_ (.A(_12165_),
    .B(_12166_),
    .C(_12167_),
    .Y(_12168_));
 sky130_vsdinv _33809_ (.A(_11888_),
    .Y(_12169_));
 sky130_fd_sc_hd__a21oi_2 _33810_ (.A1(_11885_),
    .A2(_11886_),
    .B1(_11883_),
    .Y(_12170_));
 sky130_fd_sc_hd__o21ai_2 _33811_ (.A1(_12169_),
    .A2(_12170_),
    .B1(_11887_),
    .Y(_12171_));
 sky130_fd_sc_hd__o21bai_2 _33812_ (.A1(_12164_),
    .A2(_12168_),
    .B1_N(_12171_),
    .Y(_12172_));
 sky130_fd_sc_hd__o21bai_2 _33813_ (.A1(_12166_),
    .A2(_12167_),
    .B1_N(_12163_),
    .Y(_12173_));
 sky130_fd_sc_hd__nand3_2 _33814_ (.A(_12158_),
    .B(_12163_),
    .C(_12162_),
    .Y(_12174_));
 sky130_fd_sc_hd__nand3_2 _33815_ (.A(_12173_),
    .B(_12171_),
    .C(_12174_),
    .Y(_12175_));
 sky130_fd_sc_hd__nand2_2 _33816_ (.A(_12172_),
    .B(_12175_),
    .Y(_12176_));
 sky130_fd_sc_hd__nand3_2 _33817_ (.A(_11595_),
    .B(_11594_),
    .C(_11897_),
    .Y(_12177_));
 sky130_fd_sc_hd__a31o_2 _33818_ (.A1(_10978_),
    .A2(_10979_),
    .A3(_10991_),
    .B1(_12177_),
    .X(_12178_));
 sky130_fd_sc_hd__nand3_2 _33819_ (.A(_11594_),
    .B(_11897_),
    .C(_11597_),
    .Y(_12179_));
 sky130_fd_sc_hd__nand3_2 _33820_ (.A(_11891_),
    .B(_11889_),
    .C(_11890_),
    .Y(_12180_));
 sky130_fd_sc_hd__o21a_2 _33821_ (.A1(_11592_),
    .A2(_11892_),
    .B1(_12180_),
    .X(_12181_));
 sky130_fd_sc_hd__and3_2 _33822_ (.A(_12178_),
    .B(_12179_),
    .C(_12181_),
    .X(_12182_));
 sky130_fd_sc_hd__xor2_2 _33823_ (.A(_12176_),
    .B(_12182_),
    .X(_02655_));
 sky130_fd_sc_hd__buf_1 _33824_ (.A(_10671_),
    .X(_12183_));
 sky130_fd_sc_hd__a22oi_2 _33825_ (.A1(_10669_),
    .A2(_05851_),
    .B1(_19278_),
    .B2(_12183_),
    .Y(_12184_));
 sky130_fd_sc_hd__nand2_2 _33826_ (.A(_10486_),
    .B(_08480_),
    .Y(_12185_));
 sky130_fd_sc_hd__nor3_2 _33827_ (.A(_05536_),
    .B(_11004_),
    .C(_12185_),
    .Y(_12186_));
 sky130_fd_sc_hd__and2_2 _33828_ (.A(_10266_),
    .B(_06979_),
    .X(_12187_));
 sky130_fd_sc_hd__o21bai_2 _33829_ (.A1(_12184_),
    .A2(_12186_),
    .B1_N(_12187_),
    .Y(_12188_));
 sky130_fd_sc_hd__nand3b_2 _33830_ (.A_N(_12185_),
    .B(_10672_),
    .C(_19278_),
    .Y(_12189_));
 sky130_fd_sc_hd__o21ai_2 _33831_ (.A1(_05536_),
    .A2(_11324_),
    .B1(_12185_),
    .Y(_12190_));
 sky130_fd_sc_hd__nand3_2 _33832_ (.A(_12189_),
    .B(_12187_),
    .C(_12190_),
    .Y(_12191_));
 sky130_fd_sc_hd__a21o_2 _33833_ (.A1(_11901_),
    .A2(_11902_),
    .B1(_11910_),
    .X(_12192_));
 sky130_fd_sc_hd__a21o_2 _33834_ (.A1(_12188_),
    .A2(_12191_),
    .B1(_12192_),
    .X(_12193_));
 sky130_fd_sc_hd__nand3_2 _33835_ (.A(_12192_),
    .B(_12188_),
    .C(_12191_),
    .Y(_12194_));
 sky130_fd_sc_hd__buf_1 _33836_ (.A(_12194_),
    .X(_12195_));
 sky130_fd_sc_hd__a22oi_2 _33837_ (.A1(_18710_),
    .A2(_07375_),
    .B1(_11612_),
    .B2(_05821_),
    .Y(_12196_));
 sky130_fd_sc_hd__and4_2 _33838_ (.A(_11014_),
    .B(_11612_),
    .C(_07216_),
    .D(_06074_),
    .X(_12197_));
 sky130_fd_sc_hd__and2_2 _33839_ (.A(_09605_),
    .B(_19252_),
    .X(_12198_));
 sky130_fd_sc_hd__o21bai_2 _33840_ (.A1(_12196_),
    .A2(_12197_),
    .B1_N(_12198_),
    .Y(_12199_));
 sky130_fd_sc_hd__nand2_2 _33841_ (.A(_09957_),
    .B(_07375_),
    .Y(_12200_));
 sky130_fd_sc_hd__nand3b_2 _33842_ (.A_N(_12200_),
    .B(_10253_),
    .C(_05950_),
    .Y(_12201_));
 sky130_fd_sc_hd__nand3b_2 _33843_ (.A_N(_12196_),
    .B(_12201_),
    .C(_12198_),
    .Y(_12202_));
 sky130_fd_sc_hd__nand2_2 _33844_ (.A(_12199_),
    .B(_12202_),
    .Y(_12203_));
 sky130_vsdinv _33845_ (.A(_12203_),
    .Y(_12204_));
 sky130_fd_sc_hd__a21oi_2 _33846_ (.A1(_12193_),
    .A2(_12195_),
    .B1(_12204_),
    .Y(_12205_));
 sky130_fd_sc_hd__a21oi_2 _33847_ (.A1(_12188_),
    .A2(_12191_),
    .B1(_12192_),
    .Y(_12206_));
 sky130_fd_sc_hd__nor3b_2 _33848_ (.A(_12203_),
    .B(_12206_),
    .C_N(_12195_),
    .Y(_12207_));
 sky130_fd_sc_hd__o21ai_2 _33849_ (.A1(_11921_),
    .A2(_11924_),
    .B1(_11912_),
    .Y(_12208_));
 sky130_fd_sc_hd__o21bai_2 _33850_ (.A1(_12205_),
    .A2(_12207_),
    .B1_N(_12208_),
    .Y(_12209_));
 sky130_vsdinv _33851_ (.A(_12194_),
    .Y(_12210_));
 sky130_fd_sc_hd__o21bai_2 _33852_ (.A1(_12206_),
    .A2(_12210_),
    .B1_N(_12204_),
    .Y(_12211_));
 sky130_fd_sc_hd__nand3_2 _33853_ (.A(_12193_),
    .B(_12204_),
    .C(_12195_),
    .Y(_12212_));
 sky130_fd_sc_hd__nand3_2 _33854_ (.A(_12211_),
    .B(_12212_),
    .C(_12208_),
    .Y(_12213_));
 sky130_fd_sc_hd__buf_1 _33855_ (.A(_12213_),
    .X(_12214_));
 sky130_fd_sc_hd__a22o_2 _33856_ (.A1(_09312_),
    .A2(_06203_),
    .B1(_10456_),
    .B2(_06478_),
    .X(_12215_));
 sky130_fd_sc_hd__nand2_2 _33857_ (.A(_18728_),
    .B(_09341_),
    .Y(_12216_));
 sky130_fd_sc_hd__buf_1 _33858_ (.A(_10453_),
    .X(_12217_));
 sky130_fd_sc_hd__nand3b_2 _33859_ (.A_N(_12216_),
    .B(_12217_),
    .C(_06464_),
    .Y(_12218_));
 sky130_fd_sc_hd__buf_1 _33860_ (.A(_10245_),
    .X(_12219_));
 sky130_fd_sc_hd__o2bb2ai_2 _33861_ (.A1_N(_12215_),
    .A2_N(_12218_),
    .B1(_12219_),
    .B2(_19238_),
    .Y(_12220_));
 sky130_fd_sc_hd__and2_2 _33862_ (.A(_08759_),
    .B(_06616_),
    .X(_12221_));
 sky130_fd_sc_hd__nand3_2 _33863_ (.A(_12218_),
    .B(_12215_),
    .C(_12221_),
    .Y(_12222_));
 sky130_fd_sc_hd__a21oi_2 _33864_ (.A1(_11916_),
    .A2(_11918_),
    .B1(_11915_),
    .Y(_12223_));
 sky130_vsdinv _33865_ (.A(_12223_),
    .Y(_12224_));
 sky130_fd_sc_hd__a21o_2 _33866_ (.A1(_12220_),
    .A2(_12222_),
    .B1(_12224_),
    .X(_12225_));
 sky130_fd_sc_hd__nand3_2 _33867_ (.A(_12220_),
    .B(_12224_),
    .C(_12222_),
    .Y(_12226_));
 sky130_fd_sc_hd__a21boi_2 _33868_ (.A1(_11936_),
    .A2(_11932_),
    .B1_N(_11934_),
    .Y(_12227_));
 sky130_vsdinv _33869_ (.A(_12227_),
    .Y(_12228_));
 sky130_fd_sc_hd__a21o_2 _33870_ (.A1(_12225_),
    .A2(_12226_),
    .B1(_12228_),
    .X(_12229_));
 sky130_fd_sc_hd__nand3_2 _33871_ (.A(_12225_),
    .B(_12228_),
    .C(_12226_),
    .Y(_12230_));
 sky130_fd_sc_hd__nand2_2 _33872_ (.A(_12229_),
    .B(_12230_),
    .Y(_12231_));
 sky130_fd_sc_hd__buf_1 _33873_ (.A(_12231_),
    .X(_12232_));
 sky130_fd_sc_hd__a21boi_2 _33874_ (.A1(_12209_),
    .A2(_12214_),
    .B1_N(_12232_),
    .Y(_12233_));
 sky130_fd_sc_hd__a21oi_2 _33875_ (.A1(_12211_),
    .A2(_12212_),
    .B1(_12208_),
    .Y(_12234_));
 sky130_fd_sc_hd__nor3b_2 _33876_ (.A(_12232_),
    .B(_12234_),
    .C_N(_12214_),
    .Y(_12235_));
 sky130_fd_sc_hd__o21ai_2 _33877_ (.A1(_11947_),
    .A2(_11949_),
    .B1(_11931_),
    .Y(_12236_));
 sky130_fd_sc_hd__o21bai_2 _33878_ (.A1(_12233_),
    .A2(_12235_),
    .B1_N(_12236_),
    .Y(_12237_));
 sky130_fd_sc_hd__nand2_2 _33879_ (.A(_12209_),
    .B(_12213_),
    .Y(_12238_));
 sky130_fd_sc_hd__nand2_2 _33880_ (.A(_12238_),
    .B(_12232_),
    .Y(_12239_));
 sky130_fd_sc_hd__nand3b_2 _33881_ (.A_N(_12231_),
    .B(_12209_),
    .C(_12214_),
    .Y(_12240_));
 sky130_fd_sc_hd__nand3_2 _33882_ (.A(_12239_),
    .B(_12240_),
    .C(_12236_),
    .Y(_12241_));
 sky130_fd_sc_hd__nand2_2 _33883_ (.A(_08472_),
    .B(_06453_),
    .Y(_12242_));
 sky130_fd_sc_hd__nand2_2 _33884_ (.A(_08473_),
    .B(_06745_),
    .Y(_12243_));
 sky130_fd_sc_hd__nor2_2 _33885_ (.A(_12242_),
    .B(_12243_),
    .Y(_12244_));
 sky130_fd_sc_hd__and2_2 _33886_ (.A(_08084_),
    .B(_08255_),
    .X(_12245_));
 sky130_fd_sc_hd__nand2_2 _33887_ (.A(_12242_),
    .B(_12243_),
    .Y(_12246_));
 sky130_fd_sc_hd__nand3b_2 _33888_ (.A_N(_12244_),
    .B(_12245_),
    .C(_12246_),
    .Y(_12247_));
 sky130_fd_sc_hd__a22oi_2 _33889_ (.A1(_18749_),
    .A2(_06454_),
    .B1(_11074_),
    .B2(_07913_),
    .Y(_12248_));
 sky130_fd_sc_hd__o21bai_2 _33890_ (.A1(_12248_),
    .A2(_12244_),
    .B1_N(_12245_),
    .Y(_12249_));
 sky130_fd_sc_hd__a21oi_2 _33891_ (.A1(_11966_),
    .A2(_11965_),
    .B1(_11964_),
    .Y(_12250_));
 sky130_fd_sc_hd__a21bo_2 _33892_ (.A1(_12247_),
    .A2(_12249_),
    .B1_N(_12250_),
    .X(_12251_));
 sky130_fd_sc_hd__nand3b_2 _33893_ (.A_N(_12250_),
    .B(_12247_),
    .C(_12249_),
    .Y(_12252_));
 sky130_fd_sc_hd__nand2_2 _33894_ (.A(_10745_),
    .B(_07947_),
    .Y(_12253_));
 sky130_fd_sc_hd__buf_1 _33895_ (.A(_18770_),
    .X(_12254_));
 sky130_fd_sc_hd__nand2_2 _33896_ (.A(_12254_),
    .B(_07106_),
    .Y(_12255_));
 sky130_fd_sc_hd__nand2_2 _33897_ (.A(_12253_),
    .B(_12255_),
    .Y(_12256_));
 sky130_fd_sc_hd__nor2_2 _33898_ (.A(_12253_),
    .B(_12255_),
    .Y(_12257_));
 sky130_vsdinv _33899_ (.A(_12257_),
    .Y(_12258_));
 sky130_fd_sc_hd__o2bb2ai_2 _33900_ (.A1_N(_12256_),
    .A2_N(_12258_),
    .B1(_18777_),
    .B2(_09665_),
    .Y(_12259_));
 sky130_fd_sc_hd__and2_2 _33901_ (.A(_07421_),
    .B(_08303_),
    .X(_12260_));
 sky130_fd_sc_hd__nand3b_2 _33902_ (.A_N(_12257_),
    .B(_12260_),
    .C(_12256_),
    .Y(_12261_));
 sky130_fd_sc_hd__nand2_2 _33903_ (.A(_12259_),
    .B(_12261_),
    .Y(_12262_));
 sky130_fd_sc_hd__a21boi_2 _33904_ (.A1(_12251_),
    .A2(_12252_),
    .B1_N(_12262_),
    .Y(_12263_));
 sky130_vsdinv _33905_ (.A(_12252_),
    .Y(_12264_));
 sky130_fd_sc_hd__nor3b_2 _33906_ (.A(_12262_),
    .B(_12264_),
    .C_N(_12251_),
    .Y(_12265_));
 sky130_fd_sc_hd__o21ai_2 _33907_ (.A1(_11942_),
    .A2(_11939_),
    .B1(_11940_),
    .Y(_12266_));
 sky130_fd_sc_hd__o21bai_2 _33908_ (.A1(_12263_),
    .A2(_12265_),
    .B1_N(_12266_),
    .Y(_12267_));
 sky130_fd_sc_hd__nand3b_2 _33909_ (.A_N(_12262_),
    .B(_12252_),
    .C(_12251_),
    .Y(_12268_));
 sky130_fd_sc_hd__nand3b_2 _33910_ (.A_N(_12263_),
    .B(_12266_),
    .C(_12268_),
    .Y(_12269_));
 sky130_fd_sc_hd__a21boi_2 _33911_ (.A1(_11977_),
    .A2(_11972_),
    .B1_N(_11971_),
    .Y(_12270_));
 sky130_vsdinv _33912_ (.A(_12270_),
    .Y(_12271_));
 sky130_fd_sc_hd__a21oi_2 _33913_ (.A1(_12267_),
    .A2(_12269_),
    .B1(_12271_),
    .Y(_12272_));
 sky130_fd_sc_hd__nand3_2 _33914_ (.A(_12267_),
    .B(_12269_),
    .C(_12271_),
    .Y(_12273_));
 sky130_vsdinv _33915_ (.A(_12273_),
    .Y(_12274_));
 sky130_fd_sc_hd__nor2_2 _33916_ (.A(_12272_),
    .B(_12274_),
    .Y(_12275_));
 sky130_fd_sc_hd__a21oi_2 _33917_ (.A1(_12237_),
    .A2(_12241_),
    .B1(_12275_),
    .Y(_12276_));
 sky130_fd_sc_hd__a21o_2 _33918_ (.A1(_12267_),
    .A2(_12269_),
    .B1(_12271_),
    .X(_12277_));
 sky130_fd_sc_hd__nand2_2 _33919_ (.A(_12277_),
    .B(_12273_),
    .Y(_12278_));
 sky130_fd_sc_hd__a21oi_2 _33920_ (.A1(_12239_),
    .A2(_12240_),
    .B1(_12236_),
    .Y(_12279_));
 sky130_vsdinv _33921_ (.A(_12241_),
    .Y(_12280_));
 sky130_fd_sc_hd__nor3_2 _33922_ (.A(_12278_),
    .B(_12279_),
    .C(_12280_),
    .Y(_12281_));
 sky130_fd_sc_hd__o21ai_2 _33923_ (.A1(_11988_),
    .A2(_11990_),
    .B1(_11960_),
    .Y(_12282_));
 sky130_fd_sc_hd__o21bai_2 _33924_ (.A1(_12276_),
    .A2(_12281_),
    .B1_N(_12282_),
    .Y(_12283_));
 sky130_fd_sc_hd__o21bai_2 _33925_ (.A1(_12279_),
    .A2(_12280_),
    .B1_N(_12275_),
    .Y(_12284_));
 sky130_fd_sc_hd__nand3_2 _33926_ (.A(_12237_),
    .B(_12275_),
    .C(_12241_),
    .Y(_12285_));
 sky130_fd_sc_hd__nand3_2 _33927_ (.A(_12284_),
    .B(_12285_),
    .C(_12282_),
    .Y(_12286_));
 sky130_fd_sc_hd__buf_1 _33928_ (.A(_12286_),
    .X(_12287_));
 sky130_fd_sc_hd__buf_1 _33929_ (.A(_07591_),
    .X(_12288_));
 sky130_fd_sc_hd__buf_1 _33930_ (.A(_08391_),
    .X(_12289_));
 sky130_fd_sc_hd__a22o_2 _33931_ (.A1(_18781_),
    .A2(_12288_),
    .B1(_12289_),
    .B2(_08571_),
    .X(_12290_));
 sky130_fd_sc_hd__nand2_2 _33932_ (.A(_08011_),
    .B(_07752_),
    .Y(_12291_));
 sky130_fd_sc_hd__buf_1 _33933_ (.A(_12004_),
    .X(_12292_));
 sky130_fd_sc_hd__nand3b_2 _33934_ (.A_N(_12291_),
    .B(_10774_),
    .C(_12292_),
    .Y(_12293_));
 sky130_fd_sc_hd__o2bb2ai_2 _33935_ (.A1_N(_12290_),
    .A2_N(_12293_),
    .B1(_07400_),
    .B2(_19187_),
    .Y(_12294_));
 sky130_fd_sc_hd__buf_1 _33936_ (.A(_08565_),
    .X(_12295_));
 sky130_fd_sc_hd__and2_2 _33937_ (.A(_11409_),
    .B(_12295_),
    .X(_12296_));
 sky130_fd_sc_hd__nand3_2 _33938_ (.A(_12293_),
    .B(_12290_),
    .C(_12296_),
    .Y(_12297_));
 sky130_fd_sc_hd__nand2_2 _33939_ (.A(_11974_),
    .B(_11975_),
    .Y(_12298_));
 sky130_fd_sc_hd__nor2_2 _33940_ (.A(_11974_),
    .B(_11975_),
    .Y(_12299_));
 sky130_fd_sc_hd__a21oi_2 _33941_ (.A1(_12298_),
    .A2(_11973_),
    .B1(_12299_),
    .Y(_12300_));
 sky130_vsdinv _33942_ (.A(_12300_),
    .Y(_12301_));
 sky130_fd_sc_hd__a21o_2 _33943_ (.A1(_12294_),
    .A2(_12297_),
    .B1(_12301_),
    .X(_12302_));
 sky130_fd_sc_hd__nand3_2 _33944_ (.A(_12294_),
    .B(_12301_),
    .C(_12297_),
    .Y(_12303_));
 sky130_fd_sc_hd__buf_1 _33945_ (.A(_12303_),
    .X(_12304_));
 sky130_fd_sc_hd__a21oi_2 _33946_ (.A1(_12003_),
    .A2(_12005_),
    .B1(_12001_),
    .Y(_12305_));
 sky130_vsdinv _33947_ (.A(_12305_),
    .Y(_12306_));
 sky130_fd_sc_hd__a21oi_2 _33948_ (.A1(_12302_),
    .A2(_12304_),
    .B1(_12306_),
    .Y(_12307_));
 sky130_fd_sc_hd__a21oi_2 _33949_ (.A1(_12294_),
    .A2(_12297_),
    .B1(_12301_),
    .Y(_12308_));
 sky130_fd_sc_hd__nor3b_2 _33950_ (.A(_12305_),
    .B(_12308_),
    .C_N(_12303_),
    .Y(_12309_));
 sky130_fd_sc_hd__a21oi_2 _33951_ (.A1(_12011_),
    .A2(_12007_),
    .B1(_12009_),
    .Y(_12310_));
 sky130_fd_sc_hd__o21ai_2 _33952_ (.A1(_12013_),
    .A2(_12310_),
    .B1(_12012_),
    .Y(_12311_));
 sky130_fd_sc_hd__o21bai_2 _33953_ (.A1(_12307_),
    .A2(_12309_),
    .B1_N(_12311_),
    .Y(_12312_));
 sky130_fd_sc_hd__a21o_2 _33954_ (.A1(_12302_),
    .A2(_12304_),
    .B1(_12306_),
    .X(_12313_));
 sky130_fd_sc_hd__nand3_2 _33955_ (.A(_12302_),
    .B(_12306_),
    .C(_12304_),
    .Y(_12314_));
 sky130_fd_sc_hd__nand3_2 _33956_ (.A(_12313_),
    .B(_12311_),
    .C(_12314_),
    .Y(_12315_));
 sky130_fd_sc_hd__buf_1 _33957_ (.A(_19149_),
    .X(_12316_));
 sky130_fd_sc_hd__and2_2 _33958_ (.A(_06138_),
    .B(_12316_),
    .X(_12317_));
 sky130_fd_sc_hd__nand2_2 _33959_ (.A(_06148_),
    .B(_10531_),
    .Y(_12318_));
 sky130_fd_sc_hd__nand2_2 _33960_ (.A(_06142_),
    .B(_12035_),
    .Y(_12319_));
 sky130_fd_sc_hd__xnor2_2 _33961_ (.A(_12318_),
    .B(_12319_),
    .Y(_12320_));
 sky130_fd_sc_hd__xor2_2 _33962_ (.A(_12317_),
    .B(_12320_),
    .X(_12321_));
 sky130_fd_sc_hd__nand2_2 _33963_ (.A(_08170_),
    .B(_10077_),
    .Y(_12322_));
 sky130_fd_sc_hd__nand2_2 _33964_ (.A(_06393_),
    .B(_10843_),
    .Y(_12323_));
 sky130_fd_sc_hd__nor2_2 _33965_ (.A(_12322_),
    .B(_12323_),
    .Y(_12324_));
 sky130_fd_sc_hd__buf_1 _33966_ (.A(_08818_),
    .X(_12325_));
 sky130_fd_sc_hd__and2_2 _33967_ (.A(_06551_),
    .B(_12325_),
    .X(_12326_));
 sky130_fd_sc_hd__nand2_2 _33968_ (.A(_12322_),
    .B(_12323_),
    .Y(_12327_));
 sky130_fd_sc_hd__nand3b_2 _33969_ (.A_N(_12324_),
    .B(_12326_),
    .C(_12327_),
    .Y(_12328_));
 sky130_fd_sc_hd__buf_1 _33970_ (.A(_10575_),
    .X(_12329_));
 sky130_fd_sc_hd__buf_1 _33971_ (.A(_10843_),
    .X(_12330_));
 sky130_fd_sc_hd__a22oi_2 _33972_ (.A1(_18799_),
    .A2(_12329_),
    .B1(_18804_),
    .B2(_12330_),
    .Y(_12331_));
 sky130_fd_sc_hd__o21bai_2 _33973_ (.A1(_12331_),
    .A2(_12324_),
    .B1_N(_12326_),
    .Y(_12332_));
 sky130_fd_sc_hd__nand2_2 _33974_ (.A(_12027_),
    .B(_12024_),
    .Y(_12333_));
 sky130_fd_sc_hd__a21o_2 _33975_ (.A1(_12328_),
    .A2(_12332_),
    .B1(_12333_),
    .X(_12334_));
 sky130_fd_sc_hd__nand3_2 _33976_ (.A(_12333_),
    .B(_12328_),
    .C(_12332_),
    .Y(_12335_));
 sky130_fd_sc_hd__nand2_2 _33977_ (.A(_12334_),
    .B(_12335_),
    .Y(_12336_));
 sky130_fd_sc_hd__xor2_2 _33978_ (.A(_12321_),
    .B(_12336_),
    .X(_12337_));
 sky130_fd_sc_hd__a21oi_2 _33979_ (.A1(_12312_),
    .A2(_12315_),
    .B1(_12337_),
    .Y(_12338_));
 sky130_fd_sc_hd__xnor2_2 _33980_ (.A(_12321_),
    .B(_12336_),
    .Y(_12339_));
 sky130_fd_sc_hd__nand2_2 _33981_ (.A(_12312_),
    .B(_12315_),
    .Y(_12340_));
 sky130_fd_sc_hd__nor2_2 _33982_ (.A(_12339_),
    .B(_12340_),
    .Y(_12341_));
 sky130_fd_sc_hd__a21boi_2 _33983_ (.A1(_11685_),
    .A2(_11674_),
    .B1_N(_11675_),
    .Y(_12342_));
 sky130_fd_sc_hd__o21ai_2 _33984_ (.A1(_12342_),
    .A2(_11981_),
    .B1(_11982_),
    .Y(_12343_));
 sky130_fd_sc_hd__o21bai_2 _33985_ (.A1(_12338_),
    .A2(_12341_),
    .B1_N(_12343_),
    .Y(_12344_));
 sky130_fd_sc_hd__nand2_2 _33986_ (.A(_12340_),
    .B(_12339_),
    .Y(_12345_));
 sky130_fd_sc_hd__nand3_2 _33987_ (.A(_12337_),
    .B(_12312_),
    .C(_12315_),
    .Y(_12346_));
 sky130_fd_sc_hd__nand3_2 _33988_ (.A(_12345_),
    .B(_12343_),
    .C(_12346_),
    .Y(_12347_));
 sky130_vsdinv _33989_ (.A(_12043_),
    .Y(_12348_));
 sky130_fd_sc_hd__a21boi_2 _33990_ (.A1(_12348_),
    .A2(_12019_),
    .B1_N(_12020_),
    .Y(_12349_));
 sky130_vsdinv _33991_ (.A(_12349_),
    .Y(_12350_));
 sky130_fd_sc_hd__a21oi_2 _33992_ (.A1(_12344_),
    .A2(_12347_),
    .B1(_12350_),
    .Y(_12351_));
 sky130_fd_sc_hd__nand3_2 _33993_ (.A(_12344_),
    .B(_12350_),
    .C(_12347_),
    .Y(_12352_));
 sky130_fd_sc_hd__and2b_2 _33994_ (.A_N(_12351_),
    .B(_12352_),
    .X(_12353_));
 sky130_fd_sc_hd__a21oi_2 _33995_ (.A1(_12283_),
    .A2(_12287_),
    .B1(_12353_),
    .Y(_12354_));
 sky130_fd_sc_hd__a21o_2 _33996_ (.A1(_12344_),
    .A2(_12347_),
    .B1(_12350_),
    .X(_12355_));
 sky130_fd_sc_hd__nand2_2 _33997_ (.A(_12355_),
    .B(_12352_),
    .Y(_12356_));
 sky130_fd_sc_hd__a21oi_2 _33998_ (.A1(_12284_),
    .A2(_12285_),
    .B1(_12282_),
    .Y(_12357_));
 sky130_vsdinv _33999_ (.A(_12287_),
    .Y(_12358_));
 sky130_fd_sc_hd__nor3_2 _34000_ (.A(_12356_),
    .B(_12357_),
    .C(_12358_),
    .Y(_12359_));
 sky130_fd_sc_hd__o21ai_2 _34001_ (.A1(_12056_),
    .A2(_12058_),
    .B1(_11998_),
    .Y(_12360_));
 sky130_fd_sc_hd__o21bai_2 _34002_ (.A1(_12354_),
    .A2(_12359_),
    .B1_N(_12360_),
    .Y(_12361_));
 sky130_fd_sc_hd__nand2_2 _34003_ (.A(_12283_),
    .B(_12286_),
    .Y(_12362_));
 sky130_fd_sc_hd__nand2_2 _34004_ (.A(_12362_),
    .B(_12356_),
    .Y(_12363_));
 sky130_fd_sc_hd__nand3_2 _34005_ (.A(_12353_),
    .B(_12287_),
    .C(_12283_),
    .Y(_12364_));
 sky130_fd_sc_hd__nand3_2 _34006_ (.A(_12363_),
    .B(_12364_),
    .C(_12360_),
    .Y(_12365_));
 sky130_fd_sc_hd__o21a_2 _34007_ (.A1(_05634_),
    .A2(_08291_),
    .B1(_11203_),
    .X(_12366_));
 sky130_fd_sc_hd__buf_1 _34008_ (.A(_12366_),
    .X(_12367_));
 sky130_fd_sc_hd__buf_1 _34009_ (.A(_16961_),
    .X(_12368_));
 sky130_fd_sc_hd__nand3_2 _34010_ (.A(_12368_),
    .B(_07595_),
    .C(_05504_),
    .Y(_12369_));
 sky130_fd_sc_hd__a21boi_2 _34011_ (.A1(_12367_),
    .A2(_12369_),
    .B1_N(_11188_),
    .Y(_12370_));
 sky130_fd_sc_hd__o211a_2 _34012_ (.A1(_11487_),
    .A2(_18880_),
    .B1(_12369_),
    .C1(_12366_),
    .X(_12371_));
 sky130_fd_sc_hd__o221ai_2 _34013_ (.A1(_12098_),
    .A2(_12100_),
    .B1(_12370_),
    .B2(_12371_),
    .C1(_12102_),
    .Y(_12372_));
 sky130_fd_sc_hd__nor2_2 _34014_ (.A(_12098_),
    .B(_12100_),
    .Y(_12373_));
 sky130_fd_sc_hd__nor2_2 _34015_ (.A(_10888_),
    .B(_12103_),
    .Y(_12374_));
 sky130_fd_sc_hd__nor2_2 _34016_ (.A(_12370_),
    .B(_12371_),
    .Y(_12375_));
 sky130_fd_sc_hd__o21ai_2 _34017_ (.A1(_12373_),
    .A2(_12374_),
    .B1(_12375_),
    .Y(_12376_));
 sky130_fd_sc_hd__o211a_2 _34018_ (.A1(_11832_),
    .A2(_11833_),
    .B1(_12372_),
    .C1(_12376_),
    .X(_12377_));
 sky130_fd_sc_hd__a21boi_2 _34019_ (.A1(_12108_),
    .A2(_12110_),
    .B1_N(_12109_),
    .Y(_12378_));
 sky130_vsdinv _34020_ (.A(_12378_),
    .Y(_12379_));
 sky130_fd_sc_hd__a21boi_2 _34021_ (.A1(_12376_),
    .A2(_12372_),
    .B1_N(_11835_),
    .Y(_12380_));
 sky130_vsdinv _34022_ (.A(_12380_),
    .Y(_12381_));
 sky130_fd_sc_hd__nand3b_2 _34023_ (.A_N(_12377_),
    .B(_12379_),
    .C(_12381_),
    .Y(_12382_));
 sky130_fd_sc_hd__o21ai_2 _34024_ (.A1(_12380_),
    .A2(_12377_),
    .B1(_12378_),
    .Y(_12383_));
 sky130_fd_sc_hd__nand3_2 _34025_ (.A(_12382_),
    .B(_12118_),
    .C(_12383_),
    .Y(_12384_));
 sky130_fd_sc_hd__a21o_2 _34026_ (.A1(_12382_),
    .A2(_12383_),
    .B1(_12118_),
    .X(_12385_));
 sky130_fd_sc_hd__a22o_2 _34027_ (.A1(_06311_),
    .A2(_12069_),
    .B1(_18834_),
    .B2(_10913_),
    .X(_12386_));
 sky130_fd_sc_hd__nand2_2 _34028_ (.A(_06890_),
    .B(_19139_),
    .Y(_12387_));
 sky130_fd_sc_hd__nand3b_2 _34029_ (.A_N(_12387_),
    .B(_18830_),
    .C(_10895_),
    .Y(_12388_));
 sky130_fd_sc_hd__buf_1 _34030_ (.A(_10541_),
    .X(_12389_));
 sky130_fd_sc_hd__o2bb2ai_2 _34031_ (.A1_N(_12386_),
    .A2_N(_12388_),
    .B1(_06114_),
    .B2(_12389_),
    .Y(_12390_));
 sky130_fd_sc_hd__and2_2 _34032_ (.A(_05779_),
    .B(_11201_),
    .X(_12391_));
 sky130_fd_sc_hd__nand3_2 _34033_ (.A(_12388_),
    .B(_12386_),
    .C(_12391_),
    .Y(_12392_));
 sky130_fd_sc_hd__nand2_2 _34034_ (.A(_12037_),
    .B(_12038_),
    .Y(_12393_));
 sky130_fd_sc_hd__nor2_2 _34035_ (.A(_12037_),
    .B(_12038_),
    .Y(_12394_));
 sky130_fd_sc_hd__a21oi_2 _34036_ (.A1(_12393_),
    .A2(_12036_),
    .B1(_12394_),
    .Y(_12395_));
 sky130_vsdinv _34037_ (.A(_12395_),
    .Y(_12396_));
 sky130_fd_sc_hd__a21o_2 _34038_ (.A1(_12390_),
    .A2(_12392_),
    .B1(_12396_),
    .X(_12397_));
 sky130_fd_sc_hd__nand3_2 _34039_ (.A(_12390_),
    .B(_12396_),
    .C(_12392_),
    .Y(_12398_));
 sky130_fd_sc_hd__a21boi_2 _34040_ (.A1(_12067_),
    .A2(_12072_),
    .B1_N(_12070_),
    .Y(_12399_));
 sky130_vsdinv _34041_ (.A(_12399_),
    .Y(_12400_));
 sky130_fd_sc_hd__a21oi_2 _34042_ (.A1(_12397_),
    .A2(_12398_),
    .B1(_12400_),
    .Y(_12401_));
 sky130_fd_sc_hd__nand3_2 _34043_ (.A(_12397_),
    .B(_12400_),
    .C(_12398_),
    .Y(_12402_));
 sky130_vsdinv _34044_ (.A(_12402_),
    .Y(_12403_));
 sky130_fd_sc_hd__o21ai_2 _34045_ (.A1(_12031_),
    .A2(_12040_),
    .B1(_12033_),
    .Y(_12404_));
 sky130_fd_sc_hd__o21bai_2 _34046_ (.A1(_12401_),
    .A2(_12403_),
    .B1_N(_12404_),
    .Y(_12405_));
 sky130_fd_sc_hd__a21o_2 _34047_ (.A1(_12397_),
    .A2(_12398_),
    .B1(_12400_),
    .X(_12406_));
 sky130_fd_sc_hd__nand3_2 _34048_ (.A(_12406_),
    .B(_12404_),
    .C(_12402_),
    .Y(_12407_));
 sky130_fd_sc_hd__a21boi_2 _34049_ (.A1(_12077_),
    .A2(_12081_),
    .B1_N(_12079_),
    .Y(_12408_));
 sky130_vsdinv _34050_ (.A(_12408_),
    .Y(_12409_));
 sky130_fd_sc_hd__a21oi_2 _34051_ (.A1(_12405_),
    .A2(_12407_),
    .B1(_12409_),
    .Y(_12410_));
 sky130_fd_sc_hd__nand3_2 _34052_ (.A(_12405_),
    .B(_12409_),
    .C(_12407_),
    .Y(_12411_));
 sky130_vsdinv _34053_ (.A(_12411_),
    .Y(_12412_));
 sky130_fd_sc_hd__o21ai_2 _34054_ (.A1(_12088_),
    .A2(_12085_),
    .B1(_12086_),
    .Y(_12413_));
 sky130_fd_sc_hd__o21bai_2 _34055_ (.A1(_12410_),
    .A2(_12412_),
    .B1_N(_12413_),
    .Y(_12414_));
 sky130_fd_sc_hd__a21o_2 _34056_ (.A1(_12405_),
    .A2(_12407_),
    .B1(_12409_),
    .X(_12415_));
 sky130_fd_sc_hd__nand3_2 _34057_ (.A(_12415_),
    .B(_12411_),
    .C(_12413_),
    .Y(_12416_));
 sky130_fd_sc_hd__a22oi_2 _34058_ (.A1(_12384_),
    .A2(_12385_),
    .B1(_12414_),
    .B2(_12416_),
    .Y(_12417_));
 sky130_fd_sc_hd__nand2_2 _34059_ (.A(_12385_),
    .B(_12384_),
    .Y(_12418_));
 sky130_fd_sc_hd__nand2_2 _34060_ (.A(_12414_),
    .B(_12416_),
    .Y(_12419_));
 sky130_fd_sc_hd__nor2_2 _34061_ (.A(_12418_),
    .B(_12419_),
    .Y(_12420_));
 sky130_fd_sc_hd__a21oi_2 _34062_ (.A1(_12044_),
    .A2(_12045_),
    .B1(_12049_),
    .Y(_12421_));
 sky130_fd_sc_hd__o21ai_2 _34063_ (.A1(_12052_),
    .A2(_12421_),
    .B1(_12050_),
    .Y(_12422_));
 sky130_fd_sc_hd__o21bai_2 _34064_ (.A1(_12417_),
    .A2(_12420_),
    .B1_N(_12422_),
    .Y(_12423_));
 sky130_fd_sc_hd__nand3b_2 _34065_ (.A_N(_12418_),
    .B(_12414_),
    .C(_12416_),
    .Y(_12424_));
 sky130_fd_sc_hd__nand3b_2 _34066_ (.A_N(_12417_),
    .B(_12422_),
    .C(_12424_),
    .Y(_12425_));
 sky130_fd_sc_hd__nand2_2 _34067_ (.A(_12423_),
    .B(_12425_),
    .Y(_12426_));
 sky130_fd_sc_hd__a21boi_2 _34068_ (.A1(_12122_),
    .A2(_12094_),
    .B1_N(_12096_),
    .Y(_12427_));
 sky130_fd_sc_hd__nand2_2 _34069_ (.A(_12426_),
    .B(_12427_),
    .Y(_12428_));
 sky130_fd_sc_hd__nand3b_2 _34070_ (.A_N(_12427_),
    .B(_12423_),
    .C(_12425_),
    .Y(_12429_));
 sky130_fd_sc_hd__nand2_2 _34071_ (.A(_12428_),
    .B(_12429_),
    .Y(_12430_));
 sky130_fd_sc_hd__buf_1 _34072_ (.A(_12430_),
    .X(_12431_));
 sky130_fd_sc_hd__a21boi_2 _34073_ (.A1(_12361_),
    .A2(_12365_),
    .B1_N(_12431_),
    .Y(_12432_));
 sky130_fd_sc_hd__a21oi_2 _34074_ (.A1(_12363_),
    .A2(_12364_),
    .B1(_12360_),
    .Y(_12433_));
 sky130_vsdinv _34075_ (.A(_12365_),
    .Y(_12434_));
 sky130_fd_sc_hd__nor3_2 _34076_ (.A(_12431_),
    .B(_12433_),
    .C(_12434_),
    .Y(_12435_));
 sky130_fd_sc_hd__o21ai_2 _34077_ (.A1(_12140_),
    .A2(_12141_),
    .B1(_12066_),
    .Y(_12436_));
 sky130_fd_sc_hd__o21bai_2 _34078_ (.A1(_12432_),
    .A2(_12435_),
    .B1_N(_12436_),
    .Y(_12437_));
 sky130_fd_sc_hd__o21ai_2 _34079_ (.A1(_12433_),
    .A2(_12434_),
    .B1(_12431_),
    .Y(_12438_));
 sky130_fd_sc_hd__nand3b_2 _34080_ (.A_N(_12430_),
    .B(_12365_),
    .C(_12361_),
    .Y(_12439_));
 sky130_fd_sc_hd__nand3_2 _34081_ (.A(_12438_),
    .B(_12439_),
    .C(_12436_),
    .Y(_12440_));
 sky130_fd_sc_hd__buf_1 _34082_ (.A(_12440_),
    .X(_12441_));
 sky130_fd_sc_hd__buf_1 _34083_ (.A(_12117_),
    .X(_12442_));
 sky130_fd_sc_hd__a21boi_2 _34084_ (.A1(_12114_),
    .A2(_12442_),
    .B1_N(_12115_),
    .Y(_12443_));
 sky130_fd_sc_hd__nand2_2 _34085_ (.A(_12139_),
    .B(_12131_),
    .Y(_12444_));
 sky130_fd_sc_hd__xnor2_2 _34086_ (.A(_12443_),
    .B(_12444_),
    .Y(_12445_));
 sky130_fd_sc_hd__a21oi_2 _34087_ (.A1(_12437_),
    .A2(_12441_),
    .B1(_12445_),
    .Y(_12446_));
 sky130_fd_sc_hd__nand3_2 _34088_ (.A(_12437_),
    .B(_12445_),
    .C(_12440_),
    .Y(_12447_));
 sky130_vsdinv _34089_ (.A(_12447_),
    .Y(_12448_));
 sky130_fd_sc_hd__o21ai_2 _34090_ (.A1(_12154_),
    .A2(_12155_),
    .B1(_12149_),
    .Y(_12449_));
 sky130_fd_sc_hd__o21bai_2 _34091_ (.A1(_12446_),
    .A2(_12448_),
    .B1_N(_12449_),
    .Y(_12450_));
 sky130_fd_sc_hd__nand2_2 _34092_ (.A(_12437_),
    .B(_12441_),
    .Y(_12451_));
 sky130_vsdinv _34093_ (.A(_12445_),
    .Y(_12452_));
 sky130_fd_sc_hd__nand2_2 _34094_ (.A(_12451_),
    .B(_12452_),
    .Y(_12453_));
 sky130_fd_sc_hd__nand3_2 _34095_ (.A(_12453_),
    .B(_12447_),
    .C(_12449_),
    .Y(_12454_));
 sky130_fd_sc_hd__a21oi_2 _34096_ (.A1(_11860_),
    .A2(_11856_),
    .B1(_12150_),
    .Y(_12455_));
 sky130_fd_sc_hd__a21oi_2 _34097_ (.A1(_12450_),
    .A2(_12454_),
    .B1(_12455_),
    .Y(_12456_));
 sky130_fd_sc_hd__nand3_2 _34098_ (.A(_12450_),
    .B(_12455_),
    .C(_12454_),
    .Y(_12457_));
 sky130_vsdinv _34099_ (.A(_12457_),
    .Y(_12458_));
 sky130_fd_sc_hd__o21ai_2 _34100_ (.A1(_12165_),
    .A2(_12166_),
    .B1(_12162_),
    .Y(_12459_));
 sky130_fd_sc_hd__o21bai_2 _34101_ (.A1(_12456_),
    .A2(_12458_),
    .B1_N(_12459_),
    .Y(_12460_));
 sky130_fd_sc_hd__a21o_2 _34102_ (.A1(_12450_),
    .A2(_12454_),
    .B1(_12455_),
    .X(_12461_));
 sky130_fd_sc_hd__nand3_2 _34103_ (.A(_12461_),
    .B(_12459_),
    .C(_12457_),
    .Y(_12462_));
 sky130_fd_sc_hd__nand2_2 _34104_ (.A(_12460_),
    .B(_12462_),
    .Y(_12463_));
 sky130_fd_sc_hd__o21ai_2 _34105_ (.A1(_12176_),
    .A2(_12182_),
    .B1(_12175_),
    .Y(_12464_));
 sky130_fd_sc_hd__xnor2_2 _34106_ (.A(_12463_),
    .B(_12464_),
    .Y(_02656_));
 sky130_fd_sc_hd__and2b_2 _34107_ (.A_N(_05671_),
    .B(_12183_),
    .X(_12465_));
 sky130_fd_sc_hd__and2_2 _34108_ (.A(_10669_),
    .B(_06043_),
    .X(_12466_));
 sky130_fd_sc_hd__nand2_2 _34109_ (.A(_12465_),
    .B(_12466_),
    .Y(_12467_));
 sky130_fd_sc_hd__nand2_2 _34110_ (.A(_10994_),
    .B(_05649_),
    .Y(_12468_));
 sky130_fd_sc_hd__o21ai_2 _34111_ (.A1(_06041_),
    .A2(_11331_),
    .B1(_12468_),
    .Y(_12469_));
 sky130_fd_sc_hd__and2_2 _34112_ (.A(_11326_),
    .B(_07499_),
    .X(_12470_));
 sky130_fd_sc_hd__a21oi_2 _34113_ (.A1(_12467_),
    .A2(_12469_),
    .B1(_12470_),
    .Y(_12471_));
 sky130_fd_sc_hd__nand3_2 _34114_ (.A(_12467_),
    .B(_12469_),
    .C(_12470_),
    .Y(_12472_));
 sky130_vsdinv _34115_ (.A(_12472_),
    .Y(_12473_));
 sky130_fd_sc_hd__a21oi_2 _34116_ (.A1(_12190_),
    .A2(_12187_),
    .B1(_12186_),
    .Y(_12474_));
 sky130_fd_sc_hd__o21ai_2 _34117_ (.A1(_12471_),
    .A2(_12473_),
    .B1(_12474_),
    .Y(_12475_));
 sky130_fd_sc_hd__a21o_2 _34118_ (.A1(_12187_),
    .A2(_12190_),
    .B1(_12186_),
    .X(_12476_));
 sky130_fd_sc_hd__buf_1 _34119_ (.A(_10487_),
    .X(_12477_));
 sky130_fd_sc_hd__a22oi_2 _34120_ (.A1(_12477_),
    .A2(_06486_),
    .B1(_19274_),
    .B2(_11289_),
    .Y(_12478_));
 sky130_fd_sc_hd__nor3_2 _34121_ (.A(_05671_),
    .B(_10675_),
    .C(_12468_),
    .Y(_12479_));
 sky130_fd_sc_hd__o21bai_2 _34122_ (.A1(_12478_),
    .A2(_12479_),
    .B1_N(_12470_),
    .Y(_12480_));
 sky130_fd_sc_hd__nand3_2 _34123_ (.A(_12476_),
    .B(_12480_),
    .C(_12472_),
    .Y(_12481_));
 sky130_fd_sc_hd__a22oi_2 _34124_ (.A1(_11618_),
    .A2(_05950_),
    .B1(_11340_),
    .B2(_06883_),
    .Y(_12482_));
 sky130_fd_sc_hd__and4_2 _34125_ (.A(_10683_),
    .B(_11340_),
    .C(_05935_),
    .D(_08035_),
    .X(_12483_));
 sky130_fd_sc_hd__and2_2 _34126_ (.A(_10474_),
    .B(_07060_),
    .X(_12484_));
 sky130_fd_sc_hd__o21bai_2 _34127_ (.A1(_12482_),
    .A2(_12483_),
    .B1_N(_12484_),
    .Y(_12485_));
 sky130_fd_sc_hd__nand2_2 _34128_ (.A(_11338_),
    .B(_05950_),
    .Y(_12486_));
 sky130_fd_sc_hd__nand3b_2 _34129_ (.A_N(_12486_),
    .B(_10263_),
    .C(_06444_),
    .Y(_12487_));
 sky130_fd_sc_hd__nand3b_2 _34130_ (.A_N(_12482_),
    .B(_12487_),
    .C(_12484_),
    .Y(_12488_));
 sky130_fd_sc_hd__nand2_2 _34131_ (.A(_12485_),
    .B(_12488_),
    .Y(_12489_));
 sky130_vsdinv _34132_ (.A(_12489_),
    .Y(_12490_));
 sky130_fd_sc_hd__a21oi_2 _34133_ (.A1(_12475_),
    .A2(_12481_),
    .B1(_12490_),
    .Y(_12491_));
 sky130_fd_sc_hd__a21oi_2 _34134_ (.A1(_12480_),
    .A2(_12472_),
    .B1(_12476_),
    .Y(_12492_));
 sky130_fd_sc_hd__nor3_2 _34135_ (.A(_12474_),
    .B(_12471_),
    .C(_12473_),
    .Y(_12493_));
 sky130_fd_sc_hd__nor3_2 _34136_ (.A(_12489_),
    .B(_12492_),
    .C(_12493_),
    .Y(_12494_));
 sky130_fd_sc_hd__o21ai_2 _34137_ (.A1(_12203_),
    .A2(_12206_),
    .B1(_12195_),
    .Y(_12495_));
 sky130_fd_sc_hd__o21bai_2 _34138_ (.A1(_12491_),
    .A2(_12494_),
    .B1_N(_12495_),
    .Y(_12496_));
 sky130_fd_sc_hd__o21bai_2 _34139_ (.A1(_12492_),
    .A2(_12493_),
    .B1_N(_12490_),
    .Y(_12497_));
 sky130_fd_sc_hd__nand3_2 _34140_ (.A(_12475_),
    .B(_12490_),
    .C(_12481_),
    .Y(_12498_));
 sky130_fd_sc_hd__nand3_2 _34141_ (.A(_12497_),
    .B(_12495_),
    .C(_12498_),
    .Y(_12499_));
 sky130_fd_sc_hd__buf_1 _34142_ (.A(_10229_),
    .X(_12500_));
 sky130_fd_sc_hd__a22o_2 _34143_ (.A1(_12500_),
    .A2(_06464_),
    .B1(_12217_),
    .B2(_06467_),
    .X(_12501_));
 sky130_fd_sc_hd__nand2_2 _34144_ (.A(_11636_),
    .B(_08054_),
    .Y(_12502_));
 sky130_fd_sc_hd__nand3b_2 _34145_ (.A_N(_12502_),
    .B(_12500_),
    .C(_06366_),
    .Y(_12503_));
 sky130_fd_sc_hd__o2bb2ai_2 _34146_ (.A1_N(_12501_),
    .A2_N(_12503_),
    .B1(_10246_),
    .B2(_19233_),
    .Y(_12504_));
 sky130_fd_sc_hd__and2_2 _34147_ (.A(_08759_),
    .B(_10743_),
    .X(_12505_));
 sky130_fd_sc_hd__nand3_2 _34148_ (.A(_12503_),
    .B(_12501_),
    .C(_12505_),
    .Y(_12506_));
 sky130_fd_sc_hd__o31ai_2 _34149_ (.A1(_18725_),
    .A2(_19254_),
    .A3(_12196_),
    .B1(_12201_),
    .Y(_12507_));
 sky130_fd_sc_hd__a21o_2 _34150_ (.A1(_12504_),
    .A2(_12506_),
    .B1(_12507_),
    .X(_12508_));
 sky130_fd_sc_hd__nand3_2 _34151_ (.A(_12507_),
    .B(_12504_),
    .C(_12506_),
    .Y(_12509_));
 sky130_fd_sc_hd__a21boi_2 _34152_ (.A1(_12221_),
    .A2(_12215_),
    .B1_N(_12218_),
    .Y(_12510_));
 sky130_vsdinv _34153_ (.A(_12510_),
    .Y(_12511_));
 sky130_fd_sc_hd__a21o_2 _34154_ (.A1(_12508_),
    .A2(_12509_),
    .B1(_12511_),
    .X(_12512_));
 sky130_fd_sc_hd__nand3_2 _34155_ (.A(_12508_),
    .B(_12511_),
    .C(_12509_),
    .Y(_12513_));
 sky130_fd_sc_hd__nand2_2 _34156_ (.A(_12512_),
    .B(_12513_),
    .Y(_12514_));
 sky130_fd_sc_hd__buf_1 _34157_ (.A(_12514_),
    .X(_12515_));
 sky130_fd_sc_hd__a21boi_2 _34158_ (.A1(_12496_),
    .A2(_12499_),
    .B1_N(_12515_),
    .Y(_12516_));
 sky130_fd_sc_hd__a21oi_2 _34159_ (.A1(_12497_),
    .A2(_12498_),
    .B1(_12495_),
    .Y(_12517_));
 sky130_vsdinv _34160_ (.A(_12499_),
    .Y(_12518_));
 sky130_fd_sc_hd__nor3_2 _34161_ (.A(_12515_),
    .B(_12517_),
    .C(_12518_),
    .Y(_12519_));
 sky130_fd_sc_hd__o21ai_2 _34162_ (.A1(_12232_),
    .A2(_12234_),
    .B1(_12214_),
    .Y(_12520_));
 sky130_fd_sc_hd__o21bai_2 _34163_ (.A1(_12516_),
    .A2(_12519_),
    .B1_N(_12520_),
    .Y(_12521_));
 sky130_fd_sc_hd__o21ai_2 _34164_ (.A1(_12517_),
    .A2(_12518_),
    .B1(_12515_),
    .Y(_12522_));
 sky130_fd_sc_hd__nand3b_2 _34165_ (.A_N(_12514_),
    .B(_12499_),
    .C(_12496_),
    .Y(_12523_));
 sky130_fd_sc_hd__nand3_2 _34166_ (.A(_12522_),
    .B(_12520_),
    .C(_12523_),
    .Y(_12524_));
 sky130_fd_sc_hd__buf_1 _34167_ (.A(_12524_),
    .X(_12525_));
 sky130_fd_sc_hd__a22o_2 _34168_ (.A1(_18749_),
    .A2(_07913_),
    .B1(_18754_),
    .B2(_07329_),
    .X(_12526_));
 sky130_fd_sc_hd__buf_1 _34169_ (.A(_08463_),
    .X(_12527_));
 sky130_fd_sc_hd__nand2_2 _34170_ (.A(_12527_),
    .B(_07906_),
    .Y(_12528_));
 sky130_fd_sc_hd__nand3b_2 _34171_ (.A_N(_12528_),
    .B(_10734_),
    .C(_10775_),
    .Y(_12529_));
 sky130_fd_sc_hd__o2bb2ai_2 _34172_ (.A1_N(_12526_),
    .A2_N(_12529_),
    .B1(_10736_),
    .B2(_19213_),
    .Y(_12530_));
 sky130_fd_sc_hd__buf_1 _34173_ (.A(_11080_),
    .X(_12531_));
 sky130_fd_sc_hd__and2_2 _34174_ (.A(_12531_),
    .B(_07606_),
    .X(_12532_));
 sky130_fd_sc_hd__nand3_2 _34175_ (.A(_12529_),
    .B(_12526_),
    .C(_12532_),
    .Y(_12533_));
 sky130_fd_sc_hd__a21oi_2 _34176_ (.A1(_12246_),
    .A2(_12245_),
    .B1(_12244_),
    .Y(_12534_));
 sky130_vsdinv _34177_ (.A(_12534_),
    .Y(_12535_));
 sky130_fd_sc_hd__a21o_2 _34178_ (.A1(_12530_),
    .A2(_12533_),
    .B1(_12535_),
    .X(_12536_));
 sky130_fd_sc_hd__nand3_2 _34179_ (.A(_12530_),
    .B(_12535_),
    .C(_12533_),
    .Y(_12537_));
 sky130_fd_sc_hd__buf_1 _34180_ (.A(_10436_),
    .X(_12538_));
 sky130_fd_sc_hd__and2_2 _34181_ (.A(_12538_),
    .B(_08314_),
    .X(_12539_));
 sky130_fd_sc_hd__buf_1 _34182_ (.A(_07537_),
    .X(_12540_));
 sky130_fd_sc_hd__nand2_2 _34183_ (.A(_12540_),
    .B(_10376_),
    .Y(_12541_));
 sky130_fd_sc_hd__nand2_2 _34184_ (.A(_11067_),
    .B(_08292_),
    .Y(_12542_));
 sky130_fd_sc_hd__xnor2_2 _34185_ (.A(_12541_),
    .B(_12542_),
    .Y(_12543_));
 sky130_fd_sc_hd__xnor2_2 _34186_ (.A(_12539_),
    .B(_12543_),
    .Y(_12544_));
 sky130_fd_sc_hd__a21oi_2 _34187_ (.A1(_12536_),
    .A2(_12537_),
    .B1(_12544_),
    .Y(_12545_));
 sky130_fd_sc_hd__nand3_2 _34188_ (.A(_12544_),
    .B(_12536_),
    .C(_12537_),
    .Y(_12546_));
 sky130_vsdinv _34189_ (.A(_12546_),
    .Y(_12547_));
 sky130_fd_sc_hd__nand2_2 _34190_ (.A(_12230_),
    .B(_12226_),
    .Y(_12548_));
 sky130_fd_sc_hd__o21bai_2 _34191_ (.A1(_12545_),
    .A2(_12547_),
    .B1_N(_12548_),
    .Y(_12549_));
 sky130_fd_sc_hd__a21o_2 _34192_ (.A1(_12536_),
    .A2(_12537_),
    .B1(_12544_),
    .X(_12550_));
 sky130_fd_sc_hd__nand3_2 _34193_ (.A(_12548_),
    .B(_12550_),
    .C(_12546_),
    .Y(_12551_));
 sky130_fd_sc_hd__a31oi_2 _34194_ (.A1(_12251_),
    .A2(_12261_),
    .A3(_12259_),
    .B1(_12264_),
    .Y(_12552_));
 sky130_vsdinv _34195_ (.A(_12552_),
    .Y(_12553_));
 sky130_fd_sc_hd__a21oi_2 _34196_ (.A1(_12549_),
    .A2(_12551_),
    .B1(_12553_),
    .Y(_12554_));
 sky130_fd_sc_hd__nand3_2 _34197_ (.A(_12549_),
    .B(_12553_),
    .C(_12551_),
    .Y(_12555_));
 sky130_vsdinv _34198_ (.A(_12555_),
    .Y(_12556_));
 sky130_fd_sc_hd__nor2_2 _34199_ (.A(_12554_),
    .B(_12556_),
    .Y(_12557_));
 sky130_fd_sc_hd__a21oi_2 _34200_ (.A1(_12521_),
    .A2(_12525_),
    .B1(_12557_),
    .Y(_12558_));
 sky130_fd_sc_hd__nand2_2 _34201_ (.A(_12549_),
    .B(_12551_),
    .Y(_12559_));
 sky130_fd_sc_hd__nand2_2 _34202_ (.A(_12559_),
    .B(_12552_),
    .Y(_12560_));
 sky130_fd_sc_hd__nand2_2 _34203_ (.A(_12560_),
    .B(_12555_),
    .Y(_12561_));
 sky130_fd_sc_hd__a21oi_2 _34204_ (.A1(_12522_),
    .A2(_12523_),
    .B1(_12520_),
    .Y(_12562_));
 sky130_vsdinv _34205_ (.A(_12525_),
    .Y(_12563_));
 sky130_fd_sc_hd__nor3_2 _34206_ (.A(_12561_),
    .B(_12562_),
    .C(_12563_),
    .Y(_12564_));
 sky130_fd_sc_hd__o21ai_2 _34207_ (.A1(_12278_),
    .A2(_12279_),
    .B1(_12241_),
    .Y(_12565_));
 sky130_fd_sc_hd__o21bai_2 _34208_ (.A1(_12558_),
    .A2(_12564_),
    .B1_N(_12565_),
    .Y(_12566_));
 sky130_fd_sc_hd__o2bb2ai_2 _34209_ (.A1_N(_12525_),
    .A2_N(_12521_),
    .B1(_12556_),
    .B2(_12554_),
    .Y(_12567_));
 sky130_fd_sc_hd__nand3_2 _34210_ (.A(_12557_),
    .B(_12525_),
    .C(_12521_),
    .Y(_12568_));
 sky130_fd_sc_hd__nand3_2 _34211_ (.A(_12567_),
    .B(_12565_),
    .C(_12568_),
    .Y(_12569_));
 sky130_fd_sc_hd__nand2_2 _34212_ (.A(_12566_),
    .B(_12569_),
    .Y(_12570_));
 sky130_fd_sc_hd__a22o_2 _34213_ (.A1(_10777_),
    .A2(_08310_),
    .B1(_18786_),
    .B2(_12295_),
    .X(_12571_));
 sky130_fd_sc_hd__nand2_2 _34214_ (.A(_07480_),
    .B(_09755_),
    .Y(_12572_));
 sky130_fd_sc_hd__nand3b_2 _34215_ (.A_N(_12572_),
    .B(_18781_),
    .C(_12292_),
    .Y(_12573_));
 sky130_fd_sc_hd__o2bb2ai_2 _34216_ (.A1_N(_12571_),
    .A2_N(_12573_),
    .B1(_11716_),
    .B2(_19182_),
    .Y(_12574_));
 sky130_fd_sc_hd__and2_2 _34217_ (.A(_11409_),
    .B(_10077_),
    .X(_12575_));
 sky130_fd_sc_hd__nand3_2 _34218_ (.A(_12573_),
    .B(_12571_),
    .C(_12575_),
    .Y(_12576_));
 sky130_fd_sc_hd__a21oi_2 _34219_ (.A1(_12256_),
    .A2(_12260_),
    .B1(_12257_),
    .Y(_12577_));
 sky130_fd_sc_hd__a21bo_2 _34220_ (.A1(_12574_),
    .A2(_12576_),
    .B1_N(_12577_),
    .X(_12578_));
 sky130_fd_sc_hd__nand3b_2 _34221_ (.A_N(_12577_),
    .B(_12574_),
    .C(_12576_),
    .Y(_12579_));
 sky130_fd_sc_hd__a21boi_2 _34222_ (.A1(_12290_),
    .A2(_12296_),
    .B1_N(_12293_),
    .Y(_12580_));
 sky130_vsdinv _34223_ (.A(_12580_),
    .Y(_12581_));
 sky130_fd_sc_hd__a21oi_2 _34224_ (.A1(_12578_),
    .A2(_12579_),
    .B1(_12581_),
    .Y(_12582_));
 sky130_fd_sc_hd__nand3_2 _34225_ (.A(_12578_),
    .B(_12581_),
    .C(_12579_),
    .Y(_12583_));
 sky130_fd_sc_hd__o21ai_2 _34226_ (.A1(_12305_),
    .A2(_12308_),
    .B1(_12304_),
    .Y(_12584_));
 sky130_fd_sc_hd__nand3b_2 _34227_ (.A_N(_12582_),
    .B(_12583_),
    .C(_12584_),
    .Y(_12585_));
 sky130_vsdinv _34228_ (.A(_12583_),
    .Y(_12586_));
 sky130_fd_sc_hd__o21bai_2 _34229_ (.A1(_12582_),
    .A2(_12586_),
    .B1_N(_12584_),
    .Y(_12587_));
 sky130_fd_sc_hd__and2_2 _34230_ (.A(_06680_),
    .B(_09793_),
    .X(_12588_));
 sky130_fd_sc_hd__nand2_2 _34231_ (.A(_06811_),
    .B(_10535_),
    .Y(_12589_));
 sky130_fd_sc_hd__nand2_2 _34232_ (.A(_11432_),
    .B(_09805_),
    .Y(_12590_));
 sky130_fd_sc_hd__xnor2_2 _34233_ (.A(_12589_),
    .B(_12590_),
    .Y(_12591_));
 sky130_fd_sc_hd__xor2_2 _34234_ (.A(_12588_),
    .B(_12591_),
    .X(_12592_));
 sky130_fd_sc_hd__nand2_2 _34235_ (.A(_06544_),
    .B(_08832_),
    .Y(_12593_));
 sky130_fd_sc_hd__nand2_2 _34236_ (.A(_18802_),
    .B(_08818_),
    .Y(_12594_));
 sky130_fd_sc_hd__xor2_2 _34237_ (.A(_12593_),
    .B(_12594_),
    .X(_12595_));
 sky130_fd_sc_hd__buf_1 _34238_ (.A(_19162_),
    .X(_12596_));
 sky130_fd_sc_hd__nand3_2 _34239_ (.A(_12595_),
    .B(_06276_),
    .C(_12596_),
    .Y(_12597_));
 sky130_fd_sc_hd__buf_1 _34240_ (.A(_12597_),
    .X(_12598_));
 sky130_fd_sc_hd__xnor2_2 _34241_ (.A(_12593_),
    .B(_12594_),
    .Y(_12599_));
 sky130_fd_sc_hd__o21ai_2 _34242_ (.A1(_18811_),
    .A2(_19164_),
    .B1(_12599_),
    .Y(_12600_));
 sky130_fd_sc_hd__a21oi_2 _34243_ (.A1(_12327_),
    .A2(_12326_),
    .B1(_12324_),
    .Y(_12601_));
 sky130_vsdinv _34244_ (.A(_12601_),
    .Y(_12602_));
 sky130_fd_sc_hd__a21oi_2 _34245_ (.A1(_12598_),
    .A2(_12600_),
    .B1(_12602_),
    .Y(_12603_));
 sky130_fd_sc_hd__nand3_2 _34246_ (.A(_12598_),
    .B(_12600_),
    .C(_12602_),
    .Y(_12604_));
 sky130_fd_sc_hd__nor3b_2 _34247_ (.A(_12592_),
    .B(_12603_),
    .C_N(_12604_),
    .Y(_12605_));
 sky130_fd_sc_hd__a21o_2 _34248_ (.A1(_12598_),
    .A2(_12600_),
    .B1(_12602_),
    .X(_12606_));
 sky130_fd_sc_hd__a21boi_2 _34249_ (.A1(_12606_),
    .A2(_12604_),
    .B1_N(_12592_),
    .Y(_12607_));
 sky130_fd_sc_hd__o2bb2ai_2 _34250_ (.A1_N(_12585_),
    .A2_N(_12587_),
    .B1(_12605_),
    .B2(_12607_),
    .Y(_12608_));
 sky130_fd_sc_hd__nor2_2 _34251_ (.A(_12607_),
    .B(_12605_),
    .Y(_12609_));
 sky130_fd_sc_hd__nand3_2 _34252_ (.A(_12587_),
    .B(_12609_),
    .C(_12585_),
    .Y(_12610_));
 sky130_fd_sc_hd__nand2_2 _34253_ (.A(_12273_),
    .B(_12269_),
    .Y(_12611_));
 sky130_fd_sc_hd__a21oi_2 _34254_ (.A1(_12608_),
    .A2(_12610_),
    .B1(_12611_),
    .Y(_12612_));
 sky130_fd_sc_hd__nand3_2 _34255_ (.A(_12608_),
    .B(_12611_),
    .C(_12610_),
    .Y(_12613_));
 sky130_vsdinv _34256_ (.A(_12613_),
    .Y(_12614_));
 sky130_fd_sc_hd__a21boi_2 _34257_ (.A1(_12337_),
    .A2(_12312_),
    .B1_N(_12315_),
    .Y(_12615_));
 sky130_vsdinv _34258_ (.A(_12615_),
    .Y(_12616_));
 sky130_fd_sc_hd__o21bai_2 _34259_ (.A1(_12612_),
    .A2(_12614_),
    .B1_N(_12616_),
    .Y(_12617_));
 sky130_fd_sc_hd__a21o_2 _34260_ (.A1(_12608_),
    .A2(_12610_),
    .B1(_12611_),
    .X(_12618_));
 sky130_fd_sc_hd__nand3_2 _34261_ (.A(_12618_),
    .B(_12616_),
    .C(_12613_),
    .Y(_12619_));
 sky130_fd_sc_hd__nand2_2 _34262_ (.A(_12617_),
    .B(_12619_),
    .Y(_12620_));
 sky130_fd_sc_hd__nand2_2 _34263_ (.A(_12570_),
    .B(_12620_),
    .Y(_12621_));
 sky130_fd_sc_hd__a21oi_2 _34264_ (.A1(_12618_),
    .A2(_12613_),
    .B1(_12616_),
    .Y(_12622_));
 sky130_vsdinv _34265_ (.A(_12619_),
    .Y(_12623_));
 sky130_fd_sc_hd__nor2_2 _34266_ (.A(_12622_),
    .B(_12623_),
    .Y(_12624_));
 sky130_fd_sc_hd__nand3_2 _34267_ (.A(_12624_),
    .B(_12566_),
    .C(_12569_),
    .Y(_12625_));
 sky130_fd_sc_hd__nand2_2 _34268_ (.A(_12621_),
    .B(_12625_),
    .Y(_12626_));
 sky130_fd_sc_hd__a21oi_2 _34269_ (.A1(_12353_),
    .A2(_12283_),
    .B1(_12358_),
    .Y(_12627_));
 sky130_fd_sc_hd__nand2_2 _34270_ (.A(_12626_),
    .B(_12627_),
    .Y(_12628_));
 sky130_fd_sc_hd__o21ai_2 _34271_ (.A1(_12356_),
    .A2(_12357_),
    .B1(_12287_),
    .Y(_12629_));
 sky130_fd_sc_hd__nand3_2 _34272_ (.A(_12621_),
    .B(_12629_),
    .C(_12625_),
    .Y(_12630_));
 sky130_fd_sc_hd__buf_1 _34273_ (.A(_12630_),
    .X(_12631_));
 sky130_fd_sc_hd__a22o_2 _34274_ (.A1(_05773_),
    .A2(_10897_),
    .B1(_06231_),
    .B2(_11201_),
    .X(_12632_));
 sky130_fd_sc_hd__nand2_2 _34275_ (.A(_05873_),
    .B(_12097_),
    .Y(_12633_));
 sky130_fd_sc_hd__nand3b_2 _34276_ (.A_N(_12633_),
    .B(_05773_),
    .C(_10913_),
    .Y(_12634_));
 sky130_fd_sc_hd__o2bb2ai_2 _34277_ (.A1_N(_12632_),
    .A2_N(_12634_),
    .B1(_11487_),
    .B2(_06248_),
    .Y(_12635_));
 sky130_fd_sc_hd__and2_2 _34278_ (.A(\pcpi_mul.rs1[32] ),
    .B(\pcpi_mul.rs2[6] ),
    .X(_12636_));
 sky130_fd_sc_hd__buf_1 _34279_ (.A(_12636_),
    .X(_12637_));
 sky130_fd_sc_hd__nand3_2 _34280_ (.A(_12634_),
    .B(_12632_),
    .C(_12637_),
    .Y(_12638_));
 sky130_fd_sc_hd__nand2_2 _34281_ (.A(_12318_),
    .B(_12319_),
    .Y(_12639_));
 sky130_fd_sc_hd__nor2_2 _34282_ (.A(_12318_),
    .B(_12319_),
    .Y(_12640_));
 sky130_fd_sc_hd__a21oi_2 _34283_ (.A1(_12639_),
    .A2(_12317_),
    .B1(_12640_),
    .Y(_12641_));
 sky130_vsdinv _34284_ (.A(_12641_),
    .Y(_12642_));
 sky130_fd_sc_hd__a21o_2 _34285_ (.A1(_12635_),
    .A2(_12638_),
    .B1(_12642_),
    .X(_12643_));
 sky130_fd_sc_hd__nand3_2 _34286_ (.A(_12635_),
    .B(_12642_),
    .C(_12638_),
    .Y(_12644_));
 sky130_fd_sc_hd__nand2_2 _34287_ (.A(_12643_),
    .B(_12644_),
    .Y(_12645_));
 sky130_fd_sc_hd__a21boi_2 _34288_ (.A1(_12386_),
    .A2(_12391_),
    .B1_N(_12388_),
    .Y(_12646_));
 sky130_fd_sc_hd__nand2_2 _34289_ (.A(_12645_),
    .B(_12646_),
    .Y(_12647_));
 sky130_fd_sc_hd__nand3b_2 _34290_ (.A_N(_12646_),
    .B(_12643_),
    .C(_12644_),
    .Y(_12648_));
 sky130_fd_sc_hd__a21oi_2 _34291_ (.A1(_12328_),
    .A2(_12332_),
    .B1(_12333_),
    .Y(_12649_));
 sky130_fd_sc_hd__o21ai_2 _34292_ (.A1(_12649_),
    .A2(_12321_),
    .B1(_12335_),
    .Y(_12650_));
 sky130_fd_sc_hd__a21oi_2 _34293_ (.A1(_12647_),
    .A2(_12648_),
    .B1(_12650_),
    .Y(_12651_));
 sky130_fd_sc_hd__nand3_2 _34294_ (.A(_12647_),
    .B(_12650_),
    .C(_12648_),
    .Y(_12652_));
 sky130_vsdinv _34295_ (.A(_12652_),
    .Y(_12653_));
 sky130_vsdinv _34296_ (.A(_12398_),
    .Y(_12654_));
 sky130_fd_sc_hd__a21oi_2 _34297_ (.A1(_12397_),
    .A2(_12400_),
    .B1(_12654_),
    .Y(_12655_));
 sky130_vsdinv _34298_ (.A(_12655_),
    .Y(_12656_));
 sky130_fd_sc_hd__o21bai_2 _34299_ (.A1(_12651_),
    .A2(_12653_),
    .B1_N(_12656_),
    .Y(_12657_));
 sky130_fd_sc_hd__nand3b_2 _34300_ (.A_N(_12651_),
    .B(_12656_),
    .C(_12652_),
    .Y(_12658_));
 sky130_fd_sc_hd__nand2_2 _34301_ (.A(_12657_),
    .B(_12658_),
    .Y(_12659_));
 sky130_fd_sc_hd__a21boi_2 _34302_ (.A1(_12405_),
    .A2(_12409_),
    .B1_N(_12407_),
    .Y(_12660_));
 sky130_fd_sc_hd__nand2_2 _34303_ (.A(_12659_),
    .B(_12660_),
    .Y(_12661_));
 sky130_fd_sc_hd__nand3b_2 _34304_ (.A_N(_12660_),
    .B(_12658_),
    .C(_12657_),
    .Y(_12662_));
 sky130_vsdinv _34305_ (.A(_12369_),
    .Y(_12663_));
 sky130_fd_sc_hd__nand2_2 _34306_ (.A(_12663_),
    .B(_10883_),
    .Y(_12664_));
 sky130_fd_sc_hd__o21a_2 _34307_ (.A1(_10884_),
    .A2(_12367_),
    .B1(_12664_),
    .X(_12665_));
 sky130_fd_sc_hd__xor2_2 _34308_ (.A(_12665_),
    .B(_11835_),
    .X(_12666_));
 sky130_fd_sc_hd__nand3b_2 _34309_ (.A_N(_12666_),
    .B(_12381_),
    .C(_12664_),
    .Y(_12667_));
 sky130_vsdinv _34310_ (.A(_12664_),
    .Y(_12668_));
 sky130_fd_sc_hd__o21ai_2 _34311_ (.A1(_12668_),
    .A2(_12380_),
    .B1(_12666_),
    .Y(_12669_));
 sky130_fd_sc_hd__a21o_2 _34312_ (.A1(_12667_),
    .A2(_12669_),
    .B1(_12118_),
    .X(_12670_));
 sky130_fd_sc_hd__nand3_2 _34313_ (.A(_12667_),
    .B(_12442_),
    .C(_12669_),
    .Y(_12671_));
 sky130_fd_sc_hd__nand2_2 _34314_ (.A(_12670_),
    .B(_12671_),
    .Y(_12672_));
 sky130_fd_sc_hd__a21boi_2 _34315_ (.A1(_12661_),
    .A2(_12662_),
    .B1_N(_12672_),
    .Y(_12673_));
 sky130_fd_sc_hd__nand2_2 _34316_ (.A(_12661_),
    .B(_12662_),
    .Y(_12674_));
 sky130_fd_sc_hd__nor2_2 _34317_ (.A(_12672_),
    .B(_12674_),
    .Y(_12675_));
 sky130_fd_sc_hd__a21oi_2 _34318_ (.A1(_12345_),
    .A2(_12346_),
    .B1(_12343_),
    .Y(_12676_));
 sky130_fd_sc_hd__o21ai_2 _34319_ (.A1(_12349_),
    .A2(_12676_),
    .B1(_12347_),
    .Y(_12677_));
 sky130_fd_sc_hd__o21bai_2 _34320_ (.A1(_12673_),
    .A2(_12675_),
    .B1_N(_12677_),
    .Y(_12678_));
 sky130_fd_sc_hd__nand3b_2 _34321_ (.A_N(_12672_),
    .B(_12662_),
    .C(_12661_),
    .Y(_12679_));
 sky130_fd_sc_hd__nand3b_2 _34322_ (.A_N(_12673_),
    .B(_12677_),
    .C(_12679_),
    .Y(_12680_));
 sky130_fd_sc_hd__buf_1 _34323_ (.A(_12680_),
    .X(_12681_));
 sky130_vsdinv _34324_ (.A(_12416_),
    .Y(_12682_));
 sky130_fd_sc_hd__a31oi_2 _34325_ (.A1(_12414_),
    .A2(_12384_),
    .A3(_12385_),
    .B1(_12682_),
    .Y(_12683_));
 sky130_fd_sc_hd__a21boi_2 _34326_ (.A1(_12678_),
    .A2(_12681_),
    .B1_N(_12683_),
    .Y(_12684_));
 sky130_fd_sc_hd__o211a_2 _34327_ (.A1(_12682_),
    .A2(_12420_),
    .B1(_12681_),
    .C1(_12678_),
    .X(_12685_));
 sky130_fd_sc_hd__nor2_2 _34328_ (.A(_12684_),
    .B(_12685_),
    .Y(_12686_));
 sky130_fd_sc_hd__a21oi_2 _34329_ (.A1(_12628_),
    .A2(_12631_),
    .B1(_12686_),
    .Y(_12687_));
 sky130_fd_sc_hd__nand2_2 _34330_ (.A(_12678_),
    .B(_12680_),
    .Y(_12688_));
 sky130_fd_sc_hd__nand2_2 _34331_ (.A(_12688_),
    .B(_12683_),
    .Y(_12689_));
 sky130_fd_sc_hd__nand3b_2 _34332_ (.A_N(_12683_),
    .B(_12678_),
    .C(_12680_),
    .Y(_12690_));
 sky130_fd_sc_hd__nand2_2 _34333_ (.A(_12689_),
    .B(_12690_),
    .Y(_12691_));
 sky130_fd_sc_hd__a21oi_2 _34334_ (.A1(_12621_),
    .A2(_12625_),
    .B1(_12629_),
    .Y(_12692_));
 sky130_vsdinv _34335_ (.A(_12631_),
    .Y(_12693_));
 sky130_fd_sc_hd__nor3_2 _34336_ (.A(_12691_),
    .B(_12692_),
    .C(_12693_),
    .Y(_12694_));
 sky130_fd_sc_hd__o21ai_2 _34337_ (.A1(_12431_),
    .A2(_12433_),
    .B1(_12365_),
    .Y(_12695_));
 sky130_fd_sc_hd__o21bai_2 _34338_ (.A1(_12687_),
    .A2(_12694_),
    .B1_N(_12695_),
    .Y(_12696_));
 sky130_fd_sc_hd__nand2_2 _34339_ (.A(_12628_),
    .B(_12630_),
    .Y(_12697_));
 sky130_fd_sc_hd__nand2_2 _34340_ (.A(_12697_),
    .B(_12691_),
    .Y(_12698_));
 sky130_fd_sc_hd__nand3_2 _34341_ (.A(_12686_),
    .B(_12628_),
    .C(_12631_),
    .Y(_12699_));
 sky130_fd_sc_hd__nand3_2 _34342_ (.A(_12698_),
    .B(_12695_),
    .C(_12699_),
    .Y(_12700_));
 sky130_fd_sc_hd__buf_1 _34343_ (.A(_12700_),
    .X(_12701_));
 sky130_fd_sc_hd__a21boi_2 _34344_ (.A1(_12442_),
    .A2(_12383_),
    .B1_N(_12382_),
    .Y(_12702_));
 sky130_fd_sc_hd__nand2_2 _34345_ (.A(_12429_),
    .B(_12425_),
    .Y(_12703_));
 sky130_fd_sc_hd__xnor2_2 _34346_ (.A(_12702_),
    .B(_12703_),
    .Y(_12704_));
 sky130_fd_sc_hd__a21oi_2 _34347_ (.A1(_12696_),
    .A2(_12701_),
    .B1(_12704_),
    .Y(_12705_));
 sky130_vsdinv _34348_ (.A(_12704_),
    .Y(_12706_));
 sky130_fd_sc_hd__a21oi_2 _34349_ (.A1(_12698_),
    .A2(_12699_),
    .B1(_12695_),
    .Y(_12707_));
 sky130_vsdinv _34350_ (.A(_12701_),
    .Y(_12708_));
 sky130_fd_sc_hd__nor3_2 _34351_ (.A(_12706_),
    .B(_12707_),
    .C(_12708_),
    .Y(_12709_));
 sky130_fd_sc_hd__a21oi_2 _34352_ (.A1(_12438_),
    .A2(_12439_),
    .B1(_12436_),
    .Y(_12710_));
 sky130_fd_sc_hd__o21ai_2 _34353_ (.A1(_12452_),
    .A2(_12710_),
    .B1(_12441_),
    .Y(_12711_));
 sky130_fd_sc_hd__o21bai_2 _34354_ (.A1(_12705_),
    .A2(_12709_),
    .B1_N(_12711_),
    .Y(_12712_));
 sky130_fd_sc_hd__nand2_2 _34355_ (.A(_12696_),
    .B(_12700_),
    .Y(_12713_));
 sky130_fd_sc_hd__nand2_2 _34356_ (.A(_12713_),
    .B(_12706_),
    .Y(_12714_));
 sky130_fd_sc_hd__nand3_2 _34357_ (.A(_12696_),
    .B(_12704_),
    .C(_12701_),
    .Y(_12715_));
 sky130_fd_sc_hd__nand3_2 _34358_ (.A(_12714_),
    .B(_12711_),
    .C(_12715_),
    .Y(_12716_));
 sky130_fd_sc_hd__a21oi_2 _34359_ (.A1(_12139_),
    .A2(_12131_),
    .B1(_12443_),
    .Y(_12717_));
 sky130_fd_sc_hd__a21oi_2 _34360_ (.A1(_12712_),
    .A2(_12716_),
    .B1(_12717_),
    .Y(_12718_));
 sky130_vsdinv _34361_ (.A(_12717_),
    .Y(_12719_));
 sky130_fd_sc_hd__a21oi_2 _34362_ (.A1(_12714_),
    .A2(_12715_),
    .B1(_12711_),
    .Y(_12720_));
 sky130_fd_sc_hd__a21boi_2 _34363_ (.A1(_12437_),
    .A2(_12445_),
    .B1_N(_12441_),
    .Y(_12721_));
 sky130_fd_sc_hd__nor3_2 _34364_ (.A(_12705_),
    .B(_12721_),
    .C(_12709_),
    .Y(_12722_));
 sky130_fd_sc_hd__nor3_2 _34365_ (.A(_12719_),
    .B(_12720_),
    .C(_12722_),
    .Y(_12723_));
 sky130_vsdinv _34366_ (.A(_12455_),
    .Y(_12724_));
 sky130_fd_sc_hd__a21oi_2 _34367_ (.A1(_12453_),
    .A2(_12447_),
    .B1(_12449_),
    .Y(_12725_));
 sky130_fd_sc_hd__o21ai_2 _34368_ (.A1(_12724_),
    .A2(_12725_),
    .B1(_12454_),
    .Y(_12726_));
 sky130_fd_sc_hd__o21bai_2 _34369_ (.A1(_12718_),
    .A2(_12723_),
    .B1_N(_12726_),
    .Y(_12727_));
 sky130_fd_sc_hd__o21bai_2 _34370_ (.A1(_12720_),
    .A2(_12722_),
    .B1_N(_12717_),
    .Y(_12728_));
 sky130_fd_sc_hd__nand3_2 _34371_ (.A(_12712_),
    .B(_12717_),
    .C(_12716_),
    .Y(_12729_));
 sky130_fd_sc_hd__nand3_2 _34372_ (.A(_12728_),
    .B(_12726_),
    .C(_12729_),
    .Y(_12730_));
 sky130_fd_sc_hd__and2_2 _34373_ (.A(_12727_),
    .B(_12730_),
    .X(_12731_));
 sky130_fd_sc_hd__nand2_2 _34374_ (.A(_12462_),
    .B(_12175_),
    .Y(_12732_));
 sky130_fd_sc_hd__nand2_2 _34375_ (.A(_12732_),
    .B(_12460_),
    .Y(_12733_));
 sky130_fd_sc_hd__o31ai_2 _34376_ (.A1(_12176_),
    .A2(_12463_),
    .A3(_12182_),
    .B1(_12733_),
    .Y(_12734_));
 sky130_fd_sc_hd__xor2_2 _34377_ (.A(_12731_),
    .B(_12734_),
    .X(_02657_));
 sky130_fd_sc_hd__nand2_2 _34378_ (.A(_10480_),
    .B(_05840_),
    .Y(_12735_));
 sky130_fd_sc_hd__nand3b_2 _34379_ (.A_N(_12735_),
    .B(_10996_),
    .C(_19268_),
    .Y(_12736_));
 sky130_fd_sc_hd__o21ai_2 _34380_ (.A1(_08007_),
    .A2(_11004_),
    .B1(_12735_),
    .Y(_12737_));
 sky130_fd_sc_hd__and2_2 _34381_ (.A(_10483_),
    .B(_06342_),
    .X(_12738_));
 sky130_fd_sc_hd__a21oi_2 _34382_ (.A1(_12736_),
    .A2(_12737_),
    .B1(_12738_),
    .Y(_12739_));
 sky130_fd_sc_hd__nand3_2 _34383_ (.A(_12736_),
    .B(_12738_),
    .C(_12737_),
    .Y(_12740_));
 sky130_vsdinv _34384_ (.A(_12740_),
    .Y(_12741_));
 sky130_fd_sc_hd__a21oi_2 _34385_ (.A1(_12469_),
    .A2(_12470_),
    .B1(_12479_),
    .Y(_12742_));
 sky130_fd_sc_hd__o21ai_2 _34386_ (.A1(_12739_),
    .A2(_12741_),
    .B1(_12742_),
    .Y(_12743_));
 sky130_fd_sc_hd__a21o_2 _34387_ (.A1(_12736_),
    .A2(_12737_),
    .B1(_12738_),
    .X(_12744_));
 sky130_fd_sc_hd__nand3b_2 _34388_ (.A_N(_12742_),
    .B(_12744_),
    .C(_12740_),
    .Y(_12745_));
 sky130_fd_sc_hd__nand2_2 _34389_ (.A(_09957_),
    .B(_19252_),
    .Y(_12746_));
 sky130_fd_sc_hd__nand2_2 _34390_ (.A(_18716_),
    .B(_08905_),
    .Y(_12747_));
 sky130_fd_sc_hd__nor2_2 _34391_ (.A(_12746_),
    .B(_12747_),
    .Y(_12748_));
 sky130_fd_sc_hd__and2_2 _34392_ (.A(_09605_),
    .B(_19242_),
    .X(_12749_));
 sky130_fd_sc_hd__nand2_2 _34393_ (.A(_12746_),
    .B(_12747_),
    .Y(_12750_));
 sky130_fd_sc_hd__nand3b_2 _34394_ (.A_N(_12748_),
    .B(_12749_),
    .C(_12750_),
    .Y(_12751_));
 sky130_fd_sc_hd__a22oi_2 _34395_ (.A1(_11618_),
    .A2(_09340_),
    .B1(_11340_),
    .B2(_06047_),
    .Y(_12752_));
 sky130_fd_sc_hd__o21bai_2 _34396_ (.A1(_12752_),
    .A2(_12748_),
    .B1_N(_12749_),
    .Y(_12753_));
 sky130_fd_sc_hd__nand2_2 _34397_ (.A(_12751_),
    .B(_12753_),
    .Y(_12754_));
 sky130_vsdinv _34398_ (.A(_12754_),
    .Y(_12755_));
 sky130_fd_sc_hd__a21oi_2 _34399_ (.A1(_12743_),
    .A2(_12745_),
    .B1(_12755_),
    .Y(_12756_));
 sky130_fd_sc_hd__nand3_2 _34400_ (.A(_12743_),
    .B(_12755_),
    .C(_12745_),
    .Y(_12757_));
 sky130_vsdinv _34401_ (.A(_12757_),
    .Y(_12758_));
 sky130_fd_sc_hd__o21ai_2 _34402_ (.A1(_12489_),
    .A2(_12492_),
    .B1(_12481_),
    .Y(_12759_));
 sky130_fd_sc_hd__o21bai_2 _34403_ (.A1(_12756_),
    .A2(_12758_),
    .B1_N(_12759_),
    .Y(_12760_));
 sky130_fd_sc_hd__nand2_2 _34404_ (.A(_12743_),
    .B(_12745_),
    .Y(_12761_));
 sky130_fd_sc_hd__nand2_2 _34405_ (.A(_12761_),
    .B(_12754_),
    .Y(_12762_));
 sky130_fd_sc_hd__nand3_2 _34406_ (.A(_12762_),
    .B(_12757_),
    .C(_12759_),
    .Y(_12763_));
 sky130_fd_sc_hd__a22o_2 _34407_ (.A1(_09312_),
    .A2(_08054_),
    .B1(_10456_),
    .B2(_07314_),
    .X(_12764_));
 sky130_fd_sc_hd__nand2_2 _34408_ (.A(_10452_),
    .B(_07100_),
    .Y(_12765_));
 sky130_fd_sc_hd__nand3b_2 _34409_ (.A_N(_12765_),
    .B(_12217_),
    .C(_10743_),
    .Y(_12766_));
 sky130_fd_sc_hd__o2bb2ai_2 _34410_ (.A1_N(_12764_),
    .A2_N(_12766_),
    .B1(_12219_),
    .B2(_19227_),
    .Y(_12767_));
 sky130_fd_sc_hd__and2_2 _34411_ (.A(_10703_),
    .B(_07906_),
    .X(_12768_));
 sky130_fd_sc_hd__nand3_2 _34412_ (.A(_12766_),
    .B(_12764_),
    .C(_12768_),
    .Y(_12769_));
 sky130_fd_sc_hd__o31ai_2 _34413_ (.A1(_18725_),
    .A2(_19250_),
    .A3(_12482_),
    .B1(_12487_),
    .Y(_12770_));
 sky130_fd_sc_hd__a21o_2 _34414_ (.A1(_12767_),
    .A2(_12769_),
    .B1(_12770_),
    .X(_12771_));
 sky130_fd_sc_hd__nand3_2 _34415_ (.A(_12770_),
    .B(_12767_),
    .C(_12769_),
    .Y(_12772_));
 sky130_fd_sc_hd__nand2_2 _34416_ (.A(_12771_),
    .B(_12772_),
    .Y(_12773_));
 sky130_fd_sc_hd__a21boi_2 _34417_ (.A1(_12505_),
    .A2(_12501_),
    .B1_N(_12503_),
    .Y(_12774_));
 sky130_fd_sc_hd__nand2_2 _34418_ (.A(_12773_),
    .B(_12774_),
    .Y(_12775_));
 sky130_fd_sc_hd__nand3b_2 _34419_ (.A_N(_12774_),
    .B(_12771_),
    .C(_12772_),
    .Y(_12776_));
 sky130_fd_sc_hd__nand2_2 _34420_ (.A(_12775_),
    .B(_12776_),
    .Y(_12777_));
 sky130_fd_sc_hd__buf_1 _34421_ (.A(_12777_),
    .X(_12778_));
 sky130_fd_sc_hd__a21boi_2 _34422_ (.A1(_12760_),
    .A2(_12763_),
    .B1_N(_12778_),
    .Y(_12779_));
 sky130_fd_sc_hd__a21oi_2 _34423_ (.A1(_12762_),
    .A2(_12757_),
    .B1(_12759_),
    .Y(_12780_));
 sky130_vsdinv _34424_ (.A(_12763_),
    .Y(_12781_));
 sky130_fd_sc_hd__nor3_2 _34425_ (.A(_12778_),
    .B(_12780_),
    .C(_12781_),
    .Y(_12782_));
 sky130_fd_sc_hd__o21ai_2 _34426_ (.A1(_12515_),
    .A2(_12517_),
    .B1(_12499_),
    .Y(_12783_));
 sky130_fd_sc_hd__o21bai_2 _34427_ (.A1(_12779_),
    .A2(_12782_),
    .B1_N(_12783_),
    .Y(_12784_));
 sky130_fd_sc_hd__o21ai_2 _34428_ (.A1(_12780_),
    .A2(_12781_),
    .B1(_12778_),
    .Y(_12785_));
 sky130_fd_sc_hd__nand3b_2 _34429_ (.A_N(_12778_),
    .B(_12760_),
    .C(_12763_),
    .Y(_12786_));
 sky130_fd_sc_hd__nand3_2 _34430_ (.A(_12785_),
    .B(_12786_),
    .C(_12783_),
    .Y(_12787_));
 sky130_fd_sc_hd__buf_1 _34431_ (.A(_12787_),
    .X(_12788_));
 sky130_fd_sc_hd__a21boi_2 _34432_ (.A1(_12532_),
    .A2(_12526_),
    .B1_N(_12529_),
    .Y(_12789_));
 sky130_fd_sc_hd__nand2_2 _34433_ (.A(_10417_),
    .B(_10150_),
    .Y(_12790_));
 sky130_fd_sc_hd__buf_1 _34434_ (.A(_11968_),
    .X(_12791_));
 sky130_fd_sc_hd__nand3b_2 _34435_ (.A_N(_12790_),
    .B(_12791_),
    .C(_11110_),
    .Y(_12792_));
 sky130_fd_sc_hd__and2_2 _34436_ (.A(_07845_),
    .B(_07942_),
    .X(_12793_));
 sky130_fd_sc_hd__buf_1 _34437_ (.A(_09263_),
    .X(_12794_));
 sky130_fd_sc_hd__nand2_2 _34438_ (.A(_12794_),
    .B(_06937_),
    .Y(_12795_));
 sky130_fd_sc_hd__nand2_2 _34439_ (.A(_12790_),
    .B(_12795_),
    .Y(_12796_));
 sky130_fd_sc_hd__nand3_2 _34440_ (.A(_12792_),
    .B(_12793_),
    .C(_12796_),
    .Y(_12797_));
 sky130_fd_sc_hd__o2bb2ai_2 _34441_ (.A1_N(_12796_),
    .A2_N(_12792_),
    .B1(_08232_),
    .B2(_19209_),
    .Y(_12798_));
 sky130_fd_sc_hd__nand3b_2 _34442_ (.A_N(_12789_),
    .B(_12797_),
    .C(_12798_),
    .Y(_12799_));
 sky130_fd_sc_hd__nand2_2 _34443_ (.A(_12798_),
    .B(_12797_),
    .Y(_12800_));
 sky130_fd_sc_hd__nand2_2 _34444_ (.A(_12800_),
    .B(_12789_),
    .Y(_12801_));
 sky130_fd_sc_hd__and2_2 _34445_ (.A(_07161_),
    .B(_08571_),
    .X(_12802_));
 sky130_fd_sc_hd__nand2_2 _34446_ (.A(_11067_),
    .B(_08549_),
    .Y(_12803_));
 sky130_fd_sc_hd__nand3b_2 _34447_ (.A_N(_12803_),
    .B(_10429_),
    .C(_11714_),
    .Y(_12804_));
 sky130_fd_sc_hd__buf_1 _34448_ (.A(_08074_),
    .X(_12805_));
 sky130_fd_sc_hd__buf_1 _34449_ (.A(_07853_),
    .X(_12806_));
 sky130_fd_sc_hd__a22o_2 _34450_ (.A1(_12805_),
    .A2(_11714_),
    .B1(_12806_),
    .B2(_12288_),
    .X(_12807_));
 sky130_fd_sc_hd__nand2_2 _34451_ (.A(_12804_),
    .B(_12807_),
    .Y(_12808_));
 sky130_fd_sc_hd__xnor2_2 _34452_ (.A(_12802_),
    .B(_12808_),
    .Y(_12809_));
 sky130_fd_sc_hd__a21o_2 _34453_ (.A1(_12799_),
    .A2(_12801_),
    .B1(_12809_),
    .X(_12810_));
 sky130_fd_sc_hd__nand3_2 _34454_ (.A(_12799_),
    .B(_12801_),
    .C(_12809_),
    .Y(_12811_));
 sky130_fd_sc_hd__nand2_2 _34455_ (.A(_12513_),
    .B(_12509_),
    .Y(_12812_));
 sky130_fd_sc_hd__a21o_2 _34456_ (.A1(_12810_),
    .A2(_12811_),
    .B1(_12812_),
    .X(_12813_));
 sky130_fd_sc_hd__nand3_2 _34457_ (.A(_12812_),
    .B(_12810_),
    .C(_12811_),
    .Y(_12814_));
 sky130_vsdinv _34458_ (.A(_12537_),
    .Y(_12815_));
 sky130_fd_sc_hd__a21oi_2 _34459_ (.A1(_12544_),
    .A2(_12536_),
    .B1(_12815_),
    .Y(_12816_));
 sky130_vsdinv _34460_ (.A(_12816_),
    .Y(_12817_));
 sky130_fd_sc_hd__a21oi_2 _34461_ (.A1(_12813_),
    .A2(_12814_),
    .B1(_12817_),
    .Y(_12818_));
 sky130_fd_sc_hd__nand3_2 _34462_ (.A(_12813_),
    .B(_12817_),
    .C(_12814_),
    .Y(_12819_));
 sky130_vsdinv _34463_ (.A(_12819_),
    .Y(_12820_));
 sky130_fd_sc_hd__nor2_2 _34464_ (.A(_12818_),
    .B(_12820_),
    .Y(_12821_));
 sky130_fd_sc_hd__a21oi_2 _34465_ (.A1(_12784_),
    .A2(_12788_),
    .B1(_12821_),
    .Y(_12822_));
 sky130_fd_sc_hd__a21oi_2 _34466_ (.A1(_12810_),
    .A2(_12811_),
    .B1(_12812_),
    .Y(_12823_));
 sky130_vsdinv _34467_ (.A(_12814_),
    .Y(_12824_));
 sky130_fd_sc_hd__o21bai_2 _34468_ (.A1(_12823_),
    .A2(_12824_),
    .B1_N(_12817_),
    .Y(_12825_));
 sky130_fd_sc_hd__nand2_2 _34469_ (.A(_12825_),
    .B(_12819_),
    .Y(_12826_));
 sky130_fd_sc_hd__a21oi_2 _34470_ (.A1(_12785_),
    .A2(_12786_),
    .B1(_12783_),
    .Y(_12827_));
 sky130_vsdinv _34471_ (.A(_12788_),
    .Y(_12828_));
 sky130_fd_sc_hd__nor3_2 _34472_ (.A(_12826_),
    .B(_12827_),
    .C(_12828_),
    .Y(_12829_));
 sky130_fd_sc_hd__o21ai_2 _34473_ (.A1(_12561_),
    .A2(_12562_),
    .B1(_12524_),
    .Y(_12830_));
 sky130_fd_sc_hd__o21bai_2 _34474_ (.A1(_12822_),
    .A2(_12829_),
    .B1_N(_12830_),
    .Y(_12831_));
 sky130_fd_sc_hd__o2bb2ai_2 _34475_ (.A1_N(_12788_),
    .A2_N(_12784_),
    .B1(_12820_),
    .B2(_12818_),
    .Y(_12832_));
 sky130_fd_sc_hd__nand3_2 _34476_ (.A(_12821_),
    .B(_12784_),
    .C(_12788_),
    .Y(_12833_));
 sky130_fd_sc_hd__nand3_2 _34477_ (.A(_12832_),
    .B(_12833_),
    .C(_12830_),
    .Y(_12834_));
 sky130_fd_sc_hd__nand2_2 _34478_ (.A(_12831_),
    .B(_12834_),
    .Y(_12835_));
 sky130_fd_sc_hd__buf_1 _34479_ (.A(_09495_),
    .X(_12836_));
 sky130_fd_sc_hd__a22o_2 _34480_ (.A1(_11108_),
    .A2(_07952_),
    .B1(_08142_),
    .B2(_12836_),
    .X(_12837_));
 sky130_fd_sc_hd__nand2_2 _34481_ (.A(_07392_),
    .B(_09755_),
    .Y(_12838_));
 sky130_fd_sc_hd__buf_1 _34482_ (.A(_08295_),
    .X(_12839_));
 sky130_fd_sc_hd__nand3b_2 _34483_ (.A_N(_12838_),
    .B(_12289_),
    .C(_12839_),
    .Y(_12840_));
 sky130_fd_sc_hd__o2bb2ai_2 _34484_ (.A1_N(_12837_),
    .A2_N(_12840_),
    .B1(_08918_),
    .B2(_19174_),
    .Y(_12841_));
 sky130_fd_sc_hd__buf_1 _34485_ (.A(_08556_),
    .X(_12842_));
 sky130_fd_sc_hd__and2_2 _34486_ (.A(_07402_),
    .B(_12842_),
    .X(_12843_));
 sky130_fd_sc_hd__nand3_2 _34487_ (.A(_12840_),
    .B(_12837_),
    .C(_12843_),
    .Y(_12844_));
 sky130_fd_sc_hd__buf_1 _34488_ (.A(_19197_),
    .X(_12845_));
 sky130_fd_sc_hd__a22oi_2 _34489_ (.A1(_10429_),
    .A2(_10379_),
    .B1(_08220_),
    .B2(_07967_),
    .Y(_12846_));
 sky130_fd_sc_hd__buf_1 _34490_ (.A(_18765_),
    .X(_12847_));
 sky130_fd_sc_hd__nand3b_2 _34491_ (.A_N(_12542_),
    .B(_12847_),
    .C(_10379_),
    .Y(_12848_));
 sky130_fd_sc_hd__o31ai_2 _34492_ (.A1(_18777_),
    .A2(_12845_),
    .A3(_12846_),
    .B1(_12848_),
    .Y(_12849_));
 sky130_fd_sc_hd__a21o_2 _34493_ (.A1(_12841_),
    .A2(_12844_),
    .B1(_12849_),
    .X(_12850_));
 sky130_fd_sc_hd__nand3_2 _34494_ (.A(_12849_),
    .B(_12841_),
    .C(_12844_),
    .Y(_12851_));
 sky130_fd_sc_hd__a21boi_2 _34495_ (.A1(_12571_),
    .A2(_12575_),
    .B1_N(_12573_),
    .Y(_12852_));
 sky130_vsdinv _34496_ (.A(_12852_),
    .Y(_12853_));
 sky130_fd_sc_hd__a21o_2 _34497_ (.A1(_12850_),
    .A2(_12851_),
    .B1(_12853_),
    .X(_12854_));
 sky130_fd_sc_hd__nand3_2 _34498_ (.A(_12850_),
    .B(_12853_),
    .C(_12851_),
    .Y(_12855_));
 sky130_fd_sc_hd__nand2_2 _34499_ (.A(_12583_),
    .B(_12579_),
    .Y(_12856_));
 sky130_fd_sc_hd__a21o_2 _34500_ (.A1(_12854_),
    .A2(_12855_),
    .B1(_12856_),
    .X(_12857_));
 sky130_fd_sc_hd__nand3_2 _34501_ (.A(_12856_),
    .B(_12854_),
    .C(_12855_),
    .Y(_12858_));
 sky130_fd_sc_hd__buf_1 _34502_ (.A(_09787_),
    .X(_12859_));
 sky130_fd_sc_hd__nand3b_2 _34503_ (.A_N(_12593_),
    .B(_18804_),
    .C(_12859_),
    .Y(_12860_));
 sky130_fd_sc_hd__nand2_2 _34504_ (.A(_06534_),
    .B(_08818_),
    .Y(_12861_));
 sky130_fd_sc_hd__nand2_2 _34505_ (.A(_08688_),
    .B(_10531_),
    .Y(_12862_));
 sky130_fd_sc_hd__nand2_2 _34506_ (.A(_12861_),
    .B(_12862_),
    .Y(_12863_));
 sky130_fd_sc_hd__nand3b_2 _34507_ (.A_N(_12861_),
    .B(_18803_),
    .C(_10538_),
    .Y(_12864_));
 sky130_fd_sc_hd__o2bb2ai_2 _34508_ (.A1_N(_12863_),
    .A2_N(_12864_),
    .B1(_11745_),
    .B2(_19158_),
    .Y(_12865_));
 sky130_fd_sc_hd__and2_2 _34509_ (.A(_10382_),
    .B(_10533_),
    .X(_12866_));
 sky130_fd_sc_hd__nand3_2 _34510_ (.A(_12864_),
    .B(_12866_),
    .C(_12863_),
    .Y(_12867_));
 sky130_fd_sc_hd__nand2_2 _34511_ (.A(_12865_),
    .B(_12867_),
    .Y(_12868_));
 sky130_fd_sc_hd__a21o_2 _34512_ (.A1(_12597_),
    .A2(_12860_),
    .B1(_12868_),
    .X(_12869_));
 sky130_fd_sc_hd__nand3_2 _34513_ (.A(_12868_),
    .B(_12860_),
    .C(_12598_),
    .Y(_12870_));
 sky130_fd_sc_hd__buf_1 _34514_ (.A(_19138_),
    .X(_12871_));
 sky130_fd_sc_hd__and2_2 _34515_ (.A(_06680_),
    .B(_12871_),
    .X(_12872_));
 sky130_fd_sc_hd__nand2_2 _34516_ (.A(_06671_),
    .B(_10877_),
    .Y(_12873_));
 sky130_fd_sc_hd__nand2_2 _34517_ (.A(_06674_),
    .B(_11791_),
    .Y(_12874_));
 sky130_fd_sc_hd__xnor2_2 _34518_ (.A(_12873_),
    .B(_12874_),
    .Y(_12875_));
 sky130_fd_sc_hd__xnor2_2 _34519_ (.A(_12872_),
    .B(_12875_),
    .Y(_12876_));
 sky130_fd_sc_hd__a21o_2 _34520_ (.A1(_12869_),
    .A2(_12870_),
    .B1(_12876_),
    .X(_12877_));
 sky130_fd_sc_hd__nand3_2 _34521_ (.A(_12869_),
    .B(_12870_),
    .C(_12876_),
    .Y(_12878_));
 sky130_fd_sc_hd__nand2_2 _34522_ (.A(_12877_),
    .B(_12878_),
    .Y(_12879_));
 sky130_fd_sc_hd__a21boi_2 _34523_ (.A1(_12857_),
    .A2(_12858_),
    .B1_N(_12879_),
    .Y(_12880_));
 sky130_fd_sc_hd__nand2_2 _34524_ (.A(_12857_),
    .B(_12858_),
    .Y(_12881_));
 sky130_fd_sc_hd__nor2_2 _34525_ (.A(_12879_),
    .B(_12881_),
    .Y(_12882_));
 sky130_fd_sc_hd__nand2_2 _34526_ (.A(_12555_),
    .B(_12551_),
    .Y(_12883_));
 sky130_fd_sc_hd__o21bai_2 _34527_ (.A1(_12880_),
    .A2(_12882_),
    .B1_N(_12883_),
    .Y(_12884_));
 sky130_fd_sc_hd__nand3b_2 _34528_ (.A_N(_12879_),
    .B(_12857_),
    .C(_12858_),
    .Y(_12885_));
 sky130_fd_sc_hd__nand3b_2 _34529_ (.A_N(_12880_),
    .B(_12883_),
    .C(_12885_),
    .Y(_12886_));
 sky130_fd_sc_hd__buf_1 _34530_ (.A(_12886_),
    .X(_12887_));
 sky130_fd_sc_hd__a21boi_2 _34531_ (.A1(_12587_),
    .A2(_12609_),
    .B1_N(_12585_),
    .Y(_12888_));
 sky130_vsdinv _34532_ (.A(_12888_),
    .Y(_12889_));
 sky130_fd_sc_hd__a21o_2 _34533_ (.A1(_12884_),
    .A2(_12887_),
    .B1(_12889_),
    .X(_12890_));
 sky130_fd_sc_hd__nand3_2 _34534_ (.A(_12884_),
    .B(_12886_),
    .C(_12889_),
    .Y(_12891_));
 sky130_fd_sc_hd__nand2_2 _34535_ (.A(_12890_),
    .B(_12891_),
    .Y(_12892_));
 sky130_fd_sc_hd__nand2_2 _34536_ (.A(_12835_),
    .B(_12892_),
    .Y(_12893_));
 sky130_fd_sc_hd__a21oi_2 _34537_ (.A1(_12884_),
    .A2(_12887_),
    .B1(_12889_),
    .Y(_12894_));
 sky130_vsdinv _34538_ (.A(_12891_),
    .Y(_12895_));
 sky130_fd_sc_hd__nor2_2 _34539_ (.A(_12894_),
    .B(_12895_),
    .Y(_12896_));
 sky130_fd_sc_hd__nand3_2 _34540_ (.A(_12896_),
    .B(_12834_),
    .C(_12831_),
    .Y(_12897_));
 sky130_fd_sc_hd__nand2_2 _34541_ (.A(_12893_),
    .B(_12897_),
    .Y(_12898_));
 sky130_fd_sc_hd__a21oi_2 _34542_ (.A1(_12567_),
    .A2(_12568_),
    .B1(_12565_),
    .Y(_12899_));
 sky130_fd_sc_hd__o21ai_2 _34543_ (.A1(_12620_),
    .A2(_12899_),
    .B1(_12569_),
    .Y(_12900_));
 sky130_vsdinv _34544_ (.A(_12900_),
    .Y(_12901_));
 sky130_fd_sc_hd__nand2_2 _34545_ (.A(_12898_),
    .B(_12901_),
    .Y(_12902_));
 sky130_fd_sc_hd__nand3_2 _34546_ (.A(_12893_),
    .B(_12897_),
    .C(_12900_),
    .Y(_12903_));
 sky130_fd_sc_hd__buf_1 _34547_ (.A(_12903_),
    .X(_12904_));
 sky130_fd_sc_hd__buf_1 _34548_ (.A(_19132_),
    .X(_12905_));
 sky130_fd_sc_hd__a22oi_2 _34549_ (.A1(_12368_),
    .A2(_06097_),
    .B1(_06225_),
    .B2(_12905_),
    .Y(_12906_));
 sky130_fd_sc_hd__nand2_2 _34550_ (.A(_05772_),
    .B(_10899_),
    .Y(_12907_));
 sky130_fd_sc_hd__nand2_2 _34551_ (.A(_10880_),
    .B(\pcpi_mul.rs2[7] ),
    .Y(_12908_));
 sky130_fd_sc_hd__nor2_2 _34552_ (.A(_12907_),
    .B(_12908_),
    .Y(_12909_));
 sky130_vsdinv _34553_ (.A(_12909_),
    .Y(_12910_));
 sky130_fd_sc_hd__nand3b_2 _34554_ (.A_N(_12906_),
    .B(_12910_),
    .C(_12637_),
    .Y(_12911_));
 sky130_fd_sc_hd__o21bai_2 _34555_ (.A1(_12906_),
    .A2(_12909_),
    .B1_N(_12637_),
    .Y(_12912_));
 sky130_fd_sc_hd__nand2_2 _34556_ (.A(_12589_),
    .B(_12590_),
    .Y(_12913_));
 sky130_fd_sc_hd__nor2_2 _34557_ (.A(_12589_),
    .B(_12590_),
    .Y(_12914_));
 sky130_fd_sc_hd__a21oi_2 _34558_ (.A1(_12913_),
    .A2(_12588_),
    .B1(_12914_),
    .Y(_12915_));
 sky130_vsdinv _34559_ (.A(_12915_),
    .Y(_12916_));
 sky130_fd_sc_hd__a21o_2 _34560_ (.A1(_12911_),
    .A2(_12912_),
    .B1(_12916_),
    .X(_12917_));
 sky130_fd_sc_hd__a21boi_2 _34561_ (.A1(_12632_),
    .A2(_12637_),
    .B1_N(_12634_),
    .Y(_12918_));
 sky130_vsdinv _34562_ (.A(_12918_),
    .Y(_12919_));
 sky130_fd_sc_hd__nand3_2 _34563_ (.A(_12916_),
    .B(_12911_),
    .C(_12912_),
    .Y(_12920_));
 sky130_fd_sc_hd__nand3_2 _34564_ (.A(_12917_),
    .B(_12919_),
    .C(_12920_),
    .Y(_12921_));
 sky130_vsdinv _34565_ (.A(_12921_),
    .Y(_12922_));
 sky130_fd_sc_hd__a21oi_2 _34566_ (.A1(_12917_),
    .A2(_12920_),
    .B1(_12919_),
    .Y(_12923_));
 sky130_fd_sc_hd__o21ai_2 _34567_ (.A1(_12592_),
    .A2(_12603_),
    .B1(_12604_),
    .Y(_12924_));
 sky130_fd_sc_hd__o21bai_2 _34568_ (.A1(_12922_),
    .A2(_12923_),
    .B1_N(_12924_),
    .Y(_12925_));
 sky130_fd_sc_hd__nand3b_2 _34569_ (.A_N(_12923_),
    .B(_12924_),
    .C(_12921_),
    .Y(_12926_));
 sky130_fd_sc_hd__buf_1 _34570_ (.A(_12926_),
    .X(_12927_));
 sky130_fd_sc_hd__o21a_2 _34571_ (.A1(_12646_),
    .A2(_12645_),
    .B1(_12644_),
    .X(_12928_));
 sky130_vsdinv _34572_ (.A(_12928_),
    .Y(_12929_));
 sky130_fd_sc_hd__a21oi_2 _34573_ (.A1(_12925_),
    .A2(_12927_),
    .B1(_12929_),
    .Y(_12930_));
 sky130_fd_sc_hd__nand2_2 _34574_ (.A(_12925_),
    .B(_12926_),
    .Y(_12931_));
 sky130_fd_sc_hd__nor2_2 _34575_ (.A(_12928_),
    .B(_12931_),
    .Y(_12932_));
 sky130_fd_sc_hd__o21ai_2 _34576_ (.A1(_12655_),
    .A2(_12651_),
    .B1(_12652_),
    .Y(_12933_));
 sky130_fd_sc_hd__o21bai_2 _34577_ (.A1(_12930_),
    .A2(_12932_),
    .B1_N(_12933_),
    .Y(_12934_));
 sky130_fd_sc_hd__nand2_2 _34578_ (.A(_12931_),
    .B(_12928_),
    .Y(_12935_));
 sky130_fd_sc_hd__nand3_2 _34579_ (.A(_12929_),
    .B(_12925_),
    .C(_12927_),
    .Y(_12936_));
 sky130_fd_sc_hd__nand3_2 _34580_ (.A(_12935_),
    .B(_12936_),
    .C(_12933_),
    .Y(_12937_));
 sky130_fd_sc_hd__nor3_2 _34581_ (.A(_12664_),
    .B(_11832_),
    .C(_11833_),
    .Y(_12938_));
 sky130_vsdinv _34582_ (.A(_12938_),
    .Y(_12939_));
 sky130_fd_sc_hd__o311a_2 _34583_ (.A1(_10884_),
    .A2(_12367_),
    .A3(_11835_),
    .B1(_12117_),
    .C1(_12939_),
    .X(_12940_));
 sky130_fd_sc_hd__o31ai_2 _34584_ (.A1(_10884_),
    .A2(_12367_),
    .A3(_11834_),
    .B1(_12939_),
    .Y(_12941_));
 sky130_fd_sc_hd__nand2_2 _34585_ (.A(_12941_),
    .B(_12116_),
    .Y(_12942_));
 sky130_fd_sc_hd__and2b_2 _34586_ (.A_N(_12940_),
    .B(_12942_),
    .X(_12943_));
 sky130_fd_sc_hd__buf_1 _34587_ (.A(_12943_),
    .X(_12944_));
 sky130_fd_sc_hd__a21oi_2 _34588_ (.A1(_12934_),
    .A2(_12937_),
    .B1(_12944_),
    .Y(_12945_));
 sky130_fd_sc_hd__buf_1 _34589_ (.A(_12943_),
    .X(_12946_));
 sky130_fd_sc_hd__buf_1 _34590_ (.A(_12946_),
    .X(_12947_));
 sky130_fd_sc_hd__nand3_2 _34591_ (.A(_12934_),
    .B(_12947_),
    .C(_12937_),
    .Y(_12948_));
 sky130_vsdinv _34592_ (.A(_12948_),
    .Y(_12949_));
 sky130_fd_sc_hd__o21ai_2 _34593_ (.A1(_12615_),
    .A2(_12612_),
    .B1(_12613_),
    .Y(_12950_));
 sky130_fd_sc_hd__o21bai_2 _34594_ (.A1(_12945_),
    .A2(_12949_),
    .B1_N(_12950_),
    .Y(_12951_));
 sky130_fd_sc_hd__nand3b_2 _34595_ (.A_N(_12945_),
    .B(_12950_),
    .C(_12948_),
    .Y(_12952_));
 sky130_fd_sc_hd__buf_1 _34596_ (.A(_12952_),
    .X(_12953_));
 sky130_fd_sc_hd__o21a_2 _34597_ (.A1(_12672_),
    .A2(_12674_),
    .B1(_12662_),
    .X(_12954_));
 sky130_fd_sc_hd__a21boi_2 _34598_ (.A1(_12951_),
    .A2(_12953_),
    .B1_N(_12954_),
    .Y(_12955_));
 sky130_fd_sc_hd__nand2_2 _34599_ (.A(_12951_),
    .B(_12952_),
    .Y(_12956_));
 sky130_fd_sc_hd__nor2_2 _34600_ (.A(_12954_),
    .B(_12956_),
    .Y(_12957_));
 sky130_fd_sc_hd__nor2_2 _34601_ (.A(_12955_),
    .B(_12957_),
    .Y(_12958_));
 sky130_fd_sc_hd__a21oi_2 _34602_ (.A1(_12902_),
    .A2(_12904_),
    .B1(_12958_),
    .Y(_12959_));
 sky130_fd_sc_hd__nand2_2 _34603_ (.A(_12956_),
    .B(_12954_),
    .Y(_12960_));
 sky130_fd_sc_hd__nand3b_2 _34604_ (.A_N(_12954_),
    .B(_12951_),
    .C(_12953_),
    .Y(_12961_));
 sky130_fd_sc_hd__nand2_2 _34605_ (.A(_12960_),
    .B(_12961_),
    .Y(_12962_));
 sky130_fd_sc_hd__a21oi_2 _34606_ (.A1(_12893_),
    .A2(_12897_),
    .B1(_12900_),
    .Y(_12963_));
 sky130_vsdinv _34607_ (.A(_12904_),
    .Y(_12964_));
 sky130_fd_sc_hd__nor3_2 _34608_ (.A(_12962_),
    .B(_12963_),
    .C(_12964_),
    .Y(_12965_));
 sky130_fd_sc_hd__o21ai_2 _34609_ (.A1(_12691_),
    .A2(_12692_),
    .B1(_12631_),
    .Y(_12966_));
 sky130_fd_sc_hd__o21bai_2 _34610_ (.A1(_12959_),
    .A2(_12965_),
    .B1_N(_12966_),
    .Y(_12967_));
 sky130_fd_sc_hd__nand2_2 _34611_ (.A(_12902_),
    .B(_12903_),
    .Y(_12968_));
 sky130_fd_sc_hd__nand2_2 _34612_ (.A(_12968_),
    .B(_12962_),
    .Y(_12969_));
 sky130_fd_sc_hd__nand3_2 _34613_ (.A(_12958_),
    .B(_12902_),
    .C(_12904_),
    .Y(_12970_));
 sky130_fd_sc_hd__nand3_2 _34614_ (.A(_12969_),
    .B(_12970_),
    .C(_12966_),
    .Y(_12971_));
 sky130_fd_sc_hd__buf_1 _34615_ (.A(_12971_),
    .X(_12972_));
 sky130_fd_sc_hd__a31oi_2 _34616_ (.A1(_12667_),
    .A2(_12442_),
    .A3(_12669_),
    .B1(_12938_),
    .Y(_12973_));
 sky130_fd_sc_hd__nand2_2 _34617_ (.A(_12690_),
    .B(_12681_),
    .Y(_12974_));
 sky130_fd_sc_hd__xnor2_2 _34618_ (.A(_12973_),
    .B(_12974_),
    .Y(_12975_));
 sky130_fd_sc_hd__a21oi_2 _34619_ (.A1(_12967_),
    .A2(_12972_),
    .B1(_12975_),
    .Y(_12976_));
 sky130_vsdinv _34620_ (.A(_12975_),
    .Y(_12977_));
 sky130_fd_sc_hd__a21oi_2 _34621_ (.A1(_12969_),
    .A2(_12970_),
    .B1(_12966_),
    .Y(_12978_));
 sky130_vsdinv _34622_ (.A(_12972_),
    .Y(_12979_));
 sky130_fd_sc_hd__nor3_2 _34623_ (.A(_12977_),
    .B(_12978_),
    .C(_12979_),
    .Y(_12980_));
 sky130_fd_sc_hd__o21ai_2 _34624_ (.A1(_12706_),
    .A2(_12707_),
    .B1(_12701_),
    .Y(_12981_));
 sky130_fd_sc_hd__o21bai_2 _34625_ (.A1(_12976_),
    .A2(_12980_),
    .B1_N(_12981_),
    .Y(_12982_));
 sky130_fd_sc_hd__nand2_2 _34626_ (.A(_12967_),
    .B(_12971_),
    .Y(_12983_));
 sky130_fd_sc_hd__nand2_2 _34627_ (.A(_12983_),
    .B(_12977_),
    .Y(_12984_));
 sky130_fd_sc_hd__nand3_2 _34628_ (.A(_12967_),
    .B(_12975_),
    .C(_12972_),
    .Y(_12985_));
 sky130_fd_sc_hd__nand3_2 _34629_ (.A(_12984_),
    .B(_12985_),
    .C(_12981_),
    .Y(_12986_));
 sky130_fd_sc_hd__a21oi_2 _34630_ (.A1(_12429_),
    .A2(_12425_),
    .B1(_12702_),
    .Y(_12987_));
 sky130_fd_sc_hd__a21oi_2 _34631_ (.A1(_12982_),
    .A2(_12986_),
    .B1(_12987_),
    .Y(_12988_));
 sky130_vsdinv _34632_ (.A(_12987_),
    .Y(_12989_));
 sky130_fd_sc_hd__a21oi_2 _34633_ (.A1(_12984_),
    .A2(_12985_),
    .B1(_12981_),
    .Y(_12990_));
 sky130_vsdinv _34634_ (.A(_12986_),
    .Y(_12991_));
 sky130_fd_sc_hd__nor3_2 _34635_ (.A(_12989_),
    .B(_12990_),
    .C(_12991_),
    .Y(_12992_));
 sky130_fd_sc_hd__o21ai_2 _34636_ (.A1(_12719_),
    .A2(_12720_),
    .B1(_12716_),
    .Y(_12993_));
 sky130_fd_sc_hd__o21bai_2 _34637_ (.A1(_12988_),
    .A2(_12992_),
    .B1_N(_12993_),
    .Y(_12994_));
 sky130_fd_sc_hd__o21bai_2 _34638_ (.A1(_12990_),
    .A2(_12991_),
    .B1_N(_12987_),
    .Y(_12995_));
 sky130_fd_sc_hd__nand3_2 _34639_ (.A(_12982_),
    .B(_12987_),
    .C(_12986_),
    .Y(_12996_));
 sky130_fd_sc_hd__nand3_2 _34640_ (.A(_12995_),
    .B(_12993_),
    .C(_12996_),
    .Y(_12997_));
 sky130_fd_sc_hd__nand2_2 _34641_ (.A(_12994_),
    .B(_12997_),
    .Y(_12998_));
 sky130_vsdinv _34642_ (.A(_12730_),
    .Y(_12999_));
 sky130_fd_sc_hd__a21oi_2 _34643_ (.A1(_12734_),
    .A2(_12727_),
    .B1(_12999_),
    .Y(_13000_));
 sky130_fd_sc_hd__xor2_2 _34644_ (.A(_12998_),
    .B(_13000_),
    .X(_02658_));
 sky130_fd_sc_hd__nand2_2 _34645_ (.A(_18694_),
    .B(_19257_),
    .Y(_13001_));
 sky130_fd_sc_hd__nand3b_2 _34646_ (.A_N(_13001_),
    .B(_11599_),
    .C(_19262_),
    .Y(_13002_));
 sky130_fd_sc_hd__o21ai_2 _34647_ (.A1(_05841_),
    .A2(_16969_),
    .B1(_13001_),
    .Y(_13003_));
 sky130_fd_sc_hd__and2_2 _34648_ (.A(_11326_),
    .B(_07382_),
    .X(_13004_));
 sky130_fd_sc_hd__a21o_2 _34649_ (.A1(_13002_),
    .A2(_13003_),
    .B1(_13004_),
    .X(_13005_));
 sky130_fd_sc_hd__nand3_2 _34650_ (.A(_13002_),
    .B(_13004_),
    .C(_13003_),
    .Y(_13006_));
 sky130_fd_sc_hd__nand2_2 _34651_ (.A(_12740_),
    .B(_12736_),
    .Y(_13007_));
 sky130_fd_sc_hd__a21o_2 _34652_ (.A1(_13005_),
    .A2(_13006_),
    .B1(_13007_),
    .X(_13008_));
 sky130_fd_sc_hd__nand3_2 _34653_ (.A(_13007_),
    .B(_13005_),
    .C(_13006_),
    .Y(_13009_));
 sky130_fd_sc_hd__and2_2 _34654_ (.A(_09319_),
    .B(_06350_),
    .X(_13010_));
 sky130_fd_sc_hd__a22oi_2 _34655_ (.A1(_10260_),
    .A2(_06588_),
    .B1(_10253_),
    .B2(_07264_),
    .Y(_13011_));
 sky130_fd_sc_hd__and4_2 _34656_ (.A(_10260_),
    .B(_10686_),
    .C(_06728_),
    .D(_07515_),
    .X(_13012_));
 sky130_fd_sc_hd__nor2_2 _34657_ (.A(_13011_),
    .B(_13012_),
    .Y(_13013_));
 sky130_fd_sc_hd__xor2_2 _34658_ (.A(_13010_),
    .B(_13013_),
    .X(_13014_));
 sky130_fd_sc_hd__a21oi_2 _34659_ (.A1(_13008_),
    .A2(_13009_),
    .B1(_13014_),
    .Y(_13015_));
 sky130_fd_sc_hd__nand3_2 _34660_ (.A(_13008_),
    .B(_13014_),
    .C(_13009_),
    .Y(_13016_));
 sky130_vsdinv _34661_ (.A(_13016_),
    .Y(_13017_));
 sky130_fd_sc_hd__nand2_2 _34662_ (.A(_12757_),
    .B(_12745_),
    .Y(_13018_));
 sky130_fd_sc_hd__o21bai_2 _34663_ (.A1(_13015_),
    .A2(_13017_),
    .B1_N(_13018_),
    .Y(_13019_));
 sky130_fd_sc_hd__a21o_2 _34664_ (.A1(_13008_),
    .A2(_13009_),
    .B1(_13014_),
    .X(_13020_));
 sky130_fd_sc_hd__nand3_2 _34665_ (.A(_13020_),
    .B(_13018_),
    .C(_13016_),
    .Y(_13021_));
 sky130_fd_sc_hd__nand2_2 _34666_ (.A(_13019_),
    .B(_13021_),
    .Y(_13022_));
 sky130_fd_sc_hd__nand2_2 _34667_ (.A(_11634_),
    .B(_07688_),
    .Y(_13023_));
 sky130_fd_sc_hd__nand2_2 _34668_ (.A(_10231_),
    .B(_07306_),
    .Y(_13024_));
 sky130_fd_sc_hd__xor2_2 _34669_ (.A(_13023_),
    .B(_13024_),
    .X(_13025_));
 sky130_fd_sc_hd__buf_1 _34670_ (.A(_10703_),
    .X(_13026_));
 sky130_fd_sc_hd__nand3_2 _34671_ (.A(_13025_),
    .B(_13026_),
    .C(_10775_),
    .Y(_13027_));
 sky130_fd_sc_hd__xnor2_2 _34672_ (.A(_13023_),
    .B(_13024_),
    .Y(_13028_));
 sky130_fd_sc_hd__o21ai_2 _34673_ (.A1(_11036_),
    .A2(_19218_),
    .B1(_13028_),
    .Y(_13029_));
 sky130_fd_sc_hd__a21oi_2 _34674_ (.A1(_12750_),
    .A2(_12749_),
    .B1(_12748_),
    .Y(_13030_));
 sky130_vsdinv _34675_ (.A(_13030_),
    .Y(_13031_));
 sky130_fd_sc_hd__a21o_2 _34676_ (.A1(_13027_),
    .A2(_13029_),
    .B1(_13031_),
    .X(_13032_));
 sky130_fd_sc_hd__nand3_2 _34677_ (.A(_13027_),
    .B(_13029_),
    .C(_13031_),
    .Y(_13033_));
 sky130_fd_sc_hd__a21boi_2 _34678_ (.A1(_12764_),
    .A2(_12768_),
    .B1_N(_12766_),
    .Y(_13034_));
 sky130_fd_sc_hd__a21bo_2 _34679_ (.A1(_13032_),
    .A2(_13033_),
    .B1_N(_13034_),
    .X(_13035_));
 sky130_fd_sc_hd__nand3b_2 _34680_ (.A_N(_13034_),
    .B(_13032_),
    .C(_13033_),
    .Y(_13036_));
 sky130_fd_sc_hd__nand2_2 _34681_ (.A(_13035_),
    .B(_13036_),
    .Y(_13037_));
 sky130_fd_sc_hd__nand2_2 _34682_ (.A(_13022_),
    .B(_13037_),
    .Y(_13038_));
 sky130_fd_sc_hd__nand3b_2 _34683_ (.A_N(_13037_),
    .B(_13021_),
    .C(_13019_),
    .Y(_13039_));
 sky130_fd_sc_hd__nand2_2 _34684_ (.A(_13038_),
    .B(_13039_),
    .Y(_13040_));
 sky130_fd_sc_hd__o21ai_2 _34685_ (.A1(_12777_),
    .A2(_12780_),
    .B1(_12763_),
    .Y(_13041_));
 sky130_vsdinv _34686_ (.A(_13041_),
    .Y(_13042_));
 sky130_fd_sc_hd__nand2_2 _34687_ (.A(_13040_),
    .B(_13042_),
    .Y(_13043_));
 sky130_fd_sc_hd__nand3_2 _34688_ (.A(_13038_),
    .B(_13039_),
    .C(_13041_),
    .Y(_13044_));
 sky130_fd_sc_hd__buf_1 _34689_ (.A(_13044_),
    .X(_13045_));
 sky130_fd_sc_hd__nand2_2 _34690_ (.A(_10186_),
    .B(_07605_),
    .Y(_13046_));
 sky130_fd_sc_hd__nand2_2 _34691_ (.A(_08224_),
    .B(_07748_),
    .Y(_13047_));
 sky130_fd_sc_hd__nand2_2 _34692_ (.A(_13046_),
    .B(_13047_),
    .Y(_13048_));
 sky130_fd_sc_hd__nand3b_2 _34693_ (.A_N(_13046_),
    .B(_12791_),
    .C(_08301_),
    .Y(_13049_));
 sky130_fd_sc_hd__buf_1 _34694_ (.A(_18759_),
    .X(_13050_));
 sky130_fd_sc_hd__o2bb2ai_2 _34695_ (.A1_N(_13048_),
    .A2_N(_13049_),
    .B1(_13050_),
    .B2(_19205_),
    .Y(_13051_));
 sky130_fd_sc_hd__and2_2 _34696_ (.A(_08235_),
    .B(_08302_),
    .X(_13052_));
 sky130_fd_sc_hd__nand3_2 _34697_ (.A(_13049_),
    .B(_13048_),
    .C(_13052_),
    .Y(_13053_));
 sky130_fd_sc_hd__nor2_2 _34698_ (.A(_12790_),
    .B(_12795_),
    .Y(_13054_));
 sky130_fd_sc_hd__a21oi_2 _34699_ (.A1(_12796_),
    .A2(_12793_),
    .B1(_13054_),
    .Y(_13055_));
 sky130_vsdinv _34700_ (.A(_13055_),
    .Y(_13056_));
 sky130_fd_sc_hd__a21o_2 _34701_ (.A1(_13051_),
    .A2(_13053_),
    .B1(_13056_),
    .X(_13057_));
 sky130_fd_sc_hd__nand3_2 _34702_ (.A(_13051_),
    .B(_13056_),
    .C(_13053_),
    .Y(_13058_));
 sky130_fd_sc_hd__and2_2 _34703_ (.A(_10436_),
    .B(_08826_),
    .X(_13059_));
 sky130_fd_sc_hd__nand2_2 _34704_ (.A(_08218_),
    .B(_08549_),
    .Y(_13060_));
 sky130_fd_sc_hd__nand2_2 _34705_ (.A(_10207_),
    .B(_11136_),
    .Y(_13061_));
 sky130_fd_sc_hd__xnor2_2 _34706_ (.A(_13060_),
    .B(_13061_),
    .Y(_13062_));
 sky130_fd_sc_hd__xnor2_2 _34707_ (.A(_13059_),
    .B(_13062_),
    .Y(_13063_));
 sky130_fd_sc_hd__a21oi_2 _34708_ (.A1(_13057_),
    .A2(_13058_),
    .B1(_13063_),
    .Y(_13064_));
 sky130_fd_sc_hd__nand3_2 _34709_ (.A(_13063_),
    .B(_13057_),
    .C(_13058_),
    .Y(_13065_));
 sky130_vsdinv _34710_ (.A(_13065_),
    .Y(_13066_));
 sky130_fd_sc_hd__nand2_2 _34711_ (.A(_12776_),
    .B(_12772_),
    .Y(_13067_));
 sky130_fd_sc_hd__o21bai_2 _34712_ (.A1(_13064_),
    .A2(_13066_),
    .B1_N(_13067_),
    .Y(_13068_));
 sky130_fd_sc_hd__nand3b_2 _34713_ (.A_N(_13064_),
    .B(_13067_),
    .C(_13065_),
    .Y(_13069_));
 sky130_fd_sc_hd__a21boi_2 _34714_ (.A1(_12809_),
    .A2(_12801_),
    .B1_N(_12799_),
    .Y(_13070_));
 sky130_vsdinv _34715_ (.A(_13070_),
    .Y(_13071_));
 sky130_fd_sc_hd__a21o_2 _34716_ (.A1(_13068_),
    .A2(_13069_),
    .B1(_13071_),
    .X(_13072_));
 sky130_fd_sc_hd__nand3_2 _34717_ (.A(_13068_),
    .B(_13071_),
    .C(_13069_),
    .Y(_13073_));
 sky130_fd_sc_hd__and2_2 _34718_ (.A(_13072_),
    .B(_13073_),
    .X(_13074_));
 sky130_fd_sc_hd__a21oi_2 _34719_ (.A1(_13043_),
    .A2(_13045_),
    .B1(_13074_),
    .Y(_13075_));
 sky130_fd_sc_hd__nand2_2 _34720_ (.A(_13072_),
    .B(_13073_),
    .Y(_13076_));
 sky130_fd_sc_hd__a21oi_2 _34721_ (.A1(_13038_),
    .A2(_13039_),
    .B1(_13041_),
    .Y(_13077_));
 sky130_fd_sc_hd__nor3b_2 _34722_ (.A(_13076_),
    .B(_13077_),
    .C_N(_13045_),
    .Y(_13078_));
 sky130_fd_sc_hd__o21ai_2 _34723_ (.A1(_12826_),
    .A2(_12827_),
    .B1(_12787_),
    .Y(_13079_));
 sky130_fd_sc_hd__o21bai_2 _34724_ (.A1(_13075_),
    .A2(_13078_),
    .B1_N(_13079_),
    .Y(_13080_));
 sky130_fd_sc_hd__nand2_2 _34725_ (.A(_13043_),
    .B(_13044_),
    .Y(_13081_));
 sky130_fd_sc_hd__nand2_2 _34726_ (.A(_13081_),
    .B(_13076_),
    .Y(_13082_));
 sky130_fd_sc_hd__nand3_2 _34727_ (.A(_13074_),
    .B(_13045_),
    .C(_13043_),
    .Y(_13083_));
 sky130_fd_sc_hd__nand3_2 _34728_ (.A(_13082_),
    .B(_13083_),
    .C(_13079_),
    .Y(_13084_));
 sky130_fd_sc_hd__buf_1 _34729_ (.A(_13084_),
    .X(_13085_));
 sky130_fd_sc_hd__nand2_2 _34730_ (.A(_07469_),
    .B(_10574_),
    .Y(_13086_));
 sky130_fd_sc_hd__nand2_2 _34731_ (.A(_08908_),
    .B(_19172_),
    .Y(_13087_));
 sky130_fd_sc_hd__xor2_2 _34732_ (.A(_13086_),
    .B(_13087_),
    .X(_13088_));
 sky130_fd_sc_hd__buf_1 _34733_ (.A(_11409_),
    .X(_13089_));
 sky130_fd_sc_hd__nand3_2 _34734_ (.A(_13088_),
    .B(_13089_),
    .C(_12859_),
    .Y(_13090_));
 sky130_fd_sc_hd__xnor2_2 _34735_ (.A(_13086_),
    .B(_13087_),
    .Y(_13091_));
 sky130_fd_sc_hd__o21ai_2 _34736_ (.A1(_07400_),
    .A2(_19168_),
    .B1(_13091_),
    .Y(_13092_));
 sky130_fd_sc_hd__a21boi_2 _34737_ (.A1(_12802_),
    .A2(_12807_),
    .B1_N(_12804_),
    .Y(_13093_));
 sky130_fd_sc_hd__a21bo_2 _34738_ (.A1(_13090_),
    .A2(_13092_),
    .B1_N(_13093_),
    .X(_13094_));
 sky130_fd_sc_hd__nand3b_2 _34739_ (.A_N(_13093_),
    .B(_13090_),
    .C(_13092_),
    .Y(_13095_));
 sky130_fd_sc_hd__a21boi_2 _34740_ (.A1(_12837_),
    .A2(_12843_),
    .B1_N(_12840_),
    .Y(_13096_));
 sky130_vsdinv _34741_ (.A(_13096_),
    .Y(_13097_));
 sky130_fd_sc_hd__a21oi_2 _34742_ (.A1(_13094_),
    .A2(_13095_),
    .B1(_13097_),
    .Y(_13098_));
 sky130_fd_sc_hd__nand3_2 _34743_ (.A(_13094_),
    .B(_13097_),
    .C(_13095_),
    .Y(_13099_));
 sky130_vsdinv _34744_ (.A(_13099_),
    .Y(_13100_));
 sky130_fd_sc_hd__nand2_2 _34745_ (.A(_12855_),
    .B(_12851_),
    .Y(_13101_));
 sky130_fd_sc_hd__o21bai_2 _34746_ (.A1(_13098_),
    .A2(_13100_),
    .B1_N(_13101_),
    .Y(_13102_));
 sky130_fd_sc_hd__nand3b_2 _34747_ (.A_N(_13098_),
    .B(_13099_),
    .C(_13101_),
    .Y(_13103_));
 sky130_fd_sc_hd__nand2_2 _34748_ (.A(_13102_),
    .B(_13103_),
    .Y(_13104_));
 sky130_fd_sc_hd__and2_2 _34749_ (.A(_06816_),
    .B(_12905_),
    .X(_13105_));
 sky130_fd_sc_hd__nand2_2 _34750_ (.A(_06671_),
    .B(_10894_),
    .Y(_13106_));
 sky130_fd_sc_hd__nand2_2 _34751_ (.A(_06674_),
    .B(_11198_),
    .Y(_13107_));
 sky130_fd_sc_hd__xnor2_2 _34752_ (.A(_13106_),
    .B(_13107_),
    .Y(_13108_));
 sky130_fd_sc_hd__xor2_2 _34753_ (.A(_13105_),
    .B(_13108_),
    .X(_13109_));
 sky130_fd_sc_hd__nand2_2 _34754_ (.A(_18798_),
    .B(_11221_),
    .Y(_13110_));
 sky130_fd_sc_hd__nand2_2 _34755_ (.A(_08688_),
    .B(_10533_),
    .Y(_13111_));
 sky130_fd_sc_hd__xor2_2 _34756_ (.A(_13110_),
    .B(_13111_),
    .X(_13112_));
 sky130_fd_sc_hd__buf_1 _34757_ (.A(_10551_),
    .X(_13113_));
 sky130_fd_sc_hd__and2_2 _34758_ (.A(_06551_),
    .B(_13113_),
    .X(_13114_));
 sky130_fd_sc_hd__nand2_2 _34759_ (.A(_13112_),
    .B(_13114_),
    .Y(_13115_));
 sky130_fd_sc_hd__xnor2_2 _34760_ (.A(_13110_),
    .B(_13111_),
    .Y(_13116_));
 sky130_fd_sc_hd__o21ai_2 _34761_ (.A1(_06692_),
    .A2(_19152_),
    .B1(_13116_),
    .Y(_13117_));
 sky130_fd_sc_hd__nand2_2 _34762_ (.A(_12867_),
    .B(_12864_),
    .Y(_13118_));
 sky130_fd_sc_hd__a21oi_2 _34763_ (.A1(_13115_),
    .A2(_13117_),
    .B1(_13118_),
    .Y(_13119_));
 sky130_fd_sc_hd__nand3_2 _34764_ (.A(_13115_),
    .B(_13117_),
    .C(_13118_),
    .Y(_13120_));
 sky130_fd_sc_hd__and2b_2 _34765_ (.A_N(_13119_),
    .B(_13120_),
    .X(_13121_));
 sky130_fd_sc_hd__xor2_2 _34766_ (.A(_13109_),
    .B(_13121_),
    .X(_13122_));
 sky130_fd_sc_hd__nand2_2 _34767_ (.A(_13104_),
    .B(_13122_),
    .Y(_13123_));
 sky130_vsdinv _34768_ (.A(_13109_),
    .Y(_13124_));
 sky130_fd_sc_hd__xor2_2 _34769_ (.A(_13124_),
    .B(_13121_),
    .X(_13125_));
 sky130_fd_sc_hd__nand3_2 _34770_ (.A(_13125_),
    .B(_13103_),
    .C(_13102_),
    .Y(_13126_));
 sky130_fd_sc_hd__o21ai_2 _34771_ (.A1(_12816_),
    .A2(_12823_),
    .B1(_12814_),
    .Y(_13127_));
 sky130_fd_sc_hd__a21oi_2 _34772_ (.A1(_13123_),
    .A2(_13126_),
    .B1(_13127_),
    .Y(_13128_));
 sky130_fd_sc_hd__nand3_2 _34773_ (.A(_13123_),
    .B(_13126_),
    .C(_13127_),
    .Y(_13129_));
 sky130_vsdinv _34774_ (.A(_13129_),
    .Y(_13130_));
 sky130_fd_sc_hd__o21a_2 _34775_ (.A1(_12879_),
    .A2(_12881_),
    .B1(_12858_),
    .X(_13131_));
 sky130_fd_sc_hd__o21ai_2 _34776_ (.A1(_13128_),
    .A2(_13130_),
    .B1(_13131_),
    .Y(_13132_));
 sky130_fd_sc_hd__a21o_2 _34777_ (.A1(_13123_),
    .A2(_13126_),
    .B1(_13127_),
    .X(_13133_));
 sky130_fd_sc_hd__nand3b_2 _34778_ (.A_N(_13131_),
    .B(_13133_),
    .C(_13129_),
    .Y(_13134_));
 sky130_fd_sc_hd__nand2_2 _34779_ (.A(_13132_),
    .B(_13134_),
    .Y(_13135_));
 sky130_fd_sc_hd__buf_1 _34780_ (.A(_13135_),
    .X(_13136_));
 sky130_fd_sc_hd__a21boi_2 _34781_ (.A1(_13080_),
    .A2(_13085_),
    .B1_N(_13136_),
    .Y(_13137_));
 sky130_fd_sc_hd__a21oi_2 _34782_ (.A1(_13082_),
    .A2(_13083_),
    .B1(_13079_),
    .Y(_13138_));
 sky130_vsdinv _34783_ (.A(_13085_),
    .Y(_13139_));
 sky130_fd_sc_hd__nor3_2 _34784_ (.A(_13136_),
    .B(_13138_),
    .C(_13139_),
    .Y(_13140_));
 sky130_fd_sc_hd__a21oi_2 _34785_ (.A1(_12832_),
    .A2(_12833_),
    .B1(_12830_),
    .Y(_13141_));
 sky130_fd_sc_hd__o21ai_2 _34786_ (.A1(_13141_),
    .A2(_12892_),
    .B1(_12834_),
    .Y(_13142_));
 sky130_fd_sc_hd__o21bai_2 _34787_ (.A1(_13137_),
    .A2(_13140_),
    .B1_N(_13142_),
    .Y(_13143_));
 sky130_fd_sc_hd__nand2_2 _34788_ (.A(_13080_),
    .B(_13084_),
    .Y(_13144_));
 sky130_fd_sc_hd__nand2_2 _34789_ (.A(_13144_),
    .B(_13136_),
    .Y(_13145_));
 sky130_fd_sc_hd__nand3b_2 _34790_ (.A_N(_13135_),
    .B(_13080_),
    .C(_13085_),
    .Y(_13146_));
 sky130_fd_sc_hd__nand3_2 _34791_ (.A(_13145_),
    .B(_13146_),
    .C(_13142_),
    .Y(_13147_));
 sky130_fd_sc_hd__buf_1 _34792_ (.A(_13147_),
    .X(_13148_));
 sky130_fd_sc_hd__nand2_2 _34793_ (.A(_12873_),
    .B(_12874_),
    .Y(_13149_));
 sky130_fd_sc_hd__nor2_2 _34794_ (.A(_12873_),
    .B(_12874_),
    .Y(_13150_));
 sky130_fd_sc_hd__a21oi_2 _34795_ (.A1(_13149_),
    .A2(_12872_),
    .B1(_13150_),
    .Y(_13151_));
 sky130_fd_sc_hd__nand2_2 _34796_ (.A(_10880_),
    .B(_18827_),
    .Y(_13152_));
 sky130_fd_sc_hd__nand2_2 _34797_ (.A(_12908_),
    .B(_13152_),
    .Y(_13153_));
 sky130_fd_sc_hd__nand3_2 _34798_ (.A(_10880_),
    .B(_18827_),
    .C(_05766_),
    .Y(_13154_));
 sky130_fd_sc_hd__and3_2 _34799_ (.A(_13153_),
    .B(_12636_),
    .C(_13154_),
    .X(_13155_));
 sky130_fd_sc_hd__buf_1 _34800_ (.A(_13155_),
    .X(_13156_));
 sky130_vsdinv _34801_ (.A(_13156_),
    .Y(_13157_));
 sky130_fd_sc_hd__a21oi_2 _34802_ (.A1(_13153_),
    .A2(_13154_),
    .B1(_12636_),
    .Y(_13158_));
 sky130_vsdinv _34803_ (.A(_13158_),
    .Y(_13159_));
 sky130_fd_sc_hd__nand3b_2 _34804_ (.A_N(_13151_),
    .B(_13157_),
    .C(_13159_),
    .Y(_13160_));
 sky130_fd_sc_hd__buf_1 _34805_ (.A(_13158_),
    .X(_13161_));
 sky130_fd_sc_hd__buf_1 _34806_ (.A(_13161_),
    .X(_13162_));
 sky130_fd_sc_hd__buf_1 _34807_ (.A(_13156_),
    .X(_13163_));
 sky130_fd_sc_hd__o21ai_2 _34808_ (.A1(_13162_),
    .A2(_13163_),
    .B1(_13151_),
    .Y(_13164_));
 sky130_fd_sc_hd__o31a_2 _34809_ (.A1(_11487_),
    .A2(_06114_),
    .A3(_12906_),
    .B1(_12910_),
    .X(_13165_));
 sky130_vsdinv _34810_ (.A(_13165_),
    .Y(_13166_));
 sky130_fd_sc_hd__a21oi_2 _34811_ (.A1(_13160_),
    .A2(_13164_),
    .B1(_13166_),
    .Y(_13167_));
 sky130_fd_sc_hd__and3_2 _34812_ (.A(_13160_),
    .B(_13166_),
    .C(_13164_),
    .X(_13168_));
 sky130_fd_sc_hd__nor2_2 _34813_ (.A(_13167_),
    .B(_13168_),
    .Y(_13169_));
 sky130_fd_sc_hd__nand2_2 _34814_ (.A(_12878_),
    .B(_12869_),
    .Y(_13170_));
 sky130_fd_sc_hd__nand2_2 _34815_ (.A(_13169_),
    .B(_13170_),
    .Y(_13171_));
 sky130_fd_sc_hd__o211ai_2 _34816_ (.A1(_13167_),
    .A2(_13168_),
    .B1(_12869_),
    .C1(_12878_),
    .Y(_13172_));
 sky130_fd_sc_hd__nand2_2 _34817_ (.A(_13171_),
    .B(_13172_),
    .Y(_13173_));
 sky130_vsdinv _34818_ (.A(_12920_),
    .Y(_13174_));
 sky130_fd_sc_hd__a21oi_2 _34819_ (.A1(_12917_),
    .A2(_12919_),
    .B1(_13174_),
    .Y(_13175_));
 sky130_fd_sc_hd__nand2_2 _34820_ (.A(_13173_),
    .B(_13175_),
    .Y(_13176_));
 sky130_fd_sc_hd__nand3b_2 _34821_ (.A_N(_13175_),
    .B(_13171_),
    .C(_13172_),
    .Y(_13177_));
 sky130_fd_sc_hd__nand2_2 _34822_ (.A(_13176_),
    .B(_13177_),
    .Y(_13178_));
 sky130_fd_sc_hd__a21boi_2 _34823_ (.A1(_12929_),
    .A2(_12925_),
    .B1_N(_12927_),
    .Y(_13179_));
 sky130_fd_sc_hd__nand2_2 _34824_ (.A(_13178_),
    .B(_13179_),
    .Y(_13180_));
 sky130_fd_sc_hd__nand2_2 _34825_ (.A(_12936_),
    .B(_12927_),
    .Y(_13181_));
 sky130_fd_sc_hd__nand3_2 _34826_ (.A(_13181_),
    .B(_13177_),
    .C(_13176_),
    .Y(_13182_));
 sky130_fd_sc_hd__buf_1 _34827_ (.A(_12946_),
    .X(_13183_));
 sky130_fd_sc_hd__buf_1 _34828_ (.A(_13183_),
    .X(_13184_));
 sky130_fd_sc_hd__a21oi_2 _34829_ (.A1(_13180_),
    .A2(_13182_),
    .B1(_13184_),
    .Y(_13185_));
 sky130_fd_sc_hd__nand3_2 _34830_ (.A(_13180_),
    .B(_12947_),
    .C(_13182_),
    .Y(_13186_));
 sky130_vsdinv _34831_ (.A(_13186_),
    .Y(_13187_));
 sky130_fd_sc_hd__a21boi_2 _34832_ (.A1(_12884_),
    .A2(_12889_),
    .B1_N(_12887_),
    .Y(_13188_));
 sky130_fd_sc_hd__o21ai_2 _34833_ (.A1(_13185_),
    .A2(_13187_),
    .B1(_13188_),
    .Y(_13189_));
 sky130_fd_sc_hd__nand2_2 _34834_ (.A(_12891_),
    .B(_12887_),
    .Y(_13190_));
 sky130_fd_sc_hd__a21o_2 _34835_ (.A1(_13180_),
    .A2(_13182_),
    .B1(_12947_),
    .X(_13191_));
 sky130_fd_sc_hd__nand3_2 _34836_ (.A(_13190_),
    .B(_13186_),
    .C(_13191_),
    .Y(_13192_));
 sky130_fd_sc_hd__buf_1 _34837_ (.A(_12946_),
    .X(_13193_));
 sky130_fd_sc_hd__buf_1 _34838_ (.A(_13193_),
    .X(_13194_));
 sky130_fd_sc_hd__a21boi_2 _34839_ (.A1(_12934_),
    .A2(_13194_),
    .B1_N(_12937_),
    .Y(_13195_));
 sky130_fd_sc_hd__a21bo_2 _34840_ (.A1(_13189_),
    .A2(_13192_),
    .B1_N(_13195_),
    .X(_13196_));
 sky130_fd_sc_hd__nand3b_2 _34841_ (.A_N(_13195_),
    .B(_13189_),
    .C(_13192_),
    .Y(_13197_));
 sky130_fd_sc_hd__and2_2 _34842_ (.A(_13196_),
    .B(_13197_),
    .X(_13198_));
 sky130_fd_sc_hd__a21oi_2 _34843_ (.A1(_13143_),
    .A2(_13148_),
    .B1(_13198_),
    .Y(_13199_));
 sky130_fd_sc_hd__nand2_2 _34844_ (.A(_13196_),
    .B(_13197_),
    .Y(_13200_));
 sky130_fd_sc_hd__a21oi_2 _34845_ (.A1(_13145_),
    .A2(_13146_),
    .B1(_13142_),
    .Y(_13201_));
 sky130_vsdinv _34846_ (.A(_13148_),
    .Y(_13202_));
 sky130_fd_sc_hd__nor3_2 _34847_ (.A(_13200_),
    .B(_13201_),
    .C(_13202_),
    .Y(_13203_));
 sky130_fd_sc_hd__o21ai_2 _34848_ (.A1(_12962_),
    .A2(_12963_),
    .B1(_12904_),
    .Y(_13204_));
 sky130_fd_sc_hd__o21bai_2 _34849_ (.A1(_13199_),
    .A2(_13203_),
    .B1_N(_13204_),
    .Y(_13205_));
 sky130_fd_sc_hd__nand2_2 _34850_ (.A(_13143_),
    .B(_13147_),
    .Y(_13206_));
 sky130_fd_sc_hd__nand2_2 _34851_ (.A(_13206_),
    .B(_13200_),
    .Y(_13207_));
 sky130_fd_sc_hd__nand3_2 _34852_ (.A(_13198_),
    .B(_13148_),
    .C(_13143_),
    .Y(_13208_));
 sky130_fd_sc_hd__nand3_2 _34853_ (.A(_13207_),
    .B(_13208_),
    .C(_13204_),
    .Y(_13209_));
 sky130_fd_sc_hd__buf_1 _34854_ (.A(_13209_),
    .X(_13210_));
 sky130_fd_sc_hd__nor2_2 _34855_ (.A(_12938_),
    .B(_12940_),
    .Y(_13211_));
 sky130_vsdinv _34856_ (.A(_13211_),
    .Y(_13212_));
 sky130_fd_sc_hd__buf_1 _34857_ (.A(_13212_),
    .X(_13213_));
 sky130_fd_sc_hd__nand2_2 _34858_ (.A(_12961_),
    .B(_12953_),
    .Y(_13214_));
 sky130_fd_sc_hd__xor2_2 _34859_ (.A(_13213_),
    .B(_13214_),
    .X(_13215_));
 sky130_fd_sc_hd__a21oi_2 _34860_ (.A1(_13205_),
    .A2(_13210_),
    .B1(_13215_),
    .Y(_13216_));
 sky130_vsdinv _34861_ (.A(_13215_),
    .Y(_13217_));
 sky130_fd_sc_hd__a21oi_2 _34862_ (.A1(_13207_),
    .A2(_13208_),
    .B1(_13204_),
    .Y(_13218_));
 sky130_vsdinv _34863_ (.A(_13210_),
    .Y(_13219_));
 sky130_fd_sc_hd__nor3_2 _34864_ (.A(_13217_),
    .B(_13218_),
    .C(_13219_),
    .Y(_13220_));
 sky130_fd_sc_hd__o21ai_2 _34865_ (.A1(_12977_),
    .A2(_12978_),
    .B1(_12972_),
    .Y(_13221_));
 sky130_fd_sc_hd__o21bai_2 _34866_ (.A1(_13216_),
    .A2(_13220_),
    .B1_N(_13221_),
    .Y(_13222_));
 sky130_fd_sc_hd__nand2_2 _34867_ (.A(_13205_),
    .B(_13209_),
    .Y(_13223_));
 sky130_fd_sc_hd__nand2_2 _34868_ (.A(_13223_),
    .B(_13217_),
    .Y(_13224_));
 sky130_fd_sc_hd__nand3_2 _34869_ (.A(_13205_),
    .B(_13215_),
    .C(_13210_),
    .Y(_13225_));
 sky130_fd_sc_hd__nand3_2 _34870_ (.A(_13224_),
    .B(_13221_),
    .C(_13225_),
    .Y(_13226_));
 sky130_fd_sc_hd__a21oi_2 _34871_ (.A1(_12690_),
    .A2(_12681_),
    .B1(_12973_),
    .Y(_13227_));
 sky130_fd_sc_hd__a21oi_2 _34872_ (.A1(_13222_),
    .A2(_13226_),
    .B1(_13227_),
    .Y(_13228_));
 sky130_vsdinv _34873_ (.A(_13227_),
    .Y(_13229_));
 sky130_fd_sc_hd__a21oi_2 _34874_ (.A1(_13224_),
    .A2(_13225_),
    .B1(_13221_),
    .Y(_13230_));
 sky130_vsdinv _34875_ (.A(_13226_),
    .Y(_13231_));
 sky130_fd_sc_hd__nor3_2 _34876_ (.A(_13229_),
    .B(_13230_),
    .C(_13231_),
    .Y(_13232_));
 sky130_fd_sc_hd__o21ai_2 _34877_ (.A1(_12989_),
    .A2(_12990_),
    .B1(_12986_),
    .Y(_13233_));
 sky130_fd_sc_hd__o21bai_2 _34878_ (.A1(_13228_),
    .A2(_13232_),
    .B1_N(_13233_),
    .Y(_13234_));
 sky130_fd_sc_hd__o21bai_2 _34879_ (.A1(_13230_),
    .A2(_13231_),
    .B1_N(_13227_),
    .Y(_13235_));
 sky130_fd_sc_hd__nand3_2 _34880_ (.A(_13222_),
    .B(_13227_),
    .C(_13226_),
    .Y(_13236_));
 sky130_fd_sc_hd__nand3_2 _34881_ (.A(_13235_),
    .B(_13233_),
    .C(_13236_),
    .Y(_13237_));
 sky130_fd_sc_hd__nand2_2 _34882_ (.A(_13234_),
    .B(_13237_),
    .Y(_13238_));
 sky130_fd_sc_hd__nor2_2 _34883_ (.A(_12176_),
    .B(_12463_),
    .Y(_13239_));
 sky130_fd_sc_hd__nand2_2 _34884_ (.A(_12727_),
    .B(_12730_),
    .Y(_13240_));
 sky130_fd_sc_hd__nor2_2 _34885_ (.A(_13240_),
    .B(_12998_),
    .Y(_13241_));
 sky130_fd_sc_hd__nand2_2 _34886_ (.A(_13239_),
    .B(_13241_),
    .Y(_13242_));
 sky130_fd_sc_hd__nor2_2 _34887_ (.A(_13242_),
    .B(_12177_),
    .Y(_13243_));
 sky130_fd_sc_hd__a21oi_2 _34888_ (.A1(_12179_),
    .A2(_12181_),
    .B1(_13242_),
    .Y(_13244_));
 sky130_fd_sc_hd__a21boi_2 _34889_ (.A1(_12999_),
    .A2(_12994_),
    .B1_N(_12997_),
    .Y(_13245_));
 sky130_fd_sc_hd__o31ai_2 _34890_ (.A1(_13240_),
    .A2(_12998_),
    .A3(_12733_),
    .B1(_13245_),
    .Y(_13246_));
 sky130_fd_sc_hd__a211oi_2 _34891_ (.A1(_10993_),
    .A2(_13243_),
    .B1(_13244_),
    .C1(_13246_),
    .Y(_13247_));
 sky130_fd_sc_hd__xor2_2 _34892_ (.A(_13238_),
    .B(_13247_),
    .X(_02659_));
 sky130_fd_sc_hd__nand2_2 _34893_ (.A(_10480_),
    .B(_06067_),
    .Y(_13248_));
 sky130_fd_sc_hd__nand3b_2 _34894_ (.A_N(_13248_),
    .B(_10996_),
    .C(_19258_),
    .Y(_13249_));
 sky130_fd_sc_hd__o21ai_2 _34895_ (.A1(_05958_),
    .A2(_11004_),
    .B1(_13248_),
    .Y(_13250_));
 sky130_fd_sc_hd__and2_2 _34896_ (.A(_18703_),
    .B(_08905_),
    .X(_13251_));
 sky130_fd_sc_hd__a21o_2 _34897_ (.A1(_13249_),
    .A2(_13250_),
    .B1(_13251_),
    .X(_13252_));
 sky130_fd_sc_hd__nand3_2 _34898_ (.A(_13249_),
    .B(_13251_),
    .C(_13250_),
    .Y(_13253_));
 sky130_fd_sc_hd__nand2_2 _34899_ (.A(_13006_),
    .B(_13002_),
    .Y(_13254_));
 sky130_fd_sc_hd__a21o_2 _34900_ (.A1(_13252_),
    .A2(_13253_),
    .B1(_13254_),
    .X(_13255_));
 sky130_fd_sc_hd__nand3_2 _34901_ (.A(_13254_),
    .B(_13252_),
    .C(_13253_),
    .Y(_13256_));
 sky130_fd_sc_hd__nand2_2 _34902_ (.A(_10260_),
    .B(_07264_),
    .Y(_13257_));
 sky130_fd_sc_hd__nand2_2 _34903_ (.A(_11015_),
    .B(_06350_),
    .Y(_13258_));
 sky130_fd_sc_hd__nor2_2 _34904_ (.A(_13257_),
    .B(_13258_),
    .Y(_13259_));
 sky130_fd_sc_hd__and2_2 _34905_ (.A(_09319_),
    .B(_08186_),
    .X(_13260_));
 sky130_vsdinv _34906_ (.A(_13260_),
    .Y(_13261_));
 sky130_fd_sc_hd__nand2_2 _34907_ (.A(_13257_),
    .B(_13258_),
    .Y(_13262_));
 sky130_fd_sc_hd__nor3b_2 _34908_ (.A(_13259_),
    .B(_13261_),
    .C_N(_13262_),
    .Y(_13263_));
 sky130_fd_sc_hd__xnor2_2 _34909_ (.A(_13257_),
    .B(_13258_),
    .Y(_13264_));
 sky130_fd_sc_hd__nand2_2 _34910_ (.A(_13264_),
    .B(_13261_),
    .Y(_13265_));
 sky130_fd_sc_hd__and2b_2 _34911_ (.A_N(_13263_),
    .B(_13265_),
    .X(_13266_));
 sky130_fd_sc_hd__a21oi_2 _34912_ (.A1(_13255_),
    .A2(_13256_),
    .B1(_13266_),
    .Y(_13267_));
 sky130_fd_sc_hd__nand3_2 _34913_ (.A(_13255_),
    .B(_13266_),
    .C(_13256_),
    .Y(_13268_));
 sky130_vsdinv _34914_ (.A(_13268_),
    .Y(_13269_));
 sky130_fd_sc_hd__a21oi_2 _34915_ (.A1(_13005_),
    .A2(_13006_),
    .B1(_13007_),
    .Y(_13270_));
 sky130_fd_sc_hd__xnor2_2 _34916_ (.A(_13010_),
    .B(_13013_),
    .Y(_13271_));
 sky130_fd_sc_hd__o21ai_2 _34917_ (.A1(_13270_),
    .A2(_13271_),
    .B1(_13009_),
    .Y(_13272_));
 sky130_fd_sc_hd__o21bai_2 _34918_ (.A1(_13267_),
    .A2(_13269_),
    .B1_N(_13272_),
    .Y(_13273_));
 sky130_fd_sc_hd__a21o_2 _34919_ (.A1(_13255_),
    .A2(_13256_),
    .B1(_13266_),
    .X(_13274_));
 sky130_fd_sc_hd__nand3_2 _34920_ (.A(_13274_),
    .B(_13268_),
    .C(_13272_),
    .Y(_13275_));
 sky130_fd_sc_hd__nand2_2 _34921_ (.A(_18727_),
    .B(_08261_),
    .Y(_13276_));
 sky130_fd_sc_hd__nand2_2 _34922_ (.A(_08754_),
    .B(_08254_),
    .Y(_13277_));
 sky130_fd_sc_hd__xor2_2 _34923_ (.A(_13276_),
    .B(_13277_),
    .X(_13278_));
 sky130_fd_sc_hd__nand3_2 _34924_ (.A(_13278_),
    .B(_08458_),
    .C(_07948_),
    .Y(_13279_));
 sky130_fd_sc_hd__xnor2_2 _34925_ (.A(_13276_),
    .B(_13277_),
    .Y(_13280_));
 sky130_fd_sc_hd__o21ai_2 _34926_ (.A1(_10245_),
    .A2(_08524_),
    .B1(_13280_),
    .Y(_13281_));
 sky130_vsdinv _34927_ (.A(_13011_),
    .Y(_13282_));
 sky130_fd_sc_hd__a21o_2 _34928_ (.A1(_13282_),
    .A2(_13010_),
    .B1(_13012_),
    .X(_13283_));
 sky130_fd_sc_hd__a21o_2 _34929_ (.A1(_13279_),
    .A2(_13281_),
    .B1(_13283_),
    .X(_13284_));
 sky130_fd_sc_hd__nand3_2 _34930_ (.A(_13279_),
    .B(_13283_),
    .C(_13281_),
    .Y(_13285_));
 sky130_fd_sc_hd__buf_1 _34931_ (.A(_13285_),
    .X(_13286_));
 sky130_fd_sc_hd__o21ai_2 _34932_ (.A1(_13023_),
    .A2(_13024_),
    .B1(_13027_),
    .Y(_13287_));
 sky130_fd_sc_hd__a21o_2 _34933_ (.A1(_13284_),
    .A2(_13286_),
    .B1(_13287_),
    .X(_13288_));
 sky130_fd_sc_hd__nand3_2 _34934_ (.A(_13284_),
    .B(_13287_),
    .C(_13285_),
    .Y(_13289_));
 sky130_fd_sc_hd__nand2_2 _34935_ (.A(_13288_),
    .B(_13289_),
    .Y(_13290_));
 sky130_fd_sc_hd__buf_1 _34936_ (.A(_13290_),
    .X(_13291_));
 sky130_fd_sc_hd__a21boi_2 _34937_ (.A1(_13273_),
    .A2(_13275_),
    .B1_N(_13291_),
    .Y(_13292_));
 sky130_fd_sc_hd__nand2_2 _34938_ (.A(_13273_),
    .B(_13275_),
    .Y(_13293_));
 sky130_fd_sc_hd__nor2_2 _34939_ (.A(_13291_),
    .B(_13293_),
    .Y(_13294_));
 sky130_fd_sc_hd__a21oi_2 _34940_ (.A1(_13020_),
    .A2(_13016_),
    .B1(_13018_),
    .Y(_13295_));
 sky130_fd_sc_hd__o21ai_2 _34941_ (.A1(_13037_),
    .A2(_13295_),
    .B1(_13021_),
    .Y(_13296_));
 sky130_fd_sc_hd__o21bai_2 _34942_ (.A1(_13292_),
    .A2(_13294_),
    .B1_N(_13296_),
    .Y(_13297_));
 sky130_fd_sc_hd__nand2_2 _34943_ (.A(_13293_),
    .B(_13291_),
    .Y(_13298_));
 sky130_fd_sc_hd__nand3b_2 _34944_ (.A_N(_13290_),
    .B(_13275_),
    .C(_13273_),
    .Y(_13299_));
 sky130_fd_sc_hd__nand3_2 _34945_ (.A(_13298_),
    .B(_13296_),
    .C(_13299_),
    .Y(_13300_));
 sky130_fd_sc_hd__buf_1 _34946_ (.A(_13300_),
    .X(_13301_));
 sky130_fd_sc_hd__nand2_2 _34947_ (.A(_10186_),
    .B(_07748_),
    .Y(_13302_));
 sky130_fd_sc_hd__nand2_2 _34948_ (.A(_18753_),
    .B(_08551_),
    .Y(_13303_));
 sky130_fd_sc_hd__nand2_2 _34949_ (.A(_13302_),
    .B(_13303_),
    .Y(_13304_));
 sky130_fd_sc_hd__buf_1 _34950_ (.A(_09548_),
    .X(_13305_));
 sky130_fd_sc_hd__nand3b_2 _34951_ (.A_N(_13302_),
    .B(_13305_),
    .C(_08303_),
    .Y(_13306_));
 sky130_fd_sc_hd__o2bb2ai_2 _34952_ (.A1_N(_13304_),
    .A2_N(_13306_),
    .B1(_08231_),
    .B2(_12845_),
    .Y(_13307_));
 sky130_fd_sc_hd__and2_2 _34953_ (.A(_11080_),
    .B(_10159_),
    .X(_13308_));
 sky130_fd_sc_hd__nand3_2 _34954_ (.A(_13306_),
    .B(_13304_),
    .C(_13308_),
    .Y(_13309_));
 sky130_fd_sc_hd__nor2_2 _34955_ (.A(_13046_),
    .B(_13047_),
    .Y(_13310_));
 sky130_fd_sc_hd__a21oi_2 _34956_ (.A1(_13048_),
    .A2(_13052_),
    .B1(_13310_),
    .Y(_13311_));
 sky130_vsdinv _34957_ (.A(_13311_),
    .Y(_13312_));
 sky130_fd_sc_hd__a21oi_2 _34958_ (.A1(_13307_),
    .A2(_13309_),
    .B1(_13312_),
    .Y(_13313_));
 sky130_fd_sc_hd__nand3_2 _34959_ (.A(_13307_),
    .B(_13312_),
    .C(_13309_),
    .Y(_13314_));
 sky130_vsdinv _34960_ (.A(_13314_),
    .Y(_13315_));
 sky130_fd_sc_hd__and2_2 _34961_ (.A(_11064_),
    .B(_11434_),
    .X(_13316_));
 sky130_fd_sc_hd__nand2_2 _34962_ (.A(_07851_),
    .B(_08570_),
    .Y(_13317_));
 sky130_fd_sc_hd__nand2_2 _34963_ (.A(_10207_),
    .B(_09216_),
    .Y(_13318_));
 sky130_fd_sc_hd__xnor2_2 _34964_ (.A(_13317_),
    .B(_13318_),
    .Y(_13319_));
 sky130_fd_sc_hd__xnor2_2 _34965_ (.A(_13316_),
    .B(_13319_),
    .Y(_13320_));
 sky130_fd_sc_hd__o21bai_2 _34966_ (.A1(_13313_),
    .A2(_13315_),
    .B1_N(_13320_),
    .Y(_13321_));
 sky130_fd_sc_hd__nand3b_2 _34967_ (.A_N(_13313_),
    .B(_13320_),
    .C(_13314_),
    .Y(_13322_));
 sky130_fd_sc_hd__a21oi_2 _34968_ (.A1(_13027_),
    .A2(_13029_),
    .B1(_13031_),
    .Y(_13323_));
 sky130_fd_sc_hd__o21ai_2 _34969_ (.A1(_13034_),
    .A2(_13323_),
    .B1(_13033_),
    .Y(_13324_));
 sky130_fd_sc_hd__a21o_2 _34970_ (.A1(_13321_),
    .A2(_13322_),
    .B1(_13324_),
    .X(_13325_));
 sky130_fd_sc_hd__nand3_2 _34971_ (.A(_13321_),
    .B(_13324_),
    .C(_13322_),
    .Y(_13326_));
 sky130_fd_sc_hd__a21boi_2 _34972_ (.A1(_13063_),
    .A2(_13057_),
    .B1_N(_13058_),
    .Y(_13327_));
 sky130_vsdinv _34973_ (.A(_13327_),
    .Y(_13328_));
 sky130_fd_sc_hd__a21o_2 _34974_ (.A1(_13325_),
    .A2(_13326_),
    .B1(_13328_),
    .X(_13329_));
 sky130_fd_sc_hd__nand3_2 _34975_ (.A(_13325_),
    .B(_13328_),
    .C(_13326_),
    .Y(_13330_));
 sky130_fd_sc_hd__nand2_2 _34976_ (.A(_13329_),
    .B(_13330_),
    .Y(_13331_));
 sky130_fd_sc_hd__buf_1 _34977_ (.A(_13331_),
    .X(_13332_));
 sky130_fd_sc_hd__a21boi_2 _34978_ (.A1(_13297_),
    .A2(_13301_),
    .B1_N(_13332_),
    .Y(_13333_));
 sky130_fd_sc_hd__a21oi_2 _34979_ (.A1(_13298_),
    .A2(_13299_),
    .B1(_13296_),
    .Y(_13334_));
 sky130_fd_sc_hd__nor3b_2 _34980_ (.A(_13332_),
    .B(_13334_),
    .C_N(_13301_),
    .Y(_13335_));
 sky130_fd_sc_hd__o21ai_2 _34981_ (.A1(_13076_),
    .A2(_13077_),
    .B1(_13045_),
    .Y(_13336_));
 sky130_fd_sc_hd__o21bai_2 _34982_ (.A1(_13333_),
    .A2(_13335_),
    .B1_N(_13336_),
    .Y(_13337_));
 sky130_fd_sc_hd__nand2_2 _34983_ (.A(_13297_),
    .B(_13300_),
    .Y(_13338_));
 sky130_fd_sc_hd__nand2_2 _34984_ (.A(_13338_),
    .B(_13332_),
    .Y(_13339_));
 sky130_fd_sc_hd__nand3b_2 _34985_ (.A_N(_13331_),
    .B(_13297_),
    .C(_13301_),
    .Y(_13340_));
 sky130_fd_sc_hd__nand3_2 _34986_ (.A(_13339_),
    .B(_13340_),
    .C(_13336_),
    .Y(_13341_));
 sky130_fd_sc_hd__buf_1 _34987_ (.A(_13341_),
    .X(_13342_));
 sky130_fd_sc_hd__a22o_2 _34988_ (.A1(_08011_),
    .A2(_09497_),
    .B1(_08013_),
    .B2(_11736_),
    .X(_13343_));
 sky130_fd_sc_hd__nand2_2 _34989_ (.A(_10356_),
    .B(_09493_),
    .Y(_13344_));
 sky130_fd_sc_hd__nand3b_2 _34990_ (.A_N(_13344_),
    .B(_12289_),
    .C(_12325_),
    .Y(_13345_));
 sky130_fd_sc_hd__o2bb2ai_2 _34991_ (.A1_N(_13343_),
    .A2_N(_13345_),
    .B1(_08918_),
    .B2(_19163_),
    .Y(_13346_));
 sky130_fd_sc_hd__and2_2 _34992_ (.A(_07402_),
    .B(_10042_),
    .X(_13347_));
 sky130_fd_sc_hd__nand3_2 _34993_ (.A(_13345_),
    .B(_13343_),
    .C(_13347_),
    .Y(_13348_));
 sky130_fd_sc_hd__nand2_2 _34994_ (.A(_13060_),
    .B(_13061_),
    .Y(_13349_));
 sky130_fd_sc_hd__nor2_2 _34995_ (.A(_13060_),
    .B(_13061_),
    .Y(_13350_));
 sky130_fd_sc_hd__a21oi_2 _34996_ (.A1(_13349_),
    .A2(_13059_),
    .B1(_13350_),
    .Y(_13351_));
 sky130_fd_sc_hd__a21boi_2 _34997_ (.A1(_13346_),
    .A2(_13348_),
    .B1_N(_13351_),
    .Y(_13352_));
 sky130_fd_sc_hd__nand3b_2 _34998_ (.A_N(_13351_),
    .B(_13346_),
    .C(_13348_),
    .Y(_13353_));
 sky130_vsdinv _34999_ (.A(_13353_),
    .Y(_13354_));
 sky130_fd_sc_hd__o21ai_2 _35000_ (.A1(_13086_),
    .A2(_13087_),
    .B1(_13090_),
    .Y(_13355_));
 sky130_fd_sc_hd__o21bai_2 _35001_ (.A1(_13352_),
    .A2(_13354_),
    .B1_N(_13355_),
    .Y(_13356_));
 sky130_fd_sc_hd__a21bo_2 _35002_ (.A1(_13346_),
    .A2(_13348_),
    .B1_N(_13351_),
    .X(_13357_));
 sky130_fd_sc_hd__nand3_2 _35003_ (.A(_13357_),
    .B(_13355_),
    .C(_13353_),
    .Y(_13358_));
 sky130_fd_sc_hd__a21boi_2 _35004_ (.A1(_13090_),
    .A2(_13092_),
    .B1_N(_13093_),
    .Y(_13359_));
 sky130_fd_sc_hd__o21ai_2 _35005_ (.A1(_13096_),
    .A2(_13359_),
    .B1(_13095_),
    .Y(_13360_));
 sky130_fd_sc_hd__a21o_2 _35006_ (.A1(_13356_),
    .A2(_13358_),
    .B1(_13360_),
    .X(_13361_));
 sky130_fd_sc_hd__nand3_2 _35007_ (.A(_13360_),
    .B(_13356_),
    .C(_13358_),
    .Y(_13362_));
 sky130_fd_sc_hd__and2_2 _35008_ (.A(_16960_),
    .B(_06136_),
    .X(_13363_));
 sky130_fd_sc_hd__inv_2 _35009_ (.A(_13363_),
    .Y(_13364_));
 sky130_fd_sc_hd__nand2_2 _35010_ (.A(_18815_),
    .B(_10913_),
    .Y(_13365_));
 sky130_fd_sc_hd__nand2_2 _35011_ (.A(_06268_),
    .B(_19133_),
    .Y(_13366_));
 sky130_fd_sc_hd__xnor2_2 _35012_ (.A(_13365_),
    .B(_13366_),
    .Y(_13367_));
 sky130_fd_sc_hd__xor2_2 _35013_ (.A(_13364_),
    .B(_13367_),
    .X(_13368_));
 sky130_fd_sc_hd__buf_1 _35014_ (.A(_11788_),
    .X(_13369_));
 sky130_fd_sc_hd__nand3b_2 _35015_ (.A_N(_13110_),
    .B(_18804_),
    .C(_13369_),
    .Y(_13370_));
 sky130_fd_sc_hd__nand2_2 _35016_ (.A(_13115_),
    .B(_13370_),
    .Y(_13371_));
 sky130_fd_sc_hd__a22o_2 _35017_ (.A1(_07199_),
    .A2(_10535_),
    .B1(_08034_),
    .B2(_09500_),
    .X(_13372_));
 sky130_fd_sc_hd__nand2_2 _35018_ (.A(_06544_),
    .B(_10532_),
    .Y(_13373_));
 sky130_fd_sc_hd__nand3b_2 _35019_ (.A_N(_13373_),
    .B(_07201_),
    .C(_11515_),
    .Y(_13374_));
 sky130_fd_sc_hd__o2bb2ai_2 _35020_ (.A1_N(_13372_),
    .A2_N(_13374_),
    .B1(_06692_),
    .B2(_19146_),
    .Y(_13375_));
 sky130_fd_sc_hd__and2_2 _35021_ (.A(_08039_),
    .B(_10555_),
    .X(_13376_));
 sky130_fd_sc_hd__nand3_2 _35022_ (.A(_13374_),
    .B(_13372_),
    .C(_13376_),
    .Y(_13377_));
 sky130_fd_sc_hd__nand3_2 _35023_ (.A(_13371_),
    .B(_13375_),
    .C(_13377_),
    .Y(_13378_));
 sky130_fd_sc_hd__nand2_2 _35024_ (.A(_13375_),
    .B(_13377_),
    .Y(_13379_));
 sky130_fd_sc_hd__nand3_2 _35025_ (.A(_13379_),
    .B(_13370_),
    .C(_13115_),
    .Y(_13380_));
 sky130_fd_sc_hd__nand2_2 _35026_ (.A(_13378_),
    .B(_13380_),
    .Y(_13381_));
 sky130_fd_sc_hd__xnor2_2 _35027_ (.A(_13368_),
    .B(_13381_),
    .Y(_13382_));
 sky130_fd_sc_hd__a21oi_2 _35028_ (.A1(_13361_),
    .A2(_13362_),
    .B1(_13382_),
    .Y(_13383_));
 sky130_fd_sc_hd__nand3_2 _35029_ (.A(_13382_),
    .B(_13362_),
    .C(_13361_),
    .Y(_13384_));
 sky130_vsdinv _35030_ (.A(_13384_),
    .Y(_13385_));
 sky130_fd_sc_hd__a21boi_2 _35031_ (.A1(_13068_),
    .A2(_13071_),
    .B1_N(_13069_),
    .Y(_13386_));
 sky130_fd_sc_hd__o21ai_2 _35032_ (.A1(_13383_),
    .A2(_13385_),
    .B1(_13386_),
    .Y(_13387_));
 sky130_fd_sc_hd__nand2_2 _35033_ (.A(_13073_),
    .B(_13069_),
    .Y(_13388_));
 sky130_fd_sc_hd__nand3b_2 _35034_ (.A_N(_13383_),
    .B(_13388_),
    .C(_13384_),
    .Y(_13389_));
 sky130_vsdinv _35035_ (.A(_13103_),
    .Y(_13390_));
 sky130_fd_sc_hd__a21oi_2 _35036_ (.A1(_13125_),
    .A2(_13102_),
    .B1(_13390_),
    .Y(_13391_));
 sky130_vsdinv _35037_ (.A(_13391_),
    .Y(_13392_));
 sky130_fd_sc_hd__a21oi_2 _35038_ (.A1(_13387_),
    .A2(_13389_),
    .B1(_13392_),
    .Y(_13393_));
 sky130_fd_sc_hd__nand3_2 _35039_ (.A(_13387_),
    .B(_13389_),
    .C(_13392_),
    .Y(_13394_));
 sky130_fd_sc_hd__and2b_2 _35040_ (.A_N(_13393_),
    .B(_13394_),
    .X(_13395_));
 sky130_fd_sc_hd__a21oi_2 _35041_ (.A1(_13337_),
    .A2(_13342_),
    .B1(_13395_),
    .Y(_13396_));
 sky130_fd_sc_hd__a21o_2 _35042_ (.A1(_13387_),
    .A2(_13389_),
    .B1(_13392_),
    .X(_13397_));
 sky130_fd_sc_hd__nand2_2 _35043_ (.A(_13397_),
    .B(_13394_),
    .Y(_13398_));
 sky130_fd_sc_hd__a21oi_2 _35044_ (.A1(_13339_),
    .A2(_13340_),
    .B1(_13336_),
    .Y(_13399_));
 sky130_vsdinv _35045_ (.A(_13342_),
    .Y(_13400_));
 sky130_fd_sc_hd__nor3_2 _35046_ (.A(_13398_),
    .B(_13399_),
    .C(_13400_),
    .Y(_13401_));
 sky130_fd_sc_hd__o21ai_2 _35047_ (.A1(_13136_),
    .A2(_13138_),
    .B1(_13085_),
    .Y(_13402_));
 sky130_fd_sc_hd__o21bai_2 _35048_ (.A1(_13396_),
    .A2(_13401_),
    .B1_N(_13402_),
    .Y(_13403_));
 sky130_fd_sc_hd__nand2_2 _35049_ (.A(_13337_),
    .B(_13341_),
    .Y(_13404_));
 sky130_fd_sc_hd__nand2_2 _35050_ (.A(_13404_),
    .B(_13398_),
    .Y(_13405_));
 sky130_fd_sc_hd__nand3_2 _35051_ (.A(_13395_),
    .B(_13342_),
    .C(_13337_),
    .Y(_13406_));
 sky130_fd_sc_hd__nand3_2 _35052_ (.A(_13405_),
    .B(_13402_),
    .C(_13406_),
    .Y(_13407_));
 sky130_vsdinv _35053_ (.A(_13154_),
    .Y(_13408_));
 sky130_fd_sc_hd__a21oi_2 _35054_ (.A1(_13153_),
    .A2(_12636_),
    .B1(_13408_),
    .Y(_13409_));
 sky130_fd_sc_hd__nand2_2 _35055_ (.A(_13106_),
    .B(_13107_),
    .Y(_13410_));
 sky130_fd_sc_hd__nor2_2 _35056_ (.A(_13106_),
    .B(_13107_),
    .Y(_13411_));
 sky130_fd_sc_hd__a21oi_2 _35057_ (.A1(_13410_),
    .A2(_13105_),
    .B1(_13411_),
    .Y(_13412_));
 sky130_fd_sc_hd__buf_1 _35058_ (.A(_13156_),
    .X(_13413_));
 sky130_fd_sc_hd__nor3_2 _35059_ (.A(_13161_),
    .B(_13412_),
    .C(_13413_),
    .Y(_13414_));
 sky130_fd_sc_hd__o21ai_2 _35060_ (.A1(_13161_),
    .A2(_13163_),
    .B1(_13412_),
    .Y(_13415_));
 sky130_fd_sc_hd__nor3b_2 _35061_ (.A(_13409_),
    .B(_13414_),
    .C_N(_13415_),
    .Y(_13416_));
 sky130_vsdinv _35062_ (.A(_13414_),
    .Y(_13417_));
 sky130_vsdinv _35063_ (.A(_13409_),
    .Y(_13418_));
 sky130_fd_sc_hd__buf_1 _35064_ (.A(_13418_),
    .X(_13419_));
 sky130_fd_sc_hd__a21oi_2 _35065_ (.A1(_13417_),
    .A2(_13415_),
    .B1(_13419_),
    .Y(_13420_));
 sky130_fd_sc_hd__o21ai_2 _35066_ (.A1(_13109_),
    .A2(_13119_),
    .B1(_13120_),
    .Y(_13421_));
 sky130_fd_sc_hd__o21bai_2 _35067_ (.A1(_13416_),
    .A2(_13420_),
    .B1_N(_13421_),
    .Y(_13422_));
 sky130_vsdinv _35068_ (.A(_13416_),
    .Y(_13423_));
 sky130_fd_sc_hd__nand3b_2 _35069_ (.A_N(_13420_),
    .B(_13421_),
    .C(_13423_),
    .Y(_13424_));
 sky130_fd_sc_hd__a21boi_2 _35070_ (.A1(_13166_),
    .A2(_13164_),
    .B1_N(_13160_),
    .Y(_13425_));
 sky130_vsdinv _35071_ (.A(_13425_),
    .Y(_13426_));
 sky130_fd_sc_hd__a21o_2 _35072_ (.A1(_13422_),
    .A2(_13424_),
    .B1(_13426_),
    .X(_13427_));
 sky130_fd_sc_hd__nand3_2 _35073_ (.A(_13422_),
    .B(_13426_),
    .C(_13424_),
    .Y(_13428_));
 sky130_fd_sc_hd__nand2_2 _35074_ (.A(_13177_),
    .B(_13171_),
    .Y(_13429_));
 sky130_fd_sc_hd__a21o_2 _35075_ (.A1(_13427_),
    .A2(_13428_),
    .B1(_13429_),
    .X(_13430_));
 sky130_fd_sc_hd__nand3_2 _35076_ (.A(_13429_),
    .B(_13427_),
    .C(_13428_),
    .Y(_13431_));
 sky130_fd_sc_hd__buf_1 _35077_ (.A(_12946_),
    .X(_13432_));
 sky130_fd_sc_hd__a21oi_2 _35078_ (.A1(_13430_),
    .A2(_13431_),
    .B1(_13432_),
    .Y(_13433_));
 sky130_fd_sc_hd__nand3_2 _35079_ (.A(_13430_),
    .B(_13432_),
    .C(_13431_),
    .Y(_13434_));
 sky130_vsdinv _35080_ (.A(_13434_),
    .Y(_13435_));
 sky130_fd_sc_hd__o21ai_2 _35081_ (.A1(_13131_),
    .A2(_13128_),
    .B1(_13129_),
    .Y(_13436_));
 sky130_fd_sc_hd__o21bai_2 _35082_ (.A1(_13433_),
    .A2(_13435_),
    .B1_N(_13436_),
    .Y(_13437_));
 sky130_fd_sc_hd__nand3b_2 _35083_ (.A_N(_13433_),
    .B(_13436_),
    .C(_13434_),
    .Y(_13438_));
 sky130_fd_sc_hd__nand2_2 _35084_ (.A(_13437_),
    .B(_13438_),
    .Y(_13439_));
 sky130_fd_sc_hd__buf_1 _35085_ (.A(_12944_),
    .X(_13440_));
 sky130_fd_sc_hd__a21boi_2 _35086_ (.A1(_13180_),
    .A2(_13440_),
    .B1_N(_13182_),
    .Y(_13441_));
 sky130_fd_sc_hd__nand2_2 _35087_ (.A(_13439_),
    .B(_13441_),
    .Y(_13442_));
 sky130_fd_sc_hd__nand3b_2 _35088_ (.A_N(_13441_),
    .B(_13437_),
    .C(_13438_),
    .Y(_13443_));
 sky130_fd_sc_hd__nand2_2 _35089_ (.A(_13442_),
    .B(_13443_),
    .Y(_13444_));
 sky130_fd_sc_hd__buf_1 _35090_ (.A(_13444_),
    .X(_13445_));
 sky130_fd_sc_hd__a21boi_2 _35091_ (.A1(_13403_),
    .A2(_13407_),
    .B1_N(_13445_),
    .Y(_13446_));
 sky130_fd_sc_hd__a21oi_2 _35092_ (.A1(_13405_),
    .A2(_13406_),
    .B1(_13402_),
    .Y(_13447_));
 sky130_vsdinv _35093_ (.A(_13407_),
    .Y(_13448_));
 sky130_fd_sc_hd__nor3_2 _35094_ (.A(_13445_),
    .B(_13447_),
    .C(_13448_),
    .Y(_13449_));
 sky130_fd_sc_hd__o21ai_2 _35095_ (.A1(_13200_),
    .A2(_13201_),
    .B1(_13148_),
    .Y(_13450_));
 sky130_fd_sc_hd__o21bai_2 _35096_ (.A1(_13446_),
    .A2(_13449_),
    .B1_N(_13450_),
    .Y(_13451_));
 sky130_fd_sc_hd__o21ai_2 _35097_ (.A1(_13447_),
    .A2(_13448_),
    .B1(_13445_),
    .Y(_13452_));
 sky130_fd_sc_hd__nand3b_2 _35098_ (.A_N(_13444_),
    .B(_13403_),
    .C(_13407_),
    .Y(_13453_));
 sky130_fd_sc_hd__nand3_2 _35099_ (.A(_13452_),
    .B(_13453_),
    .C(_13450_),
    .Y(_13454_));
 sky130_fd_sc_hd__buf_1 _35100_ (.A(_13454_),
    .X(_13455_));
 sky130_fd_sc_hd__buf_1 _35101_ (.A(_13211_),
    .X(_13456_));
 sky130_fd_sc_hd__a21oi_2 _35102_ (.A1(_13197_),
    .A2(_13192_),
    .B1(_13456_),
    .Y(_13457_));
 sky130_fd_sc_hd__and3_2 _35103_ (.A(_13197_),
    .B(_13456_),
    .C(_13192_),
    .X(_13458_));
 sky130_fd_sc_hd__nor2_2 _35104_ (.A(_13457_),
    .B(_13458_),
    .Y(_13459_));
 sky130_fd_sc_hd__a21oi_2 _35105_ (.A1(_13451_),
    .A2(_13455_),
    .B1(_13459_),
    .Y(_13460_));
 sky130_fd_sc_hd__nand3_2 _35106_ (.A(_13451_),
    .B(_13459_),
    .C(_13454_),
    .Y(_13461_));
 sky130_vsdinv _35107_ (.A(_13461_),
    .Y(_13462_));
 sky130_fd_sc_hd__o21ai_2 _35108_ (.A1(_13217_),
    .A2(_13218_),
    .B1(_13210_),
    .Y(_13463_));
 sky130_fd_sc_hd__o21bai_2 _35109_ (.A1(_13460_),
    .A2(_13462_),
    .B1_N(_13463_),
    .Y(_13464_));
 sky130_fd_sc_hd__o2bb2ai_2 _35110_ (.A1_N(_13455_),
    .A2_N(_13451_),
    .B1(_13457_),
    .B2(_13458_),
    .Y(_13465_));
 sky130_fd_sc_hd__nand3_2 _35111_ (.A(_13465_),
    .B(_13461_),
    .C(_13463_),
    .Y(_13466_));
 sky130_fd_sc_hd__buf_1 _35112_ (.A(_13456_),
    .X(_13467_));
 sky130_fd_sc_hd__buf_1 _35113_ (.A(_13467_),
    .X(_13468_));
 sky130_fd_sc_hd__a21oi_2 _35114_ (.A1(_12961_),
    .A2(_12953_),
    .B1(_13468_),
    .Y(_13469_));
 sky130_fd_sc_hd__a21oi_2 _35115_ (.A1(_13464_),
    .A2(_13466_),
    .B1(_13469_),
    .Y(_13470_));
 sky130_fd_sc_hd__nand3_2 _35116_ (.A(_13464_),
    .B(_13469_),
    .C(_13466_),
    .Y(_13471_));
 sky130_vsdinv _35117_ (.A(_13471_),
    .Y(_13472_));
 sky130_fd_sc_hd__o21ai_2 _35118_ (.A1(_13229_),
    .A2(_13230_),
    .B1(_13226_),
    .Y(_13473_));
 sky130_fd_sc_hd__o21bai_2 _35119_ (.A1(_13470_),
    .A2(_13472_),
    .B1_N(_13473_),
    .Y(_13474_));
 sky130_fd_sc_hd__a21o_2 _35120_ (.A1(_13464_),
    .A2(_13466_),
    .B1(_13469_),
    .X(_13475_));
 sky130_fd_sc_hd__nand3_2 _35121_ (.A(_13475_),
    .B(_13473_),
    .C(_13471_),
    .Y(_13476_));
 sky130_fd_sc_hd__nand2_2 _35122_ (.A(_13474_),
    .B(_13476_),
    .Y(_13477_));
 sky130_fd_sc_hd__o21ai_2 _35123_ (.A1(_13238_),
    .A2(_13247_),
    .B1(_13237_),
    .Y(_13478_));
 sky130_fd_sc_hd__xnor2_2 _35124_ (.A(_13477_),
    .B(_13478_),
    .Y(_02660_));
 sky130_fd_sc_hd__nand2_2 _35125_ (.A(_10486_),
    .B(_19248_),
    .Y(_13479_));
 sky130_fd_sc_hd__nand3b_2 _35126_ (.A_N(_13479_),
    .B(_12183_),
    .C(_19253_),
    .Y(_13480_));
 sky130_fd_sc_hd__o21ai_2 _35127_ (.A1(_06883_),
    .A2(_11331_),
    .B1(_13479_),
    .Y(_13481_));
 sky130_fd_sc_hd__and2_2 _35128_ (.A(_10483_),
    .B(_07264_),
    .X(_13482_));
 sky130_fd_sc_hd__a21o_2 _35129_ (.A1(_13480_),
    .A2(_13481_),
    .B1(_13482_),
    .X(_13483_));
 sky130_fd_sc_hd__nand3_2 _35130_ (.A(_13480_),
    .B(_13482_),
    .C(_13481_),
    .Y(_13484_));
 sky130_fd_sc_hd__nand2_2 _35131_ (.A(_13253_),
    .B(_13249_),
    .Y(_13485_));
 sky130_fd_sc_hd__a21o_2 _35132_ (.A1(_13483_),
    .A2(_13484_),
    .B1(_13485_),
    .X(_13486_));
 sky130_fd_sc_hd__nand3_2 _35133_ (.A(_13485_),
    .B(_13483_),
    .C(_13484_),
    .Y(_13487_));
 sky130_fd_sc_hd__and2_2 _35134_ (.A(_09320_),
    .B(_06596_),
    .X(_13488_));
 sky130_fd_sc_hd__nand2_2 _35135_ (.A(_11014_),
    .B(_08181_),
    .Y(_13489_));
 sky130_fd_sc_hd__nand2_2 _35136_ (.A(_10686_),
    .B(_07698_),
    .Y(_13490_));
 sky130_fd_sc_hd__xnor2_2 _35137_ (.A(_13489_),
    .B(_13490_),
    .Y(_13491_));
 sky130_fd_sc_hd__xnor2_2 _35138_ (.A(_13488_),
    .B(_13491_),
    .Y(_13492_));
 sky130_fd_sc_hd__a21oi_2 _35139_ (.A1(_13486_),
    .A2(_13487_),
    .B1(_13492_),
    .Y(_13493_));
 sky130_fd_sc_hd__a21oi_2 _35140_ (.A1(_13483_),
    .A2(_13484_),
    .B1(_13485_),
    .Y(_13494_));
 sky130_fd_sc_hd__xor2_2 _35141_ (.A(_13488_),
    .B(_13491_),
    .X(_13495_));
 sky130_vsdinv _35142_ (.A(_13487_),
    .Y(_13496_));
 sky130_fd_sc_hd__nor3_2 _35143_ (.A(_13494_),
    .B(_13495_),
    .C(_13496_),
    .Y(_13497_));
 sky130_fd_sc_hd__a21oi_2 _35144_ (.A1(_13252_),
    .A2(_13253_),
    .B1(_13254_),
    .Y(_13498_));
 sky130_fd_sc_hd__or2b_2 _35145_ (.A(_13263_),
    .B_N(_13265_),
    .X(_13499_));
 sky130_fd_sc_hd__o21ai_2 _35146_ (.A1(_13498_),
    .A2(_13499_),
    .B1(_13256_),
    .Y(_13500_));
 sky130_fd_sc_hd__o21bai_2 _35147_ (.A1(_13493_),
    .A2(_13497_),
    .B1_N(_13500_),
    .Y(_13501_));
 sky130_fd_sc_hd__o21bai_2 _35148_ (.A1(_13494_),
    .A2(_13496_),
    .B1_N(_13492_),
    .Y(_13502_));
 sky130_fd_sc_hd__nand3_2 _35149_ (.A(_13486_),
    .B(_13492_),
    .C(_13487_),
    .Y(_13503_));
 sky130_fd_sc_hd__nand3_2 _35150_ (.A(_13502_),
    .B(_13503_),
    .C(_13500_),
    .Y(_13504_));
 sky130_fd_sc_hd__nand2_2 _35151_ (.A(_11634_),
    .B(_07328_),
    .Y(_13505_));
 sky130_fd_sc_hd__nand2_2 _35152_ (.A(_10231_),
    .B(_07321_),
    .Y(_13506_));
 sky130_fd_sc_hd__xor2_2 _35153_ (.A(_13505_),
    .B(_13506_),
    .X(_13507_));
 sky130_fd_sc_hd__buf_1 _35154_ (.A(_08759_),
    .X(_13508_));
 sky130_fd_sc_hd__nand3_2 _35155_ (.A(_13507_),
    .B(_13508_),
    .C(_08301_),
    .Y(_13509_));
 sky130_fd_sc_hd__xnor2_2 _35156_ (.A(_13505_),
    .B(_13506_),
    .Y(_13510_));
 sky130_fd_sc_hd__o21ai_2 _35157_ (.A1(_12219_),
    .A2(_19208_),
    .B1(_13510_),
    .Y(_13511_));
 sky130_fd_sc_hd__a21oi_2 _35158_ (.A1(_13262_),
    .A2(_13260_),
    .B1(_13259_),
    .Y(_13512_));
 sky130_fd_sc_hd__a21bo_2 _35159_ (.A1(_13509_),
    .A2(_13511_),
    .B1_N(_13512_),
    .X(_13513_));
 sky130_fd_sc_hd__nand3b_2 _35160_ (.A_N(_13512_),
    .B(_13509_),
    .C(_13511_),
    .Y(_13514_));
 sky130_fd_sc_hd__o21ai_2 _35161_ (.A1(_13276_),
    .A2(_13277_),
    .B1(_13279_),
    .Y(_13515_));
 sky130_fd_sc_hd__a21oi_2 _35162_ (.A1(_13513_),
    .A2(_13514_),
    .B1(_13515_),
    .Y(_13516_));
 sky130_fd_sc_hd__nand3_2 _35163_ (.A(_13513_),
    .B(_13515_),
    .C(_13514_),
    .Y(_13517_));
 sky130_vsdinv _35164_ (.A(_13517_),
    .Y(_13518_));
 sky130_fd_sc_hd__nor2_2 _35165_ (.A(_13516_),
    .B(_13518_),
    .Y(_13519_));
 sky130_fd_sc_hd__a21oi_2 _35166_ (.A1(_13501_),
    .A2(_13504_),
    .B1(_13519_),
    .Y(_13520_));
 sky130_fd_sc_hd__a21boi_2 _35167_ (.A1(_13509_),
    .A2(_13511_),
    .B1_N(_13512_),
    .Y(_13521_));
 sky130_vsdinv _35168_ (.A(_13514_),
    .Y(_13522_));
 sky130_fd_sc_hd__o21bai_2 _35169_ (.A1(_13521_),
    .A2(_13522_),
    .B1_N(_13515_),
    .Y(_13523_));
 sky130_fd_sc_hd__nand2_2 _35170_ (.A(_13523_),
    .B(_13517_),
    .Y(_13524_));
 sky130_fd_sc_hd__a21oi_2 _35171_ (.A1(_13502_),
    .A2(_13503_),
    .B1(_13500_),
    .Y(_13525_));
 sky130_vsdinv _35172_ (.A(_13504_),
    .Y(_13526_));
 sky130_fd_sc_hd__nor3_2 _35173_ (.A(_13524_),
    .B(_13525_),
    .C(_13526_),
    .Y(_13527_));
 sky130_fd_sc_hd__a21oi_2 _35174_ (.A1(_13274_),
    .A2(_13268_),
    .B1(_13272_),
    .Y(_13528_));
 sky130_fd_sc_hd__o21ai_2 _35175_ (.A1(_13291_),
    .A2(_13528_),
    .B1(_13275_),
    .Y(_13529_));
 sky130_fd_sc_hd__o21bai_2 _35176_ (.A1(_13520_),
    .A2(_13527_),
    .B1_N(_13529_),
    .Y(_13530_));
 sky130_fd_sc_hd__o22ai_2 _35177_ (.A1(_13518_),
    .A2(_13516_),
    .B1(_13525_),
    .B2(_13526_),
    .Y(_13531_));
 sky130_fd_sc_hd__nand3_2 _35178_ (.A(_13519_),
    .B(_13501_),
    .C(_13504_),
    .Y(_13532_));
 sky130_fd_sc_hd__nand3_2 _35179_ (.A(_13531_),
    .B(_13529_),
    .C(_13532_),
    .Y(_13533_));
 sky130_fd_sc_hd__buf_1 _35180_ (.A(_13533_),
    .X(_13534_));
 sky130_fd_sc_hd__a22o_2 _35181_ (.A1(_12527_),
    .A2(_07751_),
    .B1(_10415_),
    .B2(_08553_),
    .X(_13535_));
 sky130_fd_sc_hd__nand2_2 _35182_ (.A(_08472_),
    .B(_07310_),
    .Y(_13536_));
 sky130_fd_sc_hd__nand3b_2 _35183_ (.A_N(_13536_),
    .B(_13305_),
    .C(_10162_),
    .Y(_13537_));
 sky130_fd_sc_hd__o2bb2ai_2 _35184_ (.A1_N(_13535_),
    .A2_N(_13537_),
    .B1(_08231_),
    .B2(_19192_),
    .Y(_13538_));
 sky130_fd_sc_hd__and2_2 _35185_ (.A(_07845_),
    .B(_09078_),
    .X(_13539_));
 sky130_fd_sc_hd__nand3_2 _35186_ (.A(_13537_),
    .B(_13535_),
    .C(_13539_),
    .Y(_13540_));
 sky130_fd_sc_hd__nor2_2 _35187_ (.A(_13302_),
    .B(_13303_),
    .Y(_13541_));
 sky130_fd_sc_hd__a21oi_2 _35188_ (.A1(_13304_),
    .A2(_13308_),
    .B1(_13541_),
    .Y(_13542_));
 sky130_vsdinv _35189_ (.A(_13542_),
    .Y(_13543_));
 sky130_fd_sc_hd__a21o_2 _35190_ (.A1(_13538_),
    .A2(_13540_),
    .B1(_13543_),
    .X(_13544_));
 sky130_fd_sc_hd__nand3_2 _35191_ (.A(_13538_),
    .B(_13543_),
    .C(_13540_),
    .Y(_13545_));
 sky130_fd_sc_hd__and2_2 _35192_ (.A(_07161_),
    .B(_10843_),
    .X(_13546_));
 sky130_fd_sc_hd__nand2_2 _35193_ (.A(_08215_),
    .B(_10574_),
    .Y(_13547_));
 sky130_fd_sc_hd__nand3b_2 _35194_ (.A_N(_13547_),
    .B(_12805_),
    .C(_12295_),
    .Y(_13548_));
 sky130_fd_sc_hd__a22o_2 _35195_ (.A1(_10745_),
    .A2(_08826_),
    .B1(_12254_),
    .B2(_11434_),
    .X(_13549_));
 sky130_fd_sc_hd__nand2_2 _35196_ (.A(_13548_),
    .B(_13549_),
    .Y(_13550_));
 sky130_fd_sc_hd__xnor2_2 _35197_ (.A(_13546_),
    .B(_13550_),
    .Y(_13551_));
 sky130_fd_sc_hd__a21oi_2 _35198_ (.A1(_13544_),
    .A2(_13545_),
    .B1(_13551_),
    .Y(_13552_));
 sky130_vsdinv _35199_ (.A(_13552_),
    .Y(_13553_));
 sky130_fd_sc_hd__nand3_2 _35200_ (.A(_13544_),
    .B(_13551_),
    .C(_13545_),
    .Y(_13554_));
 sky130_fd_sc_hd__nand2_2 _35201_ (.A(_13289_),
    .B(_13286_),
    .Y(_13555_));
 sky130_fd_sc_hd__a21oi_2 _35202_ (.A1(_13553_),
    .A2(_13554_),
    .B1(_13555_),
    .Y(_13556_));
 sky130_vsdinv _35203_ (.A(_13554_),
    .Y(_13557_));
 sky130_fd_sc_hd__a211oi_2 _35204_ (.A1(_13289_),
    .A2(_13286_),
    .B1(_13552_),
    .C1(_13557_),
    .Y(_13558_));
 sky130_fd_sc_hd__and2_2 _35205_ (.A(_13322_),
    .B(_13314_),
    .X(_13559_));
 sky130_fd_sc_hd__o21ai_2 _35206_ (.A1(_13556_),
    .A2(_13558_),
    .B1(_13559_),
    .Y(_13560_));
 sky130_fd_sc_hd__o211ai_2 _35207_ (.A1(_13552_),
    .A2(_13557_),
    .B1(_13286_),
    .C1(_13289_),
    .Y(_13561_));
 sky130_fd_sc_hd__nand3_2 _35208_ (.A(_13555_),
    .B(_13553_),
    .C(_13554_),
    .Y(_13562_));
 sky130_fd_sc_hd__nand3b_2 _35209_ (.A_N(_13559_),
    .B(_13561_),
    .C(_13562_),
    .Y(_13563_));
 sky130_fd_sc_hd__nand2_2 _35210_ (.A(_13560_),
    .B(_13563_),
    .Y(_13564_));
 sky130_fd_sc_hd__buf_1 _35211_ (.A(_13564_),
    .X(_13565_));
 sky130_fd_sc_hd__a21boi_2 _35212_ (.A1(_13530_),
    .A2(_13534_),
    .B1_N(_13565_),
    .Y(_13566_));
 sky130_fd_sc_hd__a21oi_2 _35213_ (.A1(_13531_),
    .A2(_13532_),
    .B1(_13529_),
    .Y(_13567_));
 sky130_vsdinv _35214_ (.A(_13534_),
    .Y(_13568_));
 sky130_fd_sc_hd__nor3_2 _35215_ (.A(_13565_),
    .B(_13567_),
    .C(_13568_),
    .Y(_13569_));
 sky130_fd_sc_hd__o21ai_2 _35216_ (.A1(_13332_),
    .A2(_13334_),
    .B1(_13301_),
    .Y(_13570_));
 sky130_fd_sc_hd__o21bai_2 _35217_ (.A1(_13566_),
    .A2(_13569_),
    .B1_N(_13570_),
    .Y(_13571_));
 sky130_fd_sc_hd__nand2_2 _35218_ (.A(_13530_),
    .B(_13533_),
    .Y(_13572_));
 sky130_fd_sc_hd__nand2_2 _35219_ (.A(_13572_),
    .B(_13565_),
    .Y(_13573_));
 sky130_fd_sc_hd__nand3b_2 _35220_ (.A_N(_13564_),
    .B(_13534_),
    .C(_13530_),
    .Y(_13574_));
 sky130_fd_sc_hd__nand3_2 _35221_ (.A(_13573_),
    .B(_13574_),
    .C(_13570_),
    .Y(_13575_));
 sky130_fd_sc_hd__buf_1 _35222_ (.A(_13575_),
    .X(_13576_));
 sky130_fd_sc_hd__nand2_2 _35223_ (.A(_18780_),
    .B(_09086_),
    .Y(_13577_));
 sky130_fd_sc_hd__nand2_2 _35224_ (.A(_07470_),
    .B(_10537_),
    .Y(_13578_));
 sky130_fd_sc_hd__xor2_2 _35225_ (.A(_13577_),
    .B(_13578_),
    .X(_13579_));
 sky130_fd_sc_hd__buf_1 _35226_ (.A(_10875_),
    .X(_13580_));
 sky130_fd_sc_hd__nand3_2 _35227_ (.A(_13579_),
    .B(_13089_),
    .C(_13580_),
    .Y(_13581_));
 sky130_fd_sc_hd__xnor2_2 _35228_ (.A(_13577_),
    .B(_13578_),
    .Y(_13582_));
 sky130_fd_sc_hd__o21ai_2 _35229_ (.A1(_11716_),
    .A2(_19158_),
    .B1(_13582_),
    .Y(_13583_));
 sky130_fd_sc_hd__nand2_2 _35230_ (.A(_13317_),
    .B(_13318_),
    .Y(_13584_));
 sky130_fd_sc_hd__nor2_2 _35231_ (.A(_13317_),
    .B(_13318_),
    .Y(_13585_));
 sky130_fd_sc_hd__a21oi_2 _35232_ (.A1(_13584_),
    .A2(_13316_),
    .B1(_13585_),
    .Y(_13586_));
 sky130_vsdinv _35233_ (.A(_13586_),
    .Y(_13587_));
 sky130_fd_sc_hd__a21o_2 _35234_ (.A1(_13581_),
    .A2(_13583_),
    .B1(_13587_),
    .X(_13588_));
 sky130_fd_sc_hd__nand3_2 _35235_ (.A(_13581_),
    .B(_13583_),
    .C(_13587_),
    .Y(_13589_));
 sky130_fd_sc_hd__a21boi_2 _35236_ (.A1(_13343_),
    .A2(_13347_),
    .B1_N(_13345_),
    .Y(_13590_));
 sky130_vsdinv _35237_ (.A(_13590_),
    .Y(_13591_));
 sky130_fd_sc_hd__a21oi_2 _35238_ (.A1(_13588_),
    .A2(_13589_),
    .B1(_13591_),
    .Y(_13592_));
 sky130_fd_sc_hd__nand3_2 _35239_ (.A(_13588_),
    .B(_13591_),
    .C(_13589_),
    .Y(_13593_));
 sky130_vsdinv _35240_ (.A(_13593_),
    .Y(_13594_));
 sky130_fd_sc_hd__a21o_2 _35241_ (.A1(_13357_),
    .A2(_13355_),
    .B1(_13354_),
    .X(_13595_));
 sky130_fd_sc_hd__o21bai_2 _35242_ (.A1(_13592_),
    .A2(_13594_),
    .B1_N(_13595_),
    .Y(_13596_));
 sky130_fd_sc_hd__a21o_2 _35243_ (.A1(_13588_),
    .A2(_13589_),
    .B1(_13591_),
    .X(_13597_));
 sky130_fd_sc_hd__nand3_2 _35244_ (.A(_13597_),
    .B(_13593_),
    .C(_13595_),
    .Y(_13598_));
 sky130_fd_sc_hd__nand2_2 _35245_ (.A(_07190_),
    .B(_09804_),
    .Y(_13599_));
 sky130_fd_sc_hd__nand2_2 _35246_ (.A(_07200_),
    .B(_10554_),
    .Y(_13600_));
 sky130_fd_sc_hd__xor2_2 _35247_ (.A(_13599_),
    .B(_13600_),
    .X(_13601_));
 sky130_fd_sc_hd__and2_2 _35248_ (.A(_06275_),
    .B(_10039_),
    .X(_13602_));
 sky130_fd_sc_hd__nand2_2 _35249_ (.A(_13601_),
    .B(_13602_),
    .Y(_13603_));
 sky130_fd_sc_hd__xnor2_2 _35250_ (.A(_13599_),
    .B(_13600_),
    .Y(_13604_));
 sky130_fd_sc_hd__o21ai_2 _35251_ (.A1(_11745_),
    .A2(_19140_),
    .B1(_13604_),
    .Y(_13605_));
 sky130_fd_sc_hd__nand2_2 _35252_ (.A(_13377_),
    .B(_13374_),
    .Y(_13606_));
 sky130_fd_sc_hd__a21oi_2 _35253_ (.A1(_13603_),
    .A2(_13605_),
    .B1(_13606_),
    .Y(_13607_));
 sky130_fd_sc_hd__nand3_2 _35254_ (.A(_13603_),
    .B(_13605_),
    .C(_13606_),
    .Y(_13608_));
 sky130_vsdinv _35255_ (.A(_13608_),
    .Y(_13609_));
 sky130_fd_sc_hd__nand2_2 _35256_ (.A(_10393_),
    .B(_12097_),
    .Y(_13610_));
 sky130_fd_sc_hd__nand2_2 _35257_ (.A(_12099_),
    .B(_06812_),
    .Y(_13611_));
 sky130_fd_sc_hd__xnor2_2 _35258_ (.A(_13610_),
    .B(_13611_),
    .Y(_13612_));
 sky130_fd_sc_hd__xor2_2 _35259_ (.A(_13364_),
    .B(_13612_),
    .X(_13613_));
 sky130_fd_sc_hd__o21bai_2 _35260_ (.A1(_13607_),
    .A2(_13609_),
    .B1_N(_13613_),
    .Y(_13614_));
 sky130_fd_sc_hd__nand3b_2 _35261_ (.A_N(_13607_),
    .B(_13613_),
    .C(_13608_),
    .Y(_13615_));
 sky130_fd_sc_hd__and2_2 _35262_ (.A(_13614_),
    .B(_13615_),
    .X(_13616_));
 sky130_fd_sc_hd__a21oi_2 _35263_ (.A1(_13596_),
    .A2(_13598_),
    .B1(_13616_),
    .Y(_13617_));
 sky130_fd_sc_hd__nand3_2 _35264_ (.A(_13596_),
    .B(_13616_),
    .C(_13598_),
    .Y(_13618_));
 sky130_vsdinv _35265_ (.A(_13618_),
    .Y(_13619_));
 sky130_fd_sc_hd__nand2_2 _35266_ (.A(_13330_),
    .B(_13326_),
    .Y(_13620_));
 sky130_fd_sc_hd__o21bai_2 _35267_ (.A1(_13617_),
    .A2(_13619_),
    .B1_N(_13620_),
    .Y(_13621_));
 sky130_fd_sc_hd__nand3b_2 _35268_ (.A_N(_13617_),
    .B(_13620_),
    .C(_13618_),
    .Y(_13622_));
 sky130_vsdinv _35269_ (.A(_13362_),
    .Y(_13623_));
 sky130_fd_sc_hd__a21oi_2 _35270_ (.A1(_13382_),
    .A2(_13361_),
    .B1(_13623_),
    .Y(_13624_));
 sky130_vsdinv _35271_ (.A(_13624_),
    .Y(_13625_));
 sky130_fd_sc_hd__a21oi_2 _35272_ (.A1(_13621_),
    .A2(_13622_),
    .B1(_13625_),
    .Y(_13626_));
 sky130_fd_sc_hd__nand3_2 _35273_ (.A(_13621_),
    .B(_13622_),
    .C(_13625_),
    .Y(_13627_));
 sky130_vsdinv _35274_ (.A(_13627_),
    .Y(_13628_));
 sky130_fd_sc_hd__nor2_2 _35275_ (.A(_13626_),
    .B(_13628_),
    .Y(_13629_));
 sky130_fd_sc_hd__a21oi_2 _35276_ (.A1(_13571_),
    .A2(_13576_),
    .B1(_13629_),
    .Y(_13630_));
 sky130_fd_sc_hd__nand2_2 _35277_ (.A(_13621_),
    .B(_13622_),
    .Y(_13631_));
 sky130_fd_sc_hd__nand2_2 _35278_ (.A(_13631_),
    .B(_13624_),
    .Y(_13632_));
 sky130_fd_sc_hd__nand2_2 _35279_ (.A(_13632_),
    .B(_13627_),
    .Y(_13633_));
 sky130_fd_sc_hd__a21oi_2 _35280_ (.A1(_13573_),
    .A2(_13574_),
    .B1(_13570_),
    .Y(_13634_));
 sky130_fd_sc_hd__nor3b_2 _35281_ (.A(_13633_),
    .B(_13634_),
    .C_N(_13576_),
    .Y(_13635_));
 sky130_fd_sc_hd__o21ai_2 _35282_ (.A1(_13398_),
    .A2(_13399_),
    .B1(_13342_),
    .Y(_13636_));
 sky130_fd_sc_hd__o21bai_2 _35283_ (.A1(_13630_),
    .A2(_13635_),
    .B1_N(_13636_),
    .Y(_13637_));
 sky130_fd_sc_hd__nand2_2 _35284_ (.A(_13571_),
    .B(_13575_),
    .Y(_13638_));
 sky130_fd_sc_hd__nand2_2 _35285_ (.A(_13638_),
    .B(_13633_),
    .Y(_13639_));
 sky130_fd_sc_hd__nand3_2 _35286_ (.A(_13629_),
    .B(_13571_),
    .C(_13576_),
    .Y(_13640_));
 sky130_fd_sc_hd__nand3_2 _35287_ (.A(_13639_),
    .B(_13636_),
    .C(_13640_),
    .Y(_13641_));
 sky130_fd_sc_hd__buf_1 _35288_ (.A(_13641_),
    .X(_13642_));
 sky130_fd_sc_hd__nand2_2 _35289_ (.A(_13365_),
    .B(_13366_),
    .Y(_13643_));
 sky130_fd_sc_hd__nor2_2 _35290_ (.A(_13365_),
    .B(_13366_),
    .Y(_13644_));
 sky130_fd_sc_hd__a21oi_2 _35291_ (.A1(_13643_),
    .A2(_13363_),
    .B1(_13644_),
    .Y(_13645_));
 sky130_fd_sc_hd__nor3_2 _35292_ (.A(_13162_),
    .B(_13645_),
    .C(_13413_),
    .Y(_13646_));
 sky130_fd_sc_hd__o21ai_2 _35293_ (.A1(_13162_),
    .A2(_13413_),
    .B1(_13645_),
    .Y(_13647_));
 sky130_fd_sc_hd__nor3b_2 _35294_ (.A(_13409_),
    .B(_13646_),
    .C_N(_13647_),
    .Y(_13648_));
 sky130_vsdinv _35295_ (.A(_13646_),
    .Y(_13649_));
 sky130_fd_sc_hd__buf_1 _35296_ (.A(_13419_),
    .X(_13650_));
 sky130_fd_sc_hd__a21oi_2 _35297_ (.A1(_13649_),
    .A2(_13647_),
    .B1(_13650_),
    .Y(_13651_));
 sky130_fd_sc_hd__a21boi_2 _35298_ (.A1(_13368_),
    .A2(_13380_),
    .B1_N(_13378_),
    .Y(_13652_));
 sky130_fd_sc_hd__nor3_2 _35299_ (.A(_13648_),
    .B(_13651_),
    .C(_13652_),
    .Y(_13653_));
 sky130_fd_sc_hd__o21ai_2 _35300_ (.A1(_13648_),
    .A2(_13651_),
    .B1(_13652_),
    .Y(_13654_));
 sky130_vsdinv _35301_ (.A(_13654_),
    .Y(_13655_));
 sky130_fd_sc_hd__a21oi_2 _35302_ (.A1(_13415_),
    .A2(_13650_),
    .B1(_13414_),
    .Y(_13656_));
 sky130_vsdinv _35303_ (.A(_13656_),
    .Y(_13657_));
 sky130_fd_sc_hd__o21bai_2 _35304_ (.A1(_13653_),
    .A2(_13655_),
    .B1_N(_13657_),
    .Y(_13658_));
 sky130_fd_sc_hd__nand3b_2 _35305_ (.A_N(_13653_),
    .B(_13654_),
    .C(_13657_),
    .Y(_13659_));
 sky130_fd_sc_hd__nand2_2 _35306_ (.A(_13428_),
    .B(_13424_),
    .Y(_13660_));
 sky130_fd_sc_hd__a21oi_2 _35307_ (.A1(_13658_),
    .A2(_13659_),
    .B1(_13660_),
    .Y(_13661_));
 sky130_fd_sc_hd__nand3_2 _35308_ (.A(_13658_),
    .B(_13659_),
    .C(_13660_),
    .Y(_13662_));
 sky130_vsdinv _35309_ (.A(_13662_),
    .Y(_13663_));
 sky130_fd_sc_hd__o21bai_2 _35310_ (.A1(_13661_),
    .A2(_13663_),
    .B1_N(_13183_),
    .Y(_13664_));
 sky130_fd_sc_hd__a21o_2 _35311_ (.A1(_13658_),
    .A2(_13659_),
    .B1(_13660_),
    .X(_13665_));
 sky130_fd_sc_hd__nand3_2 _35312_ (.A(_13665_),
    .B(_12947_),
    .C(_13662_),
    .Y(_13666_));
 sky130_fd_sc_hd__nand2_2 _35313_ (.A(_13664_),
    .B(_13666_),
    .Y(_13667_));
 sky130_fd_sc_hd__a21boi_2 _35314_ (.A1(_13387_),
    .A2(_13392_),
    .B1_N(_13389_),
    .Y(_13668_));
 sky130_fd_sc_hd__nand2_2 _35315_ (.A(_13667_),
    .B(_13668_),
    .Y(_13669_));
 sky130_fd_sc_hd__nand3b_2 _35316_ (.A_N(_13668_),
    .B(_13666_),
    .C(_13664_),
    .Y(_13670_));
 sky130_fd_sc_hd__buf_1 _35317_ (.A(_13670_),
    .X(_13671_));
 sky130_vsdinv _35318_ (.A(_13431_),
    .Y(_13672_));
 sky130_fd_sc_hd__a21oi_2 _35319_ (.A1(_13430_),
    .A2(_13440_),
    .B1(_13672_),
    .Y(_13673_));
 sky130_vsdinv _35320_ (.A(_13673_),
    .Y(_13674_));
 sky130_fd_sc_hd__a21oi_2 _35321_ (.A1(_13669_),
    .A2(_13671_),
    .B1(_13674_),
    .Y(_13675_));
 sky130_fd_sc_hd__nand3_2 _35322_ (.A(_13669_),
    .B(_13670_),
    .C(_13674_),
    .Y(_13676_));
 sky130_vsdinv _35323_ (.A(_13676_),
    .Y(_13677_));
 sky130_fd_sc_hd__nor2_2 _35324_ (.A(_13675_),
    .B(_13677_),
    .Y(_13678_));
 sky130_fd_sc_hd__a21oi_2 _35325_ (.A1(_13637_),
    .A2(_13642_),
    .B1(_13678_),
    .Y(_13679_));
 sky130_fd_sc_hd__nand2_2 _35326_ (.A(_13669_),
    .B(_13671_),
    .Y(_13680_));
 sky130_fd_sc_hd__nand2_2 _35327_ (.A(_13680_),
    .B(_13673_),
    .Y(_13681_));
 sky130_fd_sc_hd__nand2_2 _35328_ (.A(_13681_),
    .B(_13676_),
    .Y(_13682_));
 sky130_fd_sc_hd__a21oi_2 _35329_ (.A1(_13639_),
    .A2(_13640_),
    .B1(_13636_),
    .Y(_13683_));
 sky130_vsdinv _35330_ (.A(_13642_),
    .Y(_13684_));
 sky130_fd_sc_hd__nor3_2 _35331_ (.A(_13682_),
    .B(_13683_),
    .C(_13684_),
    .Y(_13685_));
 sky130_fd_sc_hd__o21ai_2 _35332_ (.A1(_13445_),
    .A2(_13447_),
    .B1(_13407_),
    .Y(_13686_));
 sky130_fd_sc_hd__o21bai_2 _35333_ (.A1(_13679_),
    .A2(_13685_),
    .B1_N(_13686_),
    .Y(_13687_));
 sky130_fd_sc_hd__nand2_2 _35334_ (.A(_13637_),
    .B(_13641_),
    .Y(_13688_));
 sky130_fd_sc_hd__nand2_2 _35335_ (.A(_13688_),
    .B(_13682_),
    .Y(_13689_));
 sky130_fd_sc_hd__nand3_2 _35336_ (.A(_13678_),
    .B(_13637_),
    .C(_13642_),
    .Y(_13690_));
 sky130_fd_sc_hd__nand3_2 _35337_ (.A(_13689_),
    .B(_13686_),
    .C(_13690_),
    .Y(_13691_));
 sky130_fd_sc_hd__nand2_2 _35338_ (.A(_13687_),
    .B(_13691_),
    .Y(_13692_));
 sky130_fd_sc_hd__buf_1 _35339_ (.A(_13212_),
    .X(_13693_));
 sky130_fd_sc_hd__nand2_2 _35340_ (.A(_13443_),
    .B(_13438_),
    .Y(_13694_));
 sky130_fd_sc_hd__xor2_2 _35341_ (.A(_13693_),
    .B(_13694_),
    .X(_13695_));
 sky130_vsdinv _35342_ (.A(_13695_),
    .Y(_13696_));
 sky130_fd_sc_hd__nand2_2 _35343_ (.A(_13692_),
    .B(_13696_),
    .Y(_13697_));
 sky130_fd_sc_hd__buf_1 _35344_ (.A(_13691_),
    .X(_13698_));
 sky130_fd_sc_hd__nand3_2 _35345_ (.A(_13687_),
    .B(_13695_),
    .C(_13698_),
    .Y(_13699_));
 sky130_vsdinv _35346_ (.A(_13459_),
    .Y(_13700_));
 sky130_fd_sc_hd__a21oi_2 _35347_ (.A1(_13452_),
    .A2(_13453_),
    .B1(_13450_),
    .Y(_13701_));
 sky130_fd_sc_hd__o21ai_2 _35348_ (.A1(_13700_),
    .A2(_13701_),
    .B1(_13455_),
    .Y(_13702_));
 sky130_fd_sc_hd__a21oi_2 _35349_ (.A1(_13697_),
    .A2(_13699_),
    .B1(_13702_),
    .Y(_13703_));
 sky130_fd_sc_hd__a21oi_2 _35350_ (.A1(_13687_),
    .A2(_13698_),
    .B1(_13695_),
    .Y(_13704_));
 sky130_fd_sc_hd__a21boi_2 _35351_ (.A1(_13451_),
    .A2(_13459_),
    .B1_N(_13455_),
    .Y(_13705_));
 sky130_fd_sc_hd__a21oi_2 _35352_ (.A1(_13689_),
    .A2(_13690_),
    .B1(_13686_),
    .Y(_13706_));
 sky130_vsdinv _35353_ (.A(_13698_),
    .Y(_13707_));
 sky130_fd_sc_hd__nor3_2 _35354_ (.A(_13696_),
    .B(_13706_),
    .C(_13707_),
    .Y(_13708_));
 sky130_fd_sc_hd__nor3_2 _35355_ (.A(_13704_),
    .B(_13705_),
    .C(_13708_),
    .Y(_13709_));
 sky130_fd_sc_hd__buf_1 _35356_ (.A(_13457_),
    .X(_13710_));
 sky130_fd_sc_hd__o21bai_2 _35357_ (.A1(_13703_),
    .A2(_13709_),
    .B1_N(_13710_),
    .Y(_13711_));
 sky130_fd_sc_hd__o21bai_2 _35358_ (.A1(_13704_),
    .A2(_13708_),
    .B1_N(_13702_),
    .Y(_13712_));
 sky130_fd_sc_hd__nand3_2 _35359_ (.A(_13697_),
    .B(_13702_),
    .C(_13699_),
    .Y(_13713_));
 sky130_fd_sc_hd__nand3_2 _35360_ (.A(_13712_),
    .B(_13710_),
    .C(_13713_),
    .Y(_13714_));
 sky130_vsdinv _35361_ (.A(_13469_),
    .Y(_13715_));
 sky130_fd_sc_hd__a21oi_2 _35362_ (.A1(_13465_),
    .A2(_13461_),
    .B1(_13463_),
    .Y(_13716_));
 sky130_fd_sc_hd__o21ai_2 _35363_ (.A1(_13715_),
    .A2(_13716_),
    .B1(_13466_),
    .Y(_13717_));
 sky130_fd_sc_hd__a21oi_2 _35364_ (.A1(_13711_),
    .A2(_13714_),
    .B1(_13717_),
    .Y(_13718_));
 sky130_fd_sc_hd__nand3_2 _35365_ (.A(_13711_),
    .B(_13717_),
    .C(_13714_),
    .Y(_13719_));
 sky130_vsdinv _35366_ (.A(_13719_),
    .Y(_13720_));
 sky130_fd_sc_hd__nor2_2 _35367_ (.A(_13718_),
    .B(_13720_),
    .Y(_13721_));
 sky130_fd_sc_hd__a21oi_2 _35368_ (.A1(_13475_),
    .A2(_13471_),
    .B1(_13473_),
    .Y(_13722_));
 sky130_fd_sc_hd__a21oi_2 _35369_ (.A1(_13237_),
    .A2(_13476_),
    .B1(_13722_),
    .Y(_13723_));
 sky130_vsdinv _35370_ (.A(_13723_),
    .Y(_13724_));
 sky130_fd_sc_hd__o31ai_2 _35371_ (.A1(_13238_),
    .A2(_13477_),
    .A3(_13247_),
    .B1(_13724_),
    .Y(_13725_));
 sky130_fd_sc_hd__xor2_2 _35372_ (.A(_13721_),
    .B(_13725_),
    .X(_02661_));
 sky130_fd_sc_hd__nand2_2 _35373_ (.A(_10486_),
    .B(_06186_),
    .Y(_13726_));
 sky130_fd_sc_hd__nand3b_2 _35374_ (.A_N(_13726_),
    .B(_12183_),
    .C(_19249_),
    .Y(_13727_));
 sky130_fd_sc_hd__o21ai_2 _35375_ (.A1(_07060_),
    .A2(_11324_),
    .B1(_13726_),
    .Y(_13728_));
 sky130_fd_sc_hd__and2_2 _35376_ (.A(_10483_),
    .B(_08181_),
    .X(_13729_));
 sky130_fd_sc_hd__a21o_2 _35377_ (.A1(_13727_),
    .A2(_13728_),
    .B1(_13729_),
    .X(_13730_));
 sky130_fd_sc_hd__nand3_2 _35378_ (.A(_13727_),
    .B(_13729_),
    .C(_13728_),
    .Y(_13731_));
 sky130_fd_sc_hd__nand2_2 _35379_ (.A(_13484_),
    .B(_13480_),
    .Y(_13732_));
 sky130_fd_sc_hd__a21o_2 _35380_ (.A1(_13730_),
    .A2(_13731_),
    .B1(_13732_),
    .X(_13733_));
 sky130_fd_sc_hd__nand3_2 _35381_ (.A(_13732_),
    .B(_13730_),
    .C(_13731_),
    .Y(_13734_));
 sky130_fd_sc_hd__and2_2 _35382_ (.A(_09605_),
    .B(_08254_),
    .X(_13735_));
 sky130_fd_sc_hd__buf_1 _35383_ (.A(_13735_),
    .X(_13736_));
 sky130_fd_sc_hd__nand2_2 _35384_ (.A(_11011_),
    .B(_07688_),
    .Y(_13737_));
 sky130_fd_sc_hd__nand2_2 _35385_ (.A(_10253_),
    .B(_06595_),
    .Y(_13738_));
 sky130_fd_sc_hd__xnor2_2 _35386_ (.A(_13737_),
    .B(_13738_),
    .Y(_13739_));
 sky130_fd_sc_hd__xnor2_2 _35387_ (.A(_13736_),
    .B(_13739_),
    .Y(_13740_));
 sky130_fd_sc_hd__a21oi_2 _35388_ (.A1(_13733_),
    .A2(_13734_),
    .B1(_13740_),
    .Y(_13741_));
 sky130_fd_sc_hd__nand3_2 _35389_ (.A(_13733_),
    .B(_13740_),
    .C(_13734_),
    .Y(_13742_));
 sky130_vsdinv _35390_ (.A(_13742_),
    .Y(_13743_));
 sky130_fd_sc_hd__o21ai_2 _35391_ (.A1(_13494_),
    .A2(_13495_),
    .B1(_13487_),
    .Y(_13744_));
 sky130_fd_sc_hd__o21bai_2 _35392_ (.A1(_13741_),
    .A2(_13743_),
    .B1_N(_13744_),
    .Y(_13745_));
 sky130_fd_sc_hd__a21o_2 _35393_ (.A1(_13733_),
    .A2(_13734_),
    .B1(_13740_),
    .X(_13746_));
 sky130_fd_sc_hd__nand3_2 _35394_ (.A(_13746_),
    .B(_13742_),
    .C(_13744_),
    .Y(_13747_));
 sky130_fd_sc_hd__nand2_2 _35395_ (.A(_09587_),
    .B(_19211_),
    .Y(_13748_));
 sky130_fd_sc_hd__nand2_2 _35396_ (.A(_09305_),
    .B(_19207_),
    .Y(_13749_));
 sky130_fd_sc_hd__xor2_2 _35397_ (.A(_13748_),
    .B(_13749_),
    .X(_13750_));
 sky130_fd_sc_hd__nand3_2 _35398_ (.A(_13750_),
    .B(_13026_),
    .C(_08304_),
    .Y(_13751_));
 sky130_fd_sc_hd__xnor2_2 _35399_ (.A(_13748_),
    .B(_13749_),
    .Y(_13752_));
 sky130_fd_sc_hd__o21ai_2 _35400_ (.A1(_18741_),
    .A2(_09665_),
    .B1(_13752_),
    .Y(_13753_));
 sky130_fd_sc_hd__a22oi_2 _35401_ (.A1(_11618_),
    .A2(_07100_),
    .B1(_18717_),
    .B2(_06607_),
    .Y(_13754_));
 sky130_fd_sc_hd__nor2_2 _35402_ (.A(_13489_),
    .B(_13490_),
    .Y(_13755_));
 sky130_vsdinv _35403_ (.A(_13755_),
    .Y(_13756_));
 sky130_fd_sc_hd__o31a_2 _35404_ (.A1(_18724_),
    .A2(_19226_),
    .A3(_13754_),
    .B1(_13756_),
    .X(_13757_));
 sky130_fd_sc_hd__a21boi_2 _35405_ (.A1(_13751_),
    .A2(_13753_),
    .B1_N(_13757_),
    .Y(_13758_));
 sky130_fd_sc_hd__nand3b_2 _35406_ (.A_N(_13757_),
    .B(_13753_),
    .C(_13751_),
    .Y(_13759_));
 sky130_vsdinv _35407_ (.A(_13759_),
    .Y(_13760_));
 sky130_fd_sc_hd__nand3b_2 _35408_ (.A_N(_13505_),
    .B(_18736_),
    .C(_11110_),
    .Y(_13761_));
 sky130_fd_sc_hd__o31a_2 _35409_ (.A1(_11036_),
    .A2(_19209_),
    .A3(_13510_),
    .B1(_13761_),
    .X(_13762_));
 sky130_fd_sc_hd__o21ai_2 _35410_ (.A1(_13758_),
    .A2(_13760_),
    .B1(_13762_),
    .Y(_13763_));
 sky130_vsdinv _35411_ (.A(_13762_),
    .Y(_13764_));
 sky130_fd_sc_hd__a21bo_2 _35412_ (.A1(_13753_),
    .A2(_13751_),
    .B1_N(_13757_),
    .X(_13765_));
 sky130_fd_sc_hd__nand3_2 _35413_ (.A(_13764_),
    .B(_13765_),
    .C(_13759_),
    .Y(_13766_));
 sky130_fd_sc_hd__nand2_2 _35414_ (.A(_13763_),
    .B(_13766_),
    .Y(_13767_));
 sky130_fd_sc_hd__buf_1 _35415_ (.A(_13767_),
    .X(_13768_));
 sky130_fd_sc_hd__a21boi_2 _35416_ (.A1(_13745_),
    .A2(_13747_),
    .B1_N(_13768_),
    .Y(_13769_));
 sky130_fd_sc_hd__a21oi_2 _35417_ (.A1(_13746_),
    .A2(_13742_),
    .B1(_13744_),
    .Y(_13770_));
 sky130_vsdinv _35418_ (.A(_13747_),
    .Y(_13771_));
 sky130_fd_sc_hd__nor3_2 _35419_ (.A(_13768_),
    .B(_13770_),
    .C(_13771_),
    .Y(_13772_));
 sky130_fd_sc_hd__o21ai_2 _35420_ (.A1(_13524_),
    .A2(_13525_),
    .B1(_13504_),
    .Y(_13773_));
 sky130_fd_sc_hd__o21bai_2 _35421_ (.A1(_13769_),
    .A2(_13772_),
    .B1_N(_13773_),
    .Y(_13774_));
 sky130_fd_sc_hd__o21ai_2 _35422_ (.A1(_13770_),
    .A2(_13771_),
    .B1(_13768_),
    .Y(_13775_));
 sky130_fd_sc_hd__nand3b_2 _35423_ (.A_N(_13767_),
    .B(_13747_),
    .C(_13745_),
    .Y(_13776_));
 sky130_fd_sc_hd__nand3_2 _35424_ (.A(_13775_),
    .B(_13776_),
    .C(_13773_),
    .Y(_13777_));
 sky130_fd_sc_hd__buf_1 _35425_ (.A(_13777_),
    .X(_13778_));
 sky130_fd_sc_hd__nand2_2 _35426_ (.A(_10421_),
    .B(_10159_),
    .Y(_13779_));
 sky130_fd_sc_hd__nand2_2 _35427_ (.A(_08473_),
    .B(_11136_),
    .Y(_13780_));
 sky130_fd_sc_hd__nor2_2 _35428_ (.A(_13779_),
    .B(_13780_),
    .Y(_13781_));
 sky130_fd_sc_hd__and2_2 _35429_ (.A(_08084_),
    .B(_09216_),
    .X(_13782_));
 sky130_vsdinv _35430_ (.A(_13782_),
    .Y(_13783_));
 sky130_fd_sc_hd__nand2_2 _35431_ (.A(_13779_),
    .B(_13780_),
    .Y(_13784_));
 sky130_fd_sc_hd__nor3b_2 _35432_ (.A(_13781_),
    .B(_13783_),
    .C_N(_13784_),
    .Y(_13785_));
 sky130_vsdinv _35433_ (.A(_13785_),
    .Y(_13786_));
 sky130_fd_sc_hd__buf_1 _35434_ (.A(_08571_),
    .X(_13787_));
 sky130_fd_sc_hd__nand3b_2 _35435_ (.A_N(_13779_),
    .B(_12791_),
    .C(_13787_),
    .Y(_13788_));
 sky130_fd_sc_hd__o2bb2ai_2 _35436_ (.A1_N(_13784_),
    .A2_N(_13788_),
    .B1(_13050_),
    .B2(_19188_),
    .Y(_13789_));
 sky130_fd_sc_hd__a21boi_2 _35437_ (.A1(_13535_),
    .A2(_13539_),
    .B1_N(_13537_),
    .Y(_13790_));
 sky130_vsdinv _35438_ (.A(_13790_),
    .Y(_13791_));
 sky130_fd_sc_hd__a21o_2 _35439_ (.A1(_13786_),
    .A2(_13789_),
    .B1(_13791_),
    .X(_13792_));
 sky130_fd_sc_hd__nand3_2 _35440_ (.A(_13791_),
    .B(_13786_),
    .C(_13789_),
    .Y(_13793_));
 sky130_fd_sc_hd__and2_2 _35441_ (.A(_07421_),
    .B(_11736_),
    .X(_13794_));
 sky130_fd_sc_hd__nand2_2 _35442_ (.A(_10745_),
    .B(_08295_),
    .Y(_13795_));
 sky130_fd_sc_hd__nand2_2 _35443_ (.A(_12254_),
    .B(_11433_),
    .Y(_13796_));
 sky130_fd_sc_hd__xnor2_2 _35444_ (.A(_13795_),
    .B(_13796_),
    .Y(_13797_));
 sky130_fd_sc_hd__xnor2_2 _35445_ (.A(_13794_),
    .B(_13797_),
    .Y(_13798_));
 sky130_fd_sc_hd__a21oi_2 _35446_ (.A1(_13792_),
    .A2(_13793_),
    .B1(_13798_),
    .Y(_13799_));
 sky130_fd_sc_hd__nand3_2 _35447_ (.A(_13792_),
    .B(_13798_),
    .C(_13793_),
    .Y(_13800_));
 sky130_vsdinv _35448_ (.A(_13800_),
    .Y(_13801_));
 sky130_fd_sc_hd__a21o_2 _35449_ (.A1(_13513_),
    .A2(_13515_),
    .B1(_13522_),
    .X(_13802_));
 sky130_fd_sc_hd__o21bai_2 _35450_ (.A1(_13799_),
    .A2(_13801_),
    .B1_N(_13802_),
    .Y(_13803_));
 sky130_fd_sc_hd__a21o_2 _35451_ (.A1(_13792_),
    .A2(_13793_),
    .B1(_13798_),
    .X(_13804_));
 sky130_fd_sc_hd__nand3_2 _35452_ (.A(_13804_),
    .B(_13802_),
    .C(_13800_),
    .Y(_13805_));
 sky130_vsdinv _35453_ (.A(_13545_),
    .Y(_13806_));
 sky130_fd_sc_hd__a21oi_2 _35454_ (.A1(_13544_),
    .A2(_13551_),
    .B1(_13806_),
    .Y(_13807_));
 sky130_vsdinv _35455_ (.A(_13807_),
    .Y(_13808_));
 sky130_fd_sc_hd__a21oi_2 _35456_ (.A1(_13803_),
    .A2(_13805_),
    .B1(_13808_),
    .Y(_13809_));
 sky130_fd_sc_hd__nand3_2 _35457_ (.A(_13803_),
    .B(_13808_),
    .C(_13805_),
    .Y(_13810_));
 sky130_vsdinv _35458_ (.A(_13810_),
    .Y(_13811_));
 sky130_fd_sc_hd__nor2_2 _35459_ (.A(_13809_),
    .B(_13811_),
    .Y(_13812_));
 sky130_fd_sc_hd__a21oi_2 _35460_ (.A1(_13774_),
    .A2(_13778_),
    .B1(_13812_),
    .Y(_13813_));
 sky130_fd_sc_hd__nand2_2 _35461_ (.A(_13803_),
    .B(_13805_),
    .Y(_13814_));
 sky130_fd_sc_hd__nand2_2 _35462_ (.A(_13814_),
    .B(_13807_),
    .Y(_13815_));
 sky130_fd_sc_hd__nand2_2 _35463_ (.A(_13815_),
    .B(_13810_),
    .Y(_13816_));
 sky130_fd_sc_hd__a21oi_2 _35464_ (.A1(_13775_),
    .A2(_13776_),
    .B1(_13773_),
    .Y(_13817_));
 sky130_vsdinv _35465_ (.A(_13778_),
    .Y(_13818_));
 sky130_fd_sc_hd__nor3_2 _35466_ (.A(_13816_),
    .B(_13817_),
    .C(_13818_),
    .Y(_13819_));
 sky130_fd_sc_hd__o21ai_2 _35467_ (.A1(_13565_),
    .A2(_13567_),
    .B1(_13534_),
    .Y(_13820_));
 sky130_fd_sc_hd__o21bai_2 _35468_ (.A1(_13813_),
    .A2(_13819_),
    .B1_N(_13820_),
    .Y(_13821_));
 sky130_fd_sc_hd__nand2_2 _35469_ (.A(_13774_),
    .B(_13777_),
    .Y(_13822_));
 sky130_fd_sc_hd__nand2_2 _35470_ (.A(_13822_),
    .B(_13816_),
    .Y(_13823_));
 sky130_fd_sc_hd__nand3_2 _35471_ (.A(_13812_),
    .B(_13778_),
    .C(_13774_),
    .Y(_13824_));
 sky130_fd_sc_hd__nand3_2 _35472_ (.A(_13823_),
    .B(_13824_),
    .C(_13820_),
    .Y(_13825_));
 sky130_fd_sc_hd__buf_1 _35473_ (.A(_13825_),
    .X(_13826_));
 sky130_fd_sc_hd__nand2_2 _35474_ (.A(_07469_),
    .B(_10537_),
    .Y(_13827_));
 sky130_fd_sc_hd__nand2_2 _35475_ (.A(_07470_),
    .B(_19156_),
    .Y(_13828_));
 sky130_fd_sc_hd__xor2_2 _35476_ (.A(_13827_),
    .B(_13828_),
    .X(_13829_));
 sky130_fd_sc_hd__buf_1 _35477_ (.A(_19149_),
    .X(_13830_));
 sky130_fd_sc_hd__buf_1 _35478_ (.A(_13830_),
    .X(_13831_));
 sky130_fd_sc_hd__nand3_2 _35479_ (.A(_13829_),
    .B(_13089_),
    .C(_13831_),
    .Y(_13832_));
 sky130_fd_sc_hd__xnor2_2 _35480_ (.A(_13827_),
    .B(_13828_),
    .Y(_13833_));
 sky130_fd_sc_hd__o21ai_2 _35481_ (.A1(_11716_),
    .A2(_19151_),
    .B1(_13833_),
    .Y(_13834_));
 sky130_fd_sc_hd__nand2_2 _35482_ (.A(_13832_),
    .B(_13834_),
    .Y(_13835_));
 sky130_fd_sc_hd__a21boi_2 _35483_ (.A1(_13549_),
    .A2(_13546_),
    .B1_N(_13548_),
    .Y(_13836_));
 sky130_fd_sc_hd__nand2_2 _35484_ (.A(_13835_),
    .B(_13836_),
    .Y(_13837_));
 sky130_fd_sc_hd__nand3b_2 _35485_ (.A_N(_13836_),
    .B(_13832_),
    .C(_13834_),
    .Y(_13838_));
 sky130_fd_sc_hd__nand2_2 _35486_ (.A(_13837_),
    .B(_13838_),
    .Y(_13839_));
 sky130_fd_sc_hd__o21a_2 _35487_ (.A1(_13577_),
    .A2(_13578_),
    .B1(_13581_),
    .X(_13840_));
 sky130_fd_sc_hd__nand2_2 _35488_ (.A(_13839_),
    .B(_13840_),
    .Y(_13841_));
 sky130_fd_sc_hd__nand3b_2 _35489_ (.A_N(_13840_),
    .B(_13838_),
    .C(_13837_),
    .Y(_13842_));
 sky130_fd_sc_hd__nand2_2 _35490_ (.A(_13593_),
    .B(_13589_),
    .Y(_13843_));
 sky130_fd_sc_hd__a21o_2 _35491_ (.A1(_13841_),
    .A2(_13842_),
    .B1(_13843_),
    .X(_13844_));
 sky130_fd_sc_hd__nand3_2 _35492_ (.A(_13843_),
    .B(_13841_),
    .C(_13842_),
    .Y(_13845_));
 sky130_fd_sc_hd__o21ai_2 _35493_ (.A1(_13599_),
    .A2(_13600_),
    .B1(_13603_),
    .Y(_13846_));
 sky130_fd_sc_hd__nand2_2 _35494_ (.A(_07190_),
    .B(_10554_),
    .Y(_13847_));
 sky130_fd_sc_hd__nand2_2 _35495_ (.A(_06392_),
    .B(_19138_),
    .Y(_13848_));
 sky130_fd_sc_hd__xnor2_2 _35496_ (.A(_13847_),
    .B(_13848_),
    .Y(_13849_));
 sky130_fd_sc_hd__o21ai_2 _35497_ (.A1(_11745_),
    .A2(_12389_),
    .B1(_13849_),
    .Y(_13850_));
 sky130_fd_sc_hd__xor2_2 _35498_ (.A(_13847_),
    .B(_13848_),
    .X(_13851_));
 sky130_fd_sc_hd__and2_2 _35499_ (.A(_10382_),
    .B(_10540_),
    .X(_13852_));
 sky130_fd_sc_hd__nand2_2 _35500_ (.A(_13851_),
    .B(_13852_),
    .Y(_13853_));
 sky130_fd_sc_hd__nand3_2 _35501_ (.A(_13846_),
    .B(_13850_),
    .C(_13853_),
    .Y(_13854_));
 sky130_fd_sc_hd__nand2_2 _35502_ (.A(_13853_),
    .B(_13850_),
    .Y(_13855_));
 sky130_fd_sc_hd__o211ai_2 _35503_ (.A1(_13599_),
    .A2(_13600_),
    .B1(_13603_),
    .C1(_13855_),
    .Y(_13856_));
 sky130_fd_sc_hd__o21ai_2 _35504_ (.A1(_06147_),
    .A2(_06673_),
    .B1(_11830_),
    .Y(_13857_));
 sky130_fd_sc_hd__nand3_2 _35505_ (.A(_10881_),
    .B(_06810_),
    .C(_07377_),
    .Y(_13858_));
 sky130_vsdinv _35506_ (.A(_13858_),
    .Y(_13859_));
 sky130_fd_sc_hd__nor3b_2 _35507_ (.A(_13857_),
    .B(_13859_),
    .C_N(_13363_),
    .Y(_13860_));
 sky130_fd_sc_hd__o21a_2 _35508_ (.A1(_13857_),
    .A2(_13859_),
    .B1(_13364_),
    .X(_13861_));
 sky130_fd_sc_hd__o2bb2ai_2 _35509_ (.A1_N(_13854_),
    .A2_N(_13856_),
    .B1(_13860_),
    .B2(_13861_),
    .Y(_13862_));
 sky130_fd_sc_hd__nor2_2 _35510_ (.A(_13861_),
    .B(_13860_),
    .Y(_13863_));
 sky130_fd_sc_hd__buf_1 _35511_ (.A(_13863_),
    .X(_13864_));
 sky130_fd_sc_hd__nand3_2 _35512_ (.A(_13856_),
    .B(_13854_),
    .C(_13864_),
    .Y(_13865_));
 sky130_fd_sc_hd__and2_2 _35513_ (.A(_13862_),
    .B(_13865_),
    .X(_13866_));
 sky130_fd_sc_hd__a21oi_2 _35514_ (.A1(_13844_),
    .A2(_13845_),
    .B1(_13866_),
    .Y(_13867_));
 sky130_fd_sc_hd__nand3_2 _35515_ (.A(_13844_),
    .B(_13866_),
    .C(_13845_),
    .Y(_13868_));
 sky130_vsdinv _35516_ (.A(_13868_),
    .Y(_13869_));
 sky130_fd_sc_hd__o21ai_2 _35517_ (.A1(_13559_),
    .A2(_13556_),
    .B1(_13562_),
    .Y(_13870_));
 sky130_fd_sc_hd__o21bai_2 _35518_ (.A1(_13867_),
    .A2(_13869_),
    .B1_N(_13870_),
    .Y(_13871_));
 sky130_fd_sc_hd__a21o_2 _35519_ (.A1(_13844_),
    .A2(_13845_),
    .B1(_13866_),
    .X(_13872_));
 sky130_fd_sc_hd__nand3_2 _35520_ (.A(_13872_),
    .B(_13870_),
    .C(_13868_),
    .Y(_13873_));
 sky130_fd_sc_hd__nand2_2 _35521_ (.A(_13871_),
    .B(_13873_),
    .Y(_13874_));
 sky130_fd_sc_hd__a21boi_2 _35522_ (.A1(_13596_),
    .A2(_13616_),
    .B1_N(_13598_),
    .Y(_13875_));
 sky130_fd_sc_hd__nand2_2 _35523_ (.A(_13874_),
    .B(_13875_),
    .Y(_13876_));
 sky130_vsdinv _35524_ (.A(_13875_),
    .Y(_13877_));
 sky130_fd_sc_hd__nand3_2 _35525_ (.A(_13871_),
    .B(_13877_),
    .C(_13873_),
    .Y(_13878_));
 sky130_fd_sc_hd__nand2_2 _35526_ (.A(_13876_),
    .B(_13878_),
    .Y(_13879_));
 sky130_fd_sc_hd__buf_1 _35527_ (.A(_13879_),
    .X(_13880_));
 sky130_fd_sc_hd__a21boi_2 _35528_ (.A1(_13821_),
    .A2(_13826_),
    .B1_N(_13880_),
    .Y(_13881_));
 sky130_fd_sc_hd__a21oi_2 _35529_ (.A1(_13823_),
    .A2(_13824_),
    .B1(_13820_),
    .Y(_13882_));
 sky130_fd_sc_hd__nor3b_2 _35530_ (.A(_13880_),
    .B(_13882_),
    .C_N(_13826_),
    .Y(_13883_));
 sky130_fd_sc_hd__o21ai_2 _35531_ (.A1(_13633_),
    .A2(_13634_),
    .B1(_13576_),
    .Y(_13884_));
 sky130_fd_sc_hd__o21bai_2 _35532_ (.A1(_13881_),
    .A2(_13883_),
    .B1_N(_13884_),
    .Y(_13885_));
 sky130_fd_sc_hd__nand2_2 _35533_ (.A(_13821_),
    .B(_13825_),
    .Y(_13886_));
 sky130_fd_sc_hd__nand2_2 _35534_ (.A(_13886_),
    .B(_13880_),
    .Y(_13887_));
 sky130_fd_sc_hd__nand3b_2 _35535_ (.A_N(_13879_),
    .B(_13826_),
    .C(_13821_),
    .Y(_13888_));
 sky130_fd_sc_hd__nand3_2 _35536_ (.A(_13887_),
    .B(_13888_),
    .C(_13884_),
    .Y(_13889_));
 sky130_fd_sc_hd__buf_1 _35537_ (.A(_13889_),
    .X(_13890_));
 sky130_fd_sc_hd__nand2_2 _35538_ (.A(_13610_),
    .B(_13611_),
    .Y(_13891_));
 sky130_fd_sc_hd__nor2_2 _35539_ (.A(_13610_),
    .B(_13611_),
    .Y(_13892_));
 sky130_fd_sc_hd__a21oi_2 _35540_ (.A1(_13891_),
    .A2(_13363_),
    .B1(_13892_),
    .Y(_13893_));
 sky130_fd_sc_hd__nor3_2 _35541_ (.A(_13162_),
    .B(_13893_),
    .C(_13413_),
    .Y(_13894_));
 sky130_vsdinv _35542_ (.A(_13894_),
    .Y(_13895_));
 sky130_fd_sc_hd__o21ai_2 _35543_ (.A1(_13161_),
    .A2(_13163_),
    .B1(_13893_),
    .Y(_13896_));
 sky130_fd_sc_hd__a21oi_2 _35544_ (.A1(_13895_),
    .A2(_13896_),
    .B1(_13419_),
    .Y(_13897_));
 sky130_fd_sc_hd__nand2_2 _35545_ (.A(_13615_),
    .B(_13608_),
    .Y(_13898_));
 sky130_fd_sc_hd__nor3b_2 _35546_ (.A(_13409_),
    .B(_13894_),
    .C_N(_13896_),
    .Y(_13899_));
 sky130_vsdinv _35547_ (.A(_13899_),
    .Y(_13900_));
 sky130_fd_sc_hd__nand3b_2 _35548_ (.A_N(_13897_),
    .B(_13898_),
    .C(_13900_),
    .Y(_13901_));
 sky130_fd_sc_hd__o211ai_2 _35549_ (.A1(_13899_),
    .A2(_13897_),
    .B1(_13608_),
    .C1(_13615_),
    .Y(_13902_));
 sky130_fd_sc_hd__a21oi_2 _35550_ (.A1(_13647_),
    .A2(_13650_),
    .B1(_13646_),
    .Y(_13903_));
 sky130_vsdinv _35551_ (.A(_13903_),
    .Y(_13904_));
 sky130_fd_sc_hd__a21oi_2 _35552_ (.A1(_13901_),
    .A2(_13902_),
    .B1(_13904_),
    .Y(_13905_));
 sky130_fd_sc_hd__nand3_2 _35553_ (.A(_13901_),
    .B(_13902_),
    .C(_13904_),
    .Y(_13906_));
 sky130_vsdinv _35554_ (.A(_13906_),
    .Y(_13907_));
 sky130_fd_sc_hd__a21o_2 _35555_ (.A1(_13654_),
    .A2(_13657_),
    .B1(_13653_),
    .X(_13908_));
 sky130_fd_sc_hd__o21bai_2 _35556_ (.A1(_13905_),
    .A2(_13907_),
    .B1_N(_13908_),
    .Y(_13909_));
 sky130_fd_sc_hd__nand3b_2 _35557_ (.A_N(_13905_),
    .B(_13906_),
    .C(_13908_),
    .Y(_13910_));
 sky130_fd_sc_hd__a21oi_2 _35558_ (.A1(_13909_),
    .A2(_13910_),
    .B1(_13184_),
    .Y(_13911_));
 sky130_fd_sc_hd__nand3_2 _35559_ (.A(_13909_),
    .B(_13910_),
    .C(_13432_),
    .Y(_13912_));
 sky130_vsdinv _35560_ (.A(_13912_),
    .Y(_13913_));
 sky130_fd_sc_hd__a21boi_2 _35561_ (.A1(_13621_),
    .A2(_13625_),
    .B1_N(_13622_),
    .Y(_13914_));
 sky130_fd_sc_hd__o21ai_2 _35562_ (.A1(_13911_),
    .A2(_13913_),
    .B1(_13914_),
    .Y(_13915_));
 sky130_fd_sc_hd__a21o_2 _35563_ (.A1(_13909_),
    .A2(_13910_),
    .B1(_13183_),
    .X(_13916_));
 sky130_fd_sc_hd__nand3b_2 _35564_ (.A_N(_13914_),
    .B(_13912_),
    .C(_13916_),
    .Y(_13917_));
 sky130_fd_sc_hd__buf_1 _35565_ (.A(_13917_),
    .X(_13918_));
 sky130_fd_sc_hd__a21oi_2 _35566_ (.A1(_13665_),
    .A2(_13184_),
    .B1(_13663_),
    .Y(_13919_));
 sky130_vsdinv _35567_ (.A(_13919_),
    .Y(_13920_));
 sky130_fd_sc_hd__a21oi_2 _35568_ (.A1(_13915_),
    .A2(_13918_),
    .B1(_13920_),
    .Y(_13921_));
 sky130_fd_sc_hd__nand3_2 _35569_ (.A(_13915_),
    .B(_13917_),
    .C(_13920_),
    .Y(_13922_));
 sky130_vsdinv _35570_ (.A(_13922_),
    .Y(_13923_));
 sky130_fd_sc_hd__nor2_2 _35571_ (.A(_13921_),
    .B(_13923_),
    .Y(_13924_));
 sky130_fd_sc_hd__a21oi_2 _35572_ (.A1(_13885_),
    .A2(_13890_),
    .B1(_13924_),
    .Y(_13925_));
 sky130_fd_sc_hd__nand2_2 _35573_ (.A(_13915_),
    .B(_13918_),
    .Y(_13926_));
 sky130_fd_sc_hd__nand2_2 _35574_ (.A(_13926_),
    .B(_13919_),
    .Y(_13927_));
 sky130_fd_sc_hd__nand2_2 _35575_ (.A(_13927_),
    .B(_13922_),
    .Y(_13928_));
 sky130_fd_sc_hd__a21oi_2 _35576_ (.A1(_13887_),
    .A2(_13888_),
    .B1(_13884_),
    .Y(_13929_));
 sky130_vsdinv _35577_ (.A(_13890_),
    .Y(_13930_));
 sky130_fd_sc_hd__nor3_2 _35578_ (.A(_13928_),
    .B(_13929_),
    .C(_13930_),
    .Y(_13931_));
 sky130_fd_sc_hd__o21ai_2 _35579_ (.A1(_13682_),
    .A2(_13683_),
    .B1(_13642_),
    .Y(_13932_));
 sky130_fd_sc_hd__o21bai_2 _35580_ (.A1(_13925_),
    .A2(_13931_),
    .B1_N(_13932_),
    .Y(_13933_));
 sky130_fd_sc_hd__nand2_2 _35581_ (.A(_13885_),
    .B(_13889_),
    .Y(_13934_));
 sky130_fd_sc_hd__nand2_2 _35582_ (.A(_13934_),
    .B(_13928_),
    .Y(_13935_));
 sky130_fd_sc_hd__nand3_2 _35583_ (.A(_13924_),
    .B(_13885_),
    .C(_13890_),
    .Y(_13936_));
 sky130_fd_sc_hd__nand3_2 _35584_ (.A(_13935_),
    .B(_13936_),
    .C(_13932_),
    .Y(_13937_));
 sky130_fd_sc_hd__buf_1 _35585_ (.A(_13937_),
    .X(_13938_));
 sky130_fd_sc_hd__nand2_2 _35586_ (.A(_13676_),
    .B(_13671_),
    .Y(_13939_));
 sky130_fd_sc_hd__xor2_2 _35587_ (.A(_13213_),
    .B(_13939_),
    .X(_13940_));
 sky130_fd_sc_hd__a21oi_2 _35588_ (.A1(_13933_),
    .A2(_13938_),
    .B1(_13940_),
    .Y(_13941_));
 sky130_vsdinv _35589_ (.A(_13940_),
    .Y(_13942_));
 sky130_fd_sc_hd__a21oi_2 _35590_ (.A1(_13935_),
    .A2(_13936_),
    .B1(_13932_),
    .Y(_13943_));
 sky130_vsdinv _35591_ (.A(_13938_),
    .Y(_13944_));
 sky130_fd_sc_hd__nor3_2 _35592_ (.A(_13942_),
    .B(_13943_),
    .C(_13944_),
    .Y(_13945_));
 sky130_fd_sc_hd__o21ai_2 _35593_ (.A1(_13696_),
    .A2(_13706_),
    .B1(_13698_),
    .Y(_13946_));
 sky130_fd_sc_hd__o21bai_2 _35594_ (.A1(_13941_),
    .A2(_13945_),
    .B1_N(_13946_),
    .Y(_13947_));
 sky130_fd_sc_hd__nand2_2 _35595_ (.A(_13933_),
    .B(_13937_),
    .Y(_13948_));
 sky130_fd_sc_hd__nand2_2 _35596_ (.A(_13948_),
    .B(_13942_),
    .Y(_13949_));
 sky130_fd_sc_hd__nand3_2 _35597_ (.A(_13933_),
    .B(_13940_),
    .C(_13938_),
    .Y(_13950_));
 sky130_fd_sc_hd__nand3_2 _35598_ (.A(_13949_),
    .B(_13950_),
    .C(_13946_),
    .Y(_13951_));
 sky130_fd_sc_hd__buf_1 _35599_ (.A(_13468_),
    .X(_13952_));
 sky130_fd_sc_hd__a21oi_2 _35600_ (.A1(_13443_),
    .A2(_13438_),
    .B1(_13952_),
    .Y(_13953_));
 sky130_fd_sc_hd__a21oi_2 _35601_ (.A1(_13947_),
    .A2(_13951_),
    .B1(_13953_),
    .Y(_13954_));
 sky130_vsdinv _35602_ (.A(_13953_),
    .Y(_13955_));
 sky130_fd_sc_hd__a21oi_2 _35603_ (.A1(_13949_),
    .A2(_13950_),
    .B1(_13946_),
    .Y(_13956_));
 sky130_vsdinv _35604_ (.A(_13951_),
    .Y(_13957_));
 sky130_fd_sc_hd__nor3_2 _35605_ (.A(_13955_),
    .B(_13956_),
    .C(_13957_),
    .Y(_13958_));
 sky130_vsdinv _35606_ (.A(_13710_),
    .Y(_13959_));
 sky130_fd_sc_hd__o21ai_2 _35607_ (.A1(_13959_),
    .A2(_13703_),
    .B1(_13713_),
    .Y(_13960_));
 sky130_fd_sc_hd__o21bai_2 _35608_ (.A1(_13954_),
    .A2(_13958_),
    .B1_N(_13960_),
    .Y(_13961_));
 sky130_fd_sc_hd__o21bai_2 _35609_ (.A1(_13956_),
    .A2(_13957_),
    .B1_N(_13953_),
    .Y(_13962_));
 sky130_fd_sc_hd__nand3_2 _35610_ (.A(_13947_),
    .B(_13953_),
    .C(_13951_),
    .Y(_13963_));
 sky130_fd_sc_hd__nand3_2 _35611_ (.A(_13962_),
    .B(_13960_),
    .C(_13963_),
    .Y(_13964_));
 sky130_fd_sc_hd__nand2_2 _35612_ (.A(_13961_),
    .B(_13964_),
    .Y(_13965_));
 sky130_fd_sc_hd__a21oi_2 _35613_ (.A1(_13712_),
    .A2(_13713_),
    .B1(_13710_),
    .Y(_13966_));
 sky130_fd_sc_hd__nor3_2 _35614_ (.A(_13959_),
    .B(_13703_),
    .C(_13709_),
    .Y(_13967_));
 sky130_fd_sc_hd__o21bai_2 _35615_ (.A1(_13966_),
    .A2(_13967_),
    .B1_N(_13717_),
    .Y(_13968_));
 sky130_fd_sc_hd__a21oi_2 _35616_ (.A1(_13725_),
    .A2(_13968_),
    .B1(_13720_),
    .Y(_13969_));
 sky130_fd_sc_hd__xor2_2 _35617_ (.A(_13965_),
    .B(_13969_),
    .X(_02662_));
 sky130_fd_sc_hd__nand2_2 _35618_ (.A(_18694_),
    .B(_07099_),
    .Y(_13970_));
 sky130_fd_sc_hd__nand3b_2 _35619_ (.A_N(_13970_),
    .B(_11599_),
    .C(_19243_),
    .Y(_13971_));
 sky130_fd_sc_hd__o21ai_2 _35620_ (.A1(_06365_),
    .A2(_16969_),
    .B1(_13970_),
    .Y(_13972_));
 sky130_fd_sc_hd__and2_2 _35621_ (.A(_11326_),
    .B(_08186_),
    .X(_13973_));
 sky130_fd_sc_hd__a21o_2 _35622_ (.A1(_13971_),
    .A2(_13972_),
    .B1(_13973_),
    .X(_13974_));
 sky130_fd_sc_hd__nand3_2 _35623_ (.A(_13971_),
    .B(_13973_),
    .C(_13972_),
    .Y(_13975_));
 sky130_fd_sc_hd__nand2_2 _35624_ (.A(_13731_),
    .B(_13727_),
    .Y(_13976_));
 sky130_fd_sc_hd__a21o_2 _35625_ (.A1(_13974_),
    .A2(_13975_),
    .B1(_13976_),
    .X(_13977_));
 sky130_fd_sc_hd__nand3_2 _35626_ (.A(_13976_),
    .B(_13974_),
    .C(_13975_),
    .Y(_13978_));
 sky130_fd_sc_hd__and2_2 _35627_ (.A(_18723_),
    .B(_07321_),
    .X(_13979_));
 sky130_fd_sc_hd__buf_1 _35628_ (.A(_13979_),
    .X(_13980_));
 sky130_fd_sc_hd__nand2_2 _35629_ (.A(_11011_),
    .B(_19225_),
    .Y(_13981_));
 sky130_fd_sc_hd__nand2_2 _35630_ (.A(_11015_),
    .B(_07328_),
    .Y(_13982_));
 sky130_fd_sc_hd__xnor2_2 _35631_ (.A(_13981_),
    .B(_13982_),
    .Y(_13983_));
 sky130_fd_sc_hd__xnor2_2 _35632_ (.A(_13980_),
    .B(_13983_),
    .Y(_13984_));
 sky130_fd_sc_hd__a21oi_2 _35633_ (.A1(_13977_),
    .A2(_13978_),
    .B1(_13984_),
    .Y(_13985_));
 sky130_fd_sc_hd__nand3_2 _35634_ (.A(_13977_),
    .B(_13984_),
    .C(_13978_),
    .Y(_13986_));
 sky130_vsdinv _35635_ (.A(_13986_),
    .Y(_13987_));
 sky130_fd_sc_hd__a21oi_2 _35636_ (.A1(_13730_),
    .A2(_13731_),
    .B1(_13732_),
    .Y(_13988_));
 sky130_fd_sc_hd__xor2_2 _35637_ (.A(_13736_),
    .B(_13739_),
    .X(_13989_));
 sky130_fd_sc_hd__o21ai_2 _35638_ (.A1(_13988_),
    .A2(_13989_),
    .B1(_13734_),
    .Y(_13990_));
 sky130_fd_sc_hd__o21bai_2 _35639_ (.A1(_13985_),
    .A2(_13987_),
    .B1_N(_13990_),
    .Y(_13991_));
 sky130_fd_sc_hd__a21o_2 _35640_ (.A1(_13977_),
    .A2(_13978_),
    .B1(_13984_),
    .X(_13992_));
 sky130_fd_sc_hd__nand3_2 _35641_ (.A(_13992_),
    .B(_13986_),
    .C(_13990_),
    .Y(_13993_));
 sky130_fd_sc_hd__nand2_2 _35642_ (.A(_10229_),
    .B(_19207_),
    .Y(_13994_));
 sky130_fd_sc_hd__nand2_2 _35643_ (.A(_18734_),
    .B(_19203_),
    .Y(_13995_));
 sky130_fd_sc_hd__xor2_2 _35644_ (.A(_13994_),
    .B(_13995_),
    .X(_13996_));
 sky130_fd_sc_hd__buf_1 _35645_ (.A(_10162_),
    .X(_13997_));
 sky130_fd_sc_hd__nand3_2 _35646_ (.A(_13996_),
    .B(_13026_),
    .C(_13997_),
    .Y(_13998_));
 sky130_fd_sc_hd__xnor2_2 _35647_ (.A(_13994_),
    .B(_13995_),
    .Y(_13999_));
 sky130_fd_sc_hd__o21ai_2 _35648_ (.A1(_12219_),
    .A2(_12845_),
    .B1(_13999_),
    .Y(_14000_));
 sky130_fd_sc_hd__nand2_2 _35649_ (.A(_13737_),
    .B(_13738_),
    .Y(_14001_));
 sky130_fd_sc_hd__nor2_2 _35650_ (.A(_13737_),
    .B(_13738_),
    .Y(_14002_));
 sky130_fd_sc_hd__a21oi_2 _35651_ (.A1(_14001_),
    .A2(_13736_),
    .B1(_14002_),
    .Y(_14003_));
 sky130_vsdinv _35652_ (.A(_14003_),
    .Y(_14004_));
 sky130_fd_sc_hd__a21oi_2 _35653_ (.A1(_13998_),
    .A2(_14000_),
    .B1(_14004_),
    .Y(_14005_));
 sky130_fd_sc_hd__o21a_2 _35654_ (.A1(_13748_),
    .A2(_13749_),
    .B1(_13751_),
    .X(_14006_));
 sky130_vsdinv _35655_ (.A(_14006_),
    .Y(_14007_));
 sky130_fd_sc_hd__nand3_2 _35656_ (.A(_13998_),
    .B(_14000_),
    .C(_14004_),
    .Y(_14008_));
 sky130_fd_sc_hd__nand3b_2 _35657_ (.A_N(_14005_),
    .B(_14007_),
    .C(_14008_),
    .Y(_14009_));
 sky130_vsdinv _35658_ (.A(_14008_),
    .Y(_14010_));
 sky130_fd_sc_hd__o21ai_2 _35659_ (.A1(_14005_),
    .A2(_14010_),
    .B1(_14006_),
    .Y(_14011_));
 sky130_fd_sc_hd__nand2_2 _35660_ (.A(_14009_),
    .B(_14011_),
    .Y(_14012_));
 sky130_fd_sc_hd__buf_1 _35661_ (.A(_14012_),
    .X(_14013_));
 sky130_fd_sc_hd__a21boi_2 _35662_ (.A1(_13991_),
    .A2(_13993_),
    .B1_N(_14013_),
    .Y(_14014_));
 sky130_fd_sc_hd__a21oi_2 _35663_ (.A1(_13992_),
    .A2(_13986_),
    .B1(_13990_),
    .Y(_14015_));
 sky130_vsdinv _35664_ (.A(_13993_),
    .Y(_14016_));
 sky130_fd_sc_hd__nor3_2 _35665_ (.A(_14013_),
    .B(_14015_),
    .C(_14016_),
    .Y(_14017_));
 sky130_fd_sc_hd__o21ai_2 _35666_ (.A1(_13768_),
    .A2(_13770_),
    .B1(_13747_),
    .Y(_14018_));
 sky130_fd_sc_hd__o21bai_2 _35667_ (.A1(_14014_),
    .A2(_14017_),
    .B1_N(_14018_),
    .Y(_14019_));
 sky130_fd_sc_hd__o21ai_2 _35668_ (.A1(_14015_),
    .A2(_14016_),
    .B1(_14013_),
    .Y(_14020_));
 sky130_fd_sc_hd__nand3b_2 _35669_ (.A_N(_14012_),
    .B(_13991_),
    .C(_13993_),
    .Y(_14021_));
 sky130_fd_sc_hd__nand3_2 _35670_ (.A(_14020_),
    .B(_14021_),
    .C(_14018_),
    .Y(_14022_));
 sky130_fd_sc_hd__nand2_2 _35671_ (.A(_10421_),
    .B(_12004_),
    .Y(_14023_));
 sky130_fd_sc_hd__nand2_2 _35672_ (.A(_12794_),
    .B(_10070_),
    .Y(_14024_));
 sky130_fd_sc_hd__nand2_2 _35673_ (.A(_14023_),
    .B(_14024_),
    .Y(_14025_));
 sky130_fd_sc_hd__nand3b_2 _35674_ (.A_N(_14023_),
    .B(_10734_),
    .C(_09104_),
    .Y(_14026_));
 sky130_fd_sc_hd__o2bb2ai_2 _35675_ (.A1_N(_14025_),
    .A2_N(_14026_),
    .B1(_18760_),
    .B2(_09092_),
    .Y(_14027_));
 sky130_fd_sc_hd__and2_2 _35676_ (.A(_12531_),
    .B(_12836_),
    .X(_14028_));
 sky130_fd_sc_hd__nand3_2 _35677_ (.A(_14026_),
    .B(_14025_),
    .C(_14028_),
    .Y(_14029_));
 sky130_fd_sc_hd__a21oi_2 _35678_ (.A1(_13784_),
    .A2(_13782_),
    .B1(_13781_),
    .Y(_14030_));
 sky130_vsdinv _35679_ (.A(_14030_),
    .Y(_14031_));
 sky130_fd_sc_hd__a21o_2 _35680_ (.A1(_14027_),
    .A2(_14029_),
    .B1(_14031_),
    .X(_14032_));
 sky130_fd_sc_hd__nand3_2 _35681_ (.A(_14027_),
    .B(_14031_),
    .C(_14029_),
    .Y(_14033_));
 sky130_fd_sc_hd__and2_2 _35682_ (.A(_12538_),
    .B(_10849_),
    .X(_14034_));
 sky130_fd_sc_hd__nand2_2 _35683_ (.A(_18771_),
    .B(_09790_),
    .Y(_14035_));
 sky130_fd_sc_hd__nand3b_2 _35684_ (.A_N(_14035_),
    .B(_08219_),
    .C(_09785_),
    .Y(_14036_));
 sky130_fd_sc_hd__a22o_2 _35685_ (.A1(_12540_),
    .A2(_12842_),
    .B1(_10433_),
    .B2(_11224_),
    .X(_14037_));
 sky130_fd_sc_hd__nand2_2 _35686_ (.A(_14036_),
    .B(_14037_),
    .Y(_14038_));
 sky130_fd_sc_hd__xnor2_2 _35687_ (.A(_14034_),
    .B(_14038_),
    .Y(_14039_));
 sky130_fd_sc_hd__a21o_2 _35688_ (.A1(_14032_),
    .A2(_14033_),
    .B1(_14039_),
    .X(_14040_));
 sky130_fd_sc_hd__nand3_2 _35689_ (.A(_14032_),
    .B(_14039_),
    .C(_14033_),
    .Y(_14041_));
 sky130_fd_sc_hd__o21ai_2 _35690_ (.A1(_13762_),
    .A2(_13758_),
    .B1(_13759_),
    .Y(_14042_));
 sky130_fd_sc_hd__a21o_2 _35691_ (.A1(_14040_),
    .A2(_14041_),
    .B1(_14042_),
    .X(_14043_));
 sky130_fd_sc_hd__nand3_2 _35692_ (.A(_14040_),
    .B(_14042_),
    .C(_14041_),
    .Y(_14044_));
 sky130_fd_sc_hd__a21boi_2 _35693_ (.A1(_13792_),
    .A2(_13798_),
    .B1_N(_13793_),
    .Y(_14045_));
 sky130_vsdinv _35694_ (.A(_14045_),
    .Y(_14046_));
 sky130_fd_sc_hd__a21o_2 _35695_ (.A1(_14043_),
    .A2(_14044_),
    .B1(_14046_),
    .X(_14047_));
 sky130_fd_sc_hd__nand3_2 _35696_ (.A(_14043_),
    .B(_14046_),
    .C(_14044_),
    .Y(_14048_));
 sky130_fd_sc_hd__nand2_2 _35697_ (.A(_14047_),
    .B(_14048_),
    .Y(_14049_));
 sky130_fd_sc_hd__buf_1 _35698_ (.A(_14049_),
    .X(_14050_));
 sky130_fd_sc_hd__a21boi_2 _35699_ (.A1(_14019_),
    .A2(_14022_),
    .B1_N(_14050_),
    .Y(_14051_));
 sky130_fd_sc_hd__a21oi_2 _35700_ (.A1(_14020_),
    .A2(_14021_),
    .B1(_14018_),
    .Y(_14052_));
 sky130_vsdinv _35701_ (.A(_14022_),
    .Y(_14053_));
 sky130_fd_sc_hd__nor3_2 _35702_ (.A(_14050_),
    .B(_14052_),
    .C(_14053_),
    .Y(_14054_));
 sky130_fd_sc_hd__o21ai_2 _35703_ (.A1(_13816_),
    .A2(_13817_),
    .B1(_13778_),
    .Y(_14055_));
 sky130_fd_sc_hd__o21bai_2 _35704_ (.A1(_14051_),
    .A2(_14054_),
    .B1_N(_14055_),
    .Y(_14056_));
 sky130_fd_sc_hd__o21ai_2 _35705_ (.A1(_14052_),
    .A2(_14053_),
    .B1(_14050_),
    .Y(_14057_));
 sky130_fd_sc_hd__nand3b_2 _35706_ (.A_N(_14049_),
    .B(_14019_),
    .C(_14022_),
    .Y(_14058_));
 sky130_fd_sc_hd__nand3_2 _35707_ (.A(_14057_),
    .B(_14058_),
    .C(_14055_),
    .Y(_14059_));
 sky130_fd_sc_hd__nand2_2 _35708_ (.A(_10120_),
    .B(_10535_),
    .Y(_14060_));
 sky130_fd_sc_hd__nand2_2 _35709_ (.A(_08391_),
    .B(_10551_),
    .Y(_14061_));
 sky130_fd_sc_hd__xor2_2 _35710_ (.A(_14060_),
    .B(_14061_),
    .X(_14062_));
 sky130_fd_sc_hd__nand3_2 _35711_ (.A(_14062_),
    .B(_13089_),
    .C(_10895_),
    .Y(_14063_));
 sky130_fd_sc_hd__xnor2_2 _35712_ (.A(_14060_),
    .B(_14061_),
    .Y(_14064_));
 sky130_fd_sc_hd__o21ai_2 _35713_ (.A1(_10780_),
    .A2(_19145_),
    .B1(_14064_),
    .Y(_14065_));
 sky130_fd_sc_hd__nand2_2 _35714_ (.A(_13795_),
    .B(_13796_),
    .Y(_14066_));
 sky130_fd_sc_hd__nor2_2 _35715_ (.A(_13795_),
    .B(_13796_),
    .Y(_14067_));
 sky130_fd_sc_hd__a21oi_2 _35716_ (.A1(_14066_),
    .A2(_13794_),
    .B1(_14067_),
    .Y(_14068_));
 sky130_vsdinv _35717_ (.A(_14068_),
    .Y(_14069_));
 sky130_fd_sc_hd__a21oi_2 _35718_ (.A1(_14063_),
    .A2(_14065_),
    .B1(_14069_),
    .Y(_14070_));
 sky130_fd_sc_hd__nand3_2 _35719_ (.A(_14063_),
    .B(_14065_),
    .C(_14069_),
    .Y(_14071_));
 sky130_vsdinv _35720_ (.A(_14071_),
    .Y(_14072_));
 sky130_fd_sc_hd__o21a_2 _35721_ (.A1(_13827_),
    .A2(_13828_),
    .B1(_13832_),
    .X(_14073_));
 sky130_fd_sc_hd__o21ai_2 _35722_ (.A1(_14070_),
    .A2(_14072_),
    .B1(_14073_),
    .Y(_14074_));
 sky130_fd_sc_hd__a21o_2 _35723_ (.A1(_14063_),
    .A2(_14065_),
    .B1(_14069_),
    .X(_14075_));
 sky130_fd_sc_hd__nand3b_2 _35724_ (.A_N(_14073_),
    .B(_14075_),
    .C(_14071_),
    .Y(_14076_));
 sky130_fd_sc_hd__a21boi_2 _35725_ (.A1(_13832_),
    .A2(_13834_),
    .B1_N(_13836_),
    .Y(_14077_));
 sky130_fd_sc_hd__o21ai_2 _35726_ (.A1(_13840_),
    .A2(_14077_),
    .B1(_13838_),
    .Y(_14078_));
 sky130_fd_sc_hd__a21o_2 _35727_ (.A1(_14074_),
    .A2(_14076_),
    .B1(_14078_),
    .X(_14079_));
 sky130_fd_sc_hd__nand3_2 _35728_ (.A(_14074_),
    .B(_14078_),
    .C(_14076_),
    .Y(_14080_));
 sky130_fd_sc_hd__nand2_2 _35729_ (.A(_08169_),
    .B(_10912_),
    .Y(_14081_));
 sky130_fd_sc_hd__nand2_2 _35730_ (.A(_09870_),
    .B(_19132_),
    .Y(_14082_));
 sky130_fd_sc_hd__xor2_2 _35731_ (.A(_14081_),
    .B(_14082_),
    .X(_14083_));
 sky130_fd_sc_hd__and2_2 _35732_ (.A(_16961_),
    .B(_07195_),
    .X(_14084_));
 sky130_fd_sc_hd__buf_1 _35733_ (.A(_14084_),
    .X(_14085_));
 sky130_fd_sc_hd__nand2_2 _35734_ (.A(_14083_),
    .B(_14085_),
    .Y(_14086_));
 sky130_fd_sc_hd__xnor2_2 _35735_ (.A(_14081_),
    .B(_14082_),
    .Y(_14087_));
 sky130_vsdinv _35736_ (.A(_14084_),
    .Y(_14088_));
 sky130_fd_sc_hd__nand2_2 _35737_ (.A(_14087_),
    .B(_14088_),
    .Y(_14089_));
 sky130_fd_sc_hd__nand2_2 _35738_ (.A(_14086_),
    .B(_14089_),
    .Y(_14090_));
 sky130_fd_sc_hd__o211ai_2 _35739_ (.A1(_13847_),
    .A2(_13848_),
    .B1(_13853_),
    .C1(_14090_),
    .Y(_14091_));
 sky130_fd_sc_hd__o21ai_2 _35740_ (.A1(_13847_),
    .A2(_13848_),
    .B1(_13853_),
    .Y(_14092_));
 sky130_fd_sc_hd__nand3_2 _35741_ (.A(_14092_),
    .B(_14089_),
    .C(_14086_),
    .Y(_14093_));
 sky130_fd_sc_hd__o2bb2ai_2 _35742_ (.A1_N(_14091_),
    .A2_N(_14093_),
    .B1(_13860_),
    .B2(_13861_),
    .Y(_14094_));
 sky130_fd_sc_hd__nand3_2 _35743_ (.A(_14091_),
    .B(_14093_),
    .C(_13864_),
    .Y(_14095_));
 sky130_fd_sc_hd__nand2_2 _35744_ (.A(_14094_),
    .B(_14095_),
    .Y(_14096_));
 sky130_vsdinv _35745_ (.A(_14096_),
    .Y(_14097_));
 sky130_fd_sc_hd__a21oi_2 _35746_ (.A1(_14079_),
    .A2(_14080_),
    .B1(_14097_),
    .Y(_14098_));
 sky130_fd_sc_hd__nand3_2 _35747_ (.A(_14097_),
    .B(_14079_),
    .C(_14080_),
    .Y(_14099_));
 sky130_vsdinv _35748_ (.A(_14099_),
    .Y(_14100_));
 sky130_fd_sc_hd__a21oi_2 _35749_ (.A1(_13804_),
    .A2(_13800_),
    .B1(_13802_),
    .Y(_14101_));
 sky130_fd_sc_hd__o21ai_2 _35750_ (.A1(_13807_),
    .A2(_14101_),
    .B1(_13805_),
    .Y(_14102_));
 sky130_fd_sc_hd__o21bai_2 _35751_ (.A1(_14098_),
    .A2(_14100_),
    .B1_N(_14102_),
    .Y(_14103_));
 sky130_fd_sc_hd__nand3b_2 _35752_ (.A_N(_14098_),
    .B(_14102_),
    .C(_14099_),
    .Y(_14104_));
 sky130_fd_sc_hd__nand2_2 _35753_ (.A(_14103_),
    .B(_14104_),
    .Y(_14105_));
 sky130_vsdinv _35754_ (.A(_13845_),
    .Y(_14106_));
 sky130_fd_sc_hd__a21oi_2 _35755_ (.A1(_13844_),
    .A2(_13866_),
    .B1(_14106_),
    .Y(_14107_));
 sky130_fd_sc_hd__nand2_2 _35756_ (.A(_14105_),
    .B(_14107_),
    .Y(_14108_));
 sky130_vsdinv _35757_ (.A(_14107_),
    .Y(_14109_));
 sky130_fd_sc_hd__nand3_2 _35758_ (.A(_14103_),
    .B(_14109_),
    .C(_14104_),
    .Y(_14110_));
 sky130_fd_sc_hd__nand2_2 _35759_ (.A(_14108_),
    .B(_14110_),
    .Y(_14111_));
 sky130_fd_sc_hd__buf_1 _35760_ (.A(_14111_),
    .X(_14112_));
 sky130_fd_sc_hd__a21boi_2 _35761_ (.A1(_14056_),
    .A2(_14059_),
    .B1_N(_14112_),
    .Y(_14113_));
 sky130_fd_sc_hd__nand2_2 _35762_ (.A(_14056_),
    .B(_14059_),
    .Y(_14114_));
 sky130_fd_sc_hd__nor2_2 _35763_ (.A(_14112_),
    .B(_14114_),
    .Y(_14115_));
 sky130_fd_sc_hd__o21ai_2 _35764_ (.A1(_13880_),
    .A2(_13882_),
    .B1(_13826_),
    .Y(_14116_));
 sky130_fd_sc_hd__o21bai_2 _35765_ (.A1(_14113_),
    .A2(_14115_),
    .B1_N(_14116_),
    .Y(_14117_));
 sky130_fd_sc_hd__nand2_2 _35766_ (.A(_14114_),
    .B(_14112_),
    .Y(_14118_));
 sky130_fd_sc_hd__nand3b_2 _35767_ (.A_N(_14111_),
    .B(_14056_),
    .C(_14059_),
    .Y(_14119_));
 sky130_fd_sc_hd__nand3_2 _35768_ (.A(_14118_),
    .B(_14119_),
    .C(_14116_),
    .Y(_14120_));
 sky130_fd_sc_hd__nand2_2 _35769_ (.A(_13865_),
    .B(_13854_),
    .Y(_14121_));
 sky130_fd_sc_hd__o21bai_2 _35770_ (.A1(_13857_),
    .A2(_13364_),
    .B1_N(_13859_),
    .Y(_14122_));
 sky130_fd_sc_hd__o21bai_2 _35771_ (.A1(_13156_),
    .A2(_13158_),
    .B1_N(_14122_),
    .Y(_14123_));
 sky130_fd_sc_hd__nand3b_2 _35772_ (.A_N(_13155_),
    .B(_13159_),
    .C(_14122_),
    .Y(_14124_));
 sky130_fd_sc_hd__a21oi_2 _35773_ (.A1(_14123_),
    .A2(_14124_),
    .B1(_13418_),
    .Y(_14125_));
 sky130_fd_sc_hd__o211a_2 _35774_ (.A1(_13408_),
    .A2(_13163_),
    .B1(_14124_),
    .C1(_14123_),
    .X(_14126_));
 sky130_fd_sc_hd__nor2_2 _35775_ (.A(_14125_),
    .B(_14126_),
    .Y(_14127_));
 sky130_fd_sc_hd__buf_1 _35776_ (.A(_14127_),
    .X(_14128_));
 sky130_fd_sc_hd__nand2_2 _35777_ (.A(_14121_),
    .B(_14128_),
    .Y(_14129_));
 sky130_fd_sc_hd__o211ai_2 _35778_ (.A1(_14125_),
    .A2(_14126_),
    .B1(_13854_),
    .C1(_13865_),
    .Y(_14130_));
 sky130_fd_sc_hd__a21oi_2 _35779_ (.A1(_13896_),
    .A2(_13650_),
    .B1(_13894_),
    .Y(_14131_));
 sky130_vsdinv _35780_ (.A(_14131_),
    .Y(_14132_));
 sky130_fd_sc_hd__a21oi_2 _35781_ (.A1(_14129_),
    .A2(_14130_),
    .B1(_14132_),
    .Y(_14133_));
 sky130_fd_sc_hd__nand3_2 _35782_ (.A(_14129_),
    .B(_14130_),
    .C(_14132_),
    .Y(_14134_));
 sky130_vsdinv _35783_ (.A(_14134_),
    .Y(_14135_));
 sky130_fd_sc_hd__o211ai_2 _35784_ (.A1(_14133_),
    .A2(_14135_),
    .B1(_13901_),
    .C1(_13906_),
    .Y(_14136_));
 sky130_fd_sc_hd__nand2_2 _35785_ (.A(_13906_),
    .B(_13901_),
    .Y(_14137_));
 sky130_fd_sc_hd__nand3b_2 _35786_ (.A_N(_14133_),
    .B(_14137_),
    .C(_14134_),
    .Y(_14138_));
 sky130_fd_sc_hd__a21oi_2 _35787_ (.A1(_14136_),
    .A2(_14138_),
    .B1(_13432_),
    .Y(_14139_));
 sky130_fd_sc_hd__nand3_2 _35788_ (.A(_14136_),
    .B(_14138_),
    .C(_13183_),
    .Y(_14140_));
 sky130_vsdinv _35789_ (.A(_14140_),
    .Y(_14141_));
 sky130_fd_sc_hd__a21boi_2 _35790_ (.A1(_13871_),
    .A2(_13877_),
    .B1_N(_13873_),
    .Y(_14142_));
 sky130_fd_sc_hd__o21ai_2 _35791_ (.A1(_14139_),
    .A2(_14141_),
    .B1(_14142_),
    .Y(_14143_));
 sky130_fd_sc_hd__nand2_2 _35792_ (.A(_13878_),
    .B(_13873_),
    .Y(_14144_));
 sky130_fd_sc_hd__nand3b_2 _35793_ (.A_N(_14139_),
    .B(_14144_),
    .C(_14140_),
    .Y(_14145_));
 sky130_fd_sc_hd__buf_1 _35794_ (.A(_14145_),
    .X(_14146_));
 sky130_fd_sc_hd__a21boi_2 _35795_ (.A1(_13909_),
    .A2(_13193_),
    .B1_N(_13910_),
    .Y(_14147_));
 sky130_vsdinv _35796_ (.A(_14147_),
    .Y(_14148_));
 sky130_fd_sc_hd__a21oi_2 _35797_ (.A1(_14143_),
    .A2(_14146_),
    .B1(_14148_),
    .Y(_14149_));
 sky130_fd_sc_hd__nand3_2 _35798_ (.A(_14143_),
    .B(_14145_),
    .C(_14148_),
    .Y(_14150_));
 sky130_vsdinv _35799_ (.A(_14150_),
    .Y(_14151_));
 sky130_fd_sc_hd__nor2_2 _35800_ (.A(_14149_),
    .B(_14151_),
    .Y(_14152_));
 sky130_fd_sc_hd__a21oi_2 _35801_ (.A1(_14117_),
    .A2(_14120_),
    .B1(_14152_),
    .Y(_14153_));
 sky130_fd_sc_hd__a21o_2 _35802_ (.A1(_14143_),
    .A2(_14146_),
    .B1(_14148_),
    .X(_14154_));
 sky130_fd_sc_hd__nand2_2 _35803_ (.A(_14154_),
    .B(_14150_),
    .Y(_14155_));
 sky130_fd_sc_hd__a21oi_2 _35804_ (.A1(_14118_),
    .A2(_14119_),
    .B1(_14116_),
    .Y(_14156_));
 sky130_vsdinv _35805_ (.A(_14120_),
    .Y(_14157_));
 sky130_fd_sc_hd__nor3_2 _35806_ (.A(_14155_),
    .B(_14156_),
    .C(_14157_),
    .Y(_14158_));
 sky130_fd_sc_hd__o21ai_2 _35807_ (.A1(_13928_),
    .A2(_13929_),
    .B1(_13890_),
    .Y(_14159_));
 sky130_fd_sc_hd__o21bai_2 _35808_ (.A1(_14153_),
    .A2(_14158_),
    .B1_N(_14159_),
    .Y(_14160_));
 sky130_fd_sc_hd__o22ai_2 _35809_ (.A1(_14151_),
    .A2(_14149_),
    .B1(_14156_),
    .B2(_14157_),
    .Y(_14161_));
 sky130_fd_sc_hd__nand3_2 _35810_ (.A(_14152_),
    .B(_14117_),
    .C(_14120_),
    .Y(_14162_));
 sky130_fd_sc_hd__nand3_2 _35811_ (.A(_14161_),
    .B(_14162_),
    .C(_14159_),
    .Y(_14163_));
 sky130_fd_sc_hd__nand2_2 _35812_ (.A(_14160_),
    .B(_14163_),
    .Y(_14164_));
 sky130_fd_sc_hd__nand2_2 _35813_ (.A(_13922_),
    .B(_13918_),
    .Y(_14165_));
 sky130_fd_sc_hd__xor2_2 _35814_ (.A(_13213_),
    .B(_14165_),
    .X(_14166_));
 sky130_vsdinv _35815_ (.A(_14166_),
    .Y(_14167_));
 sky130_fd_sc_hd__nand2_2 _35816_ (.A(_14164_),
    .B(_14167_),
    .Y(_14168_));
 sky130_fd_sc_hd__buf_1 _35817_ (.A(_14163_),
    .X(_14169_));
 sky130_fd_sc_hd__nand3_2 _35818_ (.A(_14160_),
    .B(_14166_),
    .C(_14169_),
    .Y(_14170_));
 sky130_fd_sc_hd__o21ai_2 _35819_ (.A1(_13942_),
    .A2(_13943_),
    .B1(_13938_),
    .Y(_14171_));
 sky130_fd_sc_hd__a21oi_2 _35820_ (.A1(_14168_),
    .A2(_14170_),
    .B1(_14171_),
    .Y(_14172_));
 sky130_fd_sc_hd__nand3_2 _35821_ (.A(_14168_),
    .B(_14170_),
    .C(_14171_),
    .Y(_14173_));
 sky130_vsdinv _35822_ (.A(_14173_),
    .Y(_14174_));
 sky130_fd_sc_hd__a21oi_2 _35823_ (.A1(_13676_),
    .A2(_13671_),
    .B1(_13952_),
    .Y(_14175_));
 sky130_fd_sc_hd__o21bai_2 _35824_ (.A1(_14172_),
    .A2(_14174_),
    .B1_N(_14175_),
    .Y(_14176_));
 sky130_fd_sc_hd__a21oi_2 _35825_ (.A1(_14160_),
    .A2(_14169_),
    .B1(_14166_),
    .Y(_14177_));
 sky130_fd_sc_hd__a21oi_2 _35826_ (.A1(_14161_),
    .A2(_14162_),
    .B1(_14159_),
    .Y(_14178_));
 sky130_fd_sc_hd__nor3b_2 _35827_ (.A(_14167_),
    .B(_14178_),
    .C_N(_14169_),
    .Y(_14179_));
 sky130_fd_sc_hd__o21bai_2 _35828_ (.A1(_14177_),
    .A2(_14179_),
    .B1_N(_14171_),
    .Y(_14180_));
 sky130_fd_sc_hd__nand3_2 _35829_ (.A(_14180_),
    .B(_14175_),
    .C(_14173_),
    .Y(_14181_));
 sky130_fd_sc_hd__o21ai_2 _35830_ (.A1(_13955_),
    .A2(_13956_),
    .B1(_13951_),
    .Y(_14182_));
 sky130_fd_sc_hd__a21oi_2 _35831_ (.A1(_14176_),
    .A2(_14181_),
    .B1(_14182_),
    .Y(_14183_));
 sky130_fd_sc_hd__nand3_2 _35832_ (.A(_14176_),
    .B(_14181_),
    .C(_14182_),
    .Y(_14184_));
 sky130_vsdinv _35833_ (.A(_14184_),
    .Y(_14185_));
 sky130_fd_sc_hd__nor2_2 _35834_ (.A(_14183_),
    .B(_14185_),
    .Y(_14186_));
 sky130_fd_sc_hd__nor2_2 _35835_ (.A(_13238_),
    .B(_13477_),
    .Y(_14187_));
 sky130_fd_sc_hd__nand2_2 _35836_ (.A(_13968_),
    .B(_13719_),
    .Y(_14188_));
 sky130_fd_sc_hd__nor2_2 _35837_ (.A(_14188_),
    .B(_13965_),
    .Y(_14189_));
 sky130_fd_sc_hd__nand2_2 _35838_ (.A(_14187_),
    .B(_14189_),
    .Y(_14190_));
 sky130_fd_sc_hd__nand3b_2 _35839_ (.A_N(_13965_),
    .B(_13723_),
    .C(_13721_),
    .Y(_14191_));
 sky130_fd_sc_hd__a21boi_2 _35840_ (.A1(_13720_),
    .A2(_13961_),
    .B1_N(_13964_),
    .Y(_14192_));
 sky130_fd_sc_hd__nand2_2 _35841_ (.A(_14191_),
    .B(_14192_),
    .Y(_14193_));
 sky130_fd_sc_hd__o21bai_2 _35842_ (.A1(_14190_),
    .A2(_13247_),
    .B1_N(_14193_),
    .Y(_14194_));
 sky130_fd_sc_hd__xor2_2 _35843_ (.A(_14186_),
    .B(_14194_),
    .X(_02663_));
 sky130_fd_sc_hd__nand2_2 _35844_ (.A(_10669_),
    .B(_07698_),
    .Y(_14195_));
 sky130_fd_sc_hd__nand3b_2 _35845_ (.A_N(_14195_),
    .B(_11322_),
    .C(_19238_),
    .Y(_14196_));
 sky130_fd_sc_hd__o21ai_2 _35846_ (.A1(_06616_),
    .A2(_11005_),
    .B1(_14195_),
    .Y(_14197_));
 sky130_fd_sc_hd__and2_2 _35847_ (.A(_10267_),
    .B(_06745_),
    .X(_14198_));
 sky130_fd_sc_hd__a21o_2 _35848_ (.A1(_14196_),
    .A2(_14197_),
    .B1(_14198_),
    .X(_14199_));
 sky130_fd_sc_hd__nand3_2 _35849_ (.A(_14196_),
    .B(_14198_),
    .C(_14197_),
    .Y(_14200_));
 sky130_fd_sc_hd__nand2_2 _35850_ (.A(_13975_),
    .B(_13971_),
    .Y(_14201_));
 sky130_fd_sc_hd__a21o_2 _35851_ (.A1(_14199_),
    .A2(_14200_),
    .B1(_14201_),
    .X(_14202_));
 sky130_fd_sc_hd__nand3_2 _35852_ (.A(_14201_),
    .B(_14199_),
    .C(_14200_),
    .Y(_14203_));
 sky130_fd_sc_hd__and2_2 _35853_ (.A(_10474_),
    .B(_09364_),
    .X(_14204_));
 sky130_fd_sc_hd__buf_1 _35854_ (.A(_14204_),
    .X(_14205_));
 sky130_fd_sc_hd__nand2_2 _35855_ (.A(_09958_),
    .B(_19216_),
    .Y(_14206_));
 sky130_fd_sc_hd__nand2_2 _35856_ (.A(_10262_),
    .B(_08258_),
    .Y(_14207_));
 sky130_fd_sc_hd__xnor2_2 _35857_ (.A(_14206_),
    .B(_14207_),
    .Y(_14208_));
 sky130_fd_sc_hd__xnor2_2 _35858_ (.A(_14205_),
    .B(_14208_),
    .Y(_14209_));
 sky130_fd_sc_hd__a21oi_2 _35859_ (.A1(_14202_),
    .A2(_14203_),
    .B1(_14209_),
    .Y(_14210_));
 sky130_fd_sc_hd__nand3_2 _35860_ (.A(_14202_),
    .B(_14209_),
    .C(_14203_),
    .Y(_14211_));
 sky130_vsdinv _35861_ (.A(_14211_),
    .Y(_14212_));
 sky130_fd_sc_hd__a21oi_2 _35862_ (.A1(_13974_),
    .A2(_13975_),
    .B1(_13976_),
    .Y(_14213_));
 sky130_fd_sc_hd__xor2_2 _35863_ (.A(_13980_),
    .B(_13983_),
    .X(_14214_));
 sky130_fd_sc_hd__o21ai_2 _35864_ (.A1(_14213_),
    .A2(_14214_),
    .B1(_13978_),
    .Y(_14215_));
 sky130_fd_sc_hd__o21bai_2 _35865_ (.A1(_14210_),
    .A2(_14212_),
    .B1_N(_14215_),
    .Y(_14216_));
 sky130_fd_sc_hd__a21o_2 _35866_ (.A1(_14202_),
    .A2(_14203_),
    .B1(_14209_),
    .X(_14217_));
 sky130_fd_sc_hd__nand3_2 _35867_ (.A(_14217_),
    .B(_14211_),
    .C(_14215_),
    .Y(_14218_));
 sky130_fd_sc_hd__nand2_2 _35868_ (.A(_10452_),
    .B(_07310_),
    .Y(_14219_));
 sky130_fd_sc_hd__nand2_2 _35869_ (.A(_10453_),
    .B(_10159_),
    .Y(_14220_));
 sky130_fd_sc_hd__xor2_2 _35870_ (.A(_14219_),
    .B(_14220_),
    .X(_14221_));
 sky130_fd_sc_hd__nand3_2 _35871_ (.A(_14221_),
    .B(_13508_),
    .C(_13787_),
    .Y(_14222_));
 sky130_fd_sc_hd__xnor2_2 _35872_ (.A(_14219_),
    .B(_14220_),
    .Y(_14223_));
 sky130_fd_sc_hd__o21ai_2 _35873_ (.A1(_10246_),
    .A2(_19193_),
    .B1(_14223_),
    .Y(_14224_));
 sky130_fd_sc_hd__nand2_2 _35874_ (.A(_13981_),
    .B(_13982_),
    .Y(_14225_));
 sky130_fd_sc_hd__nor2_2 _35875_ (.A(_13981_),
    .B(_13982_),
    .Y(_14226_));
 sky130_fd_sc_hd__a21oi_2 _35876_ (.A1(_14225_),
    .A2(_13980_),
    .B1(_14226_),
    .Y(_14227_));
 sky130_fd_sc_hd__a21bo_2 _35877_ (.A1(_14222_),
    .A2(_14224_),
    .B1_N(_14227_),
    .X(_14228_));
 sky130_fd_sc_hd__nand3b_2 _35878_ (.A_N(_14227_),
    .B(_14222_),
    .C(_14224_),
    .Y(_14229_));
 sky130_fd_sc_hd__o21ai_2 _35879_ (.A1(_13994_),
    .A2(_13995_),
    .B1(_13998_),
    .Y(_14230_));
 sky130_fd_sc_hd__a21o_2 _35880_ (.A1(_14228_),
    .A2(_14229_),
    .B1(_14230_),
    .X(_14231_));
 sky130_fd_sc_hd__nand3_2 _35881_ (.A(_14228_),
    .B(_14230_),
    .C(_14229_),
    .Y(_14232_));
 sky130_fd_sc_hd__nand2_2 _35882_ (.A(_14231_),
    .B(_14232_),
    .Y(_14233_));
 sky130_fd_sc_hd__buf_1 _35883_ (.A(_14233_),
    .X(_14234_));
 sky130_fd_sc_hd__a21boi_2 _35884_ (.A1(_14216_),
    .A2(_14218_),
    .B1_N(_14234_),
    .Y(_14235_));
 sky130_fd_sc_hd__a21oi_2 _35885_ (.A1(_14217_),
    .A2(_14211_),
    .B1(_14215_),
    .Y(_14236_));
 sky130_vsdinv _35886_ (.A(_14218_),
    .Y(_14237_));
 sky130_fd_sc_hd__nor3_2 _35887_ (.A(_14234_),
    .B(_14236_),
    .C(_14237_),
    .Y(_14238_));
 sky130_fd_sc_hd__o21ai_2 _35888_ (.A1(_14013_),
    .A2(_14015_),
    .B1(_13993_),
    .Y(_14239_));
 sky130_fd_sc_hd__o21bai_2 _35889_ (.A1(_14235_),
    .A2(_14238_),
    .B1_N(_14239_),
    .Y(_14240_));
 sky130_fd_sc_hd__o21ai_2 _35890_ (.A1(_14236_),
    .A2(_14237_),
    .B1(_14234_),
    .Y(_14241_));
 sky130_fd_sc_hd__nand3b_2 _35891_ (.A_N(_14233_),
    .B(_14218_),
    .C(_14216_),
    .Y(_14242_));
 sky130_fd_sc_hd__nand3_2 _35892_ (.A(_14241_),
    .B(_14242_),
    .C(_14239_),
    .Y(_14243_));
 sky130_fd_sc_hd__buf_1 _35893_ (.A(_14243_),
    .X(_14244_));
 sky130_fd_sc_hd__buf_1 _35894_ (.A(_10186_),
    .X(_14245_));
 sky130_fd_sc_hd__nand2_2 _35895_ (.A(_14245_),
    .B(_07952_),
    .Y(_14246_));
 sky130_fd_sc_hd__nand2_2 _35896_ (.A(_13305_),
    .B(_12836_),
    .Y(_14247_));
 sky130_fd_sc_hd__nand2_2 _35897_ (.A(_14246_),
    .B(_14247_),
    .Y(_14248_));
 sky130_fd_sc_hd__nor2_2 _35898_ (.A(_14246_),
    .B(_14247_),
    .Y(_14249_));
 sky130_vsdinv _35899_ (.A(_14249_),
    .Y(_14250_));
 sky130_fd_sc_hd__o2bb2ai_2 _35900_ (.A1_N(_14248_),
    .A2_N(_14250_),
    .B1(_13050_),
    .B2(_19175_),
    .Y(_14251_));
 sky130_fd_sc_hd__and2_2 _35901_ (.A(_08085_),
    .B(_10576_),
    .X(_14252_));
 sky130_fd_sc_hd__nand3b_2 _35902_ (.A_N(_14249_),
    .B(_14248_),
    .C(_14252_),
    .Y(_14253_));
 sky130_fd_sc_hd__nor2_2 _35903_ (.A(_14023_),
    .B(_14024_),
    .Y(_14254_));
 sky130_fd_sc_hd__a21oi_2 _35904_ (.A1(_14025_),
    .A2(_14028_),
    .B1(_14254_),
    .Y(_14255_));
 sky130_vsdinv _35905_ (.A(_14255_),
    .Y(_14256_));
 sky130_fd_sc_hd__a21o_2 _35906_ (.A1(_14251_),
    .A2(_14253_),
    .B1(_14256_),
    .X(_14257_));
 sky130_fd_sc_hd__nand3_2 _35907_ (.A(_14251_),
    .B(_14253_),
    .C(_14256_),
    .Y(_14258_));
 sky130_fd_sc_hd__and2_2 _35908_ (.A(_12538_),
    .B(_10052_),
    .X(_14259_));
 sky130_fd_sc_hd__nand2_2 _35909_ (.A(_10433_),
    .B(_10531_),
    .Y(_14260_));
 sky130_fd_sc_hd__nand3b_2 _35910_ (.A_N(_14260_),
    .B(_18766_),
    .C(_09787_),
    .Y(_14261_));
 sky130_fd_sc_hd__a22o_2 _35911_ (.A1(_12805_),
    .A2(_12325_),
    .B1(_08220_),
    .B2(_10538_),
    .X(_14262_));
 sky130_fd_sc_hd__nand2_2 _35912_ (.A(_14261_),
    .B(_14262_),
    .Y(_14263_));
 sky130_fd_sc_hd__xnor2_2 _35913_ (.A(_14259_),
    .B(_14263_),
    .Y(_14264_));
 sky130_fd_sc_hd__a21oi_2 _35914_ (.A1(_14257_),
    .A2(_14258_),
    .B1(_14264_),
    .Y(_14265_));
 sky130_fd_sc_hd__nand3_2 _35915_ (.A(_14257_),
    .B(_14264_),
    .C(_14258_),
    .Y(_14266_));
 sky130_vsdinv _35916_ (.A(_14266_),
    .Y(_14267_));
 sky130_fd_sc_hd__o21ai_2 _35917_ (.A1(_14006_),
    .A2(_14005_),
    .B1(_14008_),
    .Y(_14268_));
 sky130_fd_sc_hd__o21bai_2 _35918_ (.A1(_14265_),
    .A2(_14267_),
    .B1_N(_14268_),
    .Y(_14269_));
 sky130_fd_sc_hd__nand3b_2 _35919_ (.A_N(_14265_),
    .B(_14268_),
    .C(_14266_),
    .Y(_14270_));
 sky130_fd_sc_hd__a21boi_2 _35920_ (.A1(_14032_),
    .A2(_14039_),
    .B1_N(_14033_),
    .Y(_14271_));
 sky130_vsdinv _35921_ (.A(_14271_),
    .Y(_14272_));
 sky130_fd_sc_hd__a21o_2 _35922_ (.A1(_14269_),
    .A2(_14270_),
    .B1(_14272_),
    .X(_14273_));
 sky130_fd_sc_hd__nand3_2 _35923_ (.A(_14269_),
    .B(_14270_),
    .C(_14272_),
    .Y(_14274_));
 sky130_fd_sc_hd__nand2_2 _35924_ (.A(_14273_),
    .B(_14274_),
    .Y(_14275_));
 sky130_fd_sc_hd__buf_1 _35925_ (.A(_14275_),
    .X(_14276_));
 sky130_fd_sc_hd__a21boi_2 _35926_ (.A1(_14240_),
    .A2(_14244_),
    .B1_N(_14276_),
    .Y(_14277_));
 sky130_fd_sc_hd__a21oi_2 _35927_ (.A1(_14241_),
    .A2(_14242_),
    .B1(_14239_),
    .Y(_14278_));
 sky130_fd_sc_hd__nor3b_2 _35928_ (.A(_14276_),
    .B(_14278_),
    .C_N(_14244_),
    .Y(_14279_));
 sky130_fd_sc_hd__o21ai_2 _35929_ (.A1(_14050_),
    .A2(_14052_),
    .B1(_14022_),
    .Y(_14280_));
 sky130_fd_sc_hd__o21bai_2 _35930_ (.A1(_14277_),
    .A2(_14279_),
    .B1_N(_14280_),
    .Y(_14281_));
 sky130_fd_sc_hd__nand2_2 _35931_ (.A(_14240_),
    .B(_14243_),
    .Y(_14282_));
 sky130_fd_sc_hd__nand2_2 _35932_ (.A(_14282_),
    .B(_14276_),
    .Y(_14283_));
 sky130_fd_sc_hd__nand3b_2 _35933_ (.A_N(_14275_),
    .B(_14240_),
    .C(_14244_),
    .Y(_14284_));
 sky130_fd_sc_hd__nand3_2 _35934_ (.A(_14283_),
    .B(_14284_),
    .C(_14280_),
    .Y(_14285_));
 sky130_fd_sc_hd__buf_1 _35935_ (.A(_14285_),
    .X(_14286_));
 sky130_fd_sc_hd__nand2_2 _35936_ (.A(_10356_),
    .B(_10551_),
    .Y(_14287_));
 sky130_fd_sc_hd__nand2_2 _35937_ (.A(_07474_),
    .B(_11791_),
    .Y(_14288_));
 sky130_fd_sc_hd__xor2_2 _35938_ (.A(_14287_),
    .B(_14288_),
    .X(_14289_));
 sky130_fd_sc_hd__nand3_2 _35939_ (.A(_14289_),
    .B(_06668_),
    .C(_10914_),
    .Y(_14290_));
 sky130_fd_sc_hd__xnor2_2 _35940_ (.A(_14287_),
    .B(_14288_),
    .Y(_14291_));
 sky130_fd_sc_hd__o21ai_2 _35941_ (.A1(_10780_),
    .A2(_19141_),
    .B1(_14291_),
    .Y(_14292_));
 sky130_fd_sc_hd__nand2_2 _35942_ (.A(_14290_),
    .B(_14292_),
    .Y(_14293_));
 sky130_fd_sc_hd__a21boi_2 _35943_ (.A1(_14037_),
    .A2(_14034_),
    .B1_N(_14036_),
    .Y(_14294_));
 sky130_fd_sc_hd__nand2_2 _35944_ (.A(_14293_),
    .B(_14294_),
    .Y(_14295_));
 sky130_fd_sc_hd__nand3b_2 _35945_ (.A_N(_14294_),
    .B(_14290_),
    .C(_14292_),
    .Y(_14296_));
 sky130_fd_sc_hd__o21ai_2 _35946_ (.A1(_14060_),
    .A2(_14061_),
    .B1(_14063_),
    .Y(_14297_));
 sky130_fd_sc_hd__a21oi_2 _35947_ (.A1(_14295_),
    .A2(_14296_),
    .B1(_14297_),
    .Y(_14298_));
 sky130_fd_sc_hd__nand3_2 _35948_ (.A(_14295_),
    .B(_14297_),
    .C(_14296_),
    .Y(_14299_));
 sky130_vsdinv _35949_ (.A(_14299_),
    .Y(_14300_));
 sky130_fd_sc_hd__o21ai_2 _35950_ (.A1(_14073_),
    .A2(_14070_),
    .B1(_14071_),
    .Y(_14301_));
 sky130_fd_sc_hd__o21bai_2 _35951_ (.A1(_14298_),
    .A2(_14300_),
    .B1_N(_14301_),
    .Y(_14302_));
 sky130_fd_sc_hd__nand3b_2 _35952_ (.A_N(_14298_),
    .B(_14299_),
    .C(_14301_),
    .Y(_14303_));
 sky130_fd_sc_hd__nand2_2 _35953_ (.A(_08414_),
    .B(_19132_),
    .Y(_14304_));
 sky130_fd_sc_hd__nand3b_2 _35954_ (.A_N(_14304_),
    .B(_12368_),
    .C(_06393_),
    .Y(_14305_));
 sky130_fd_sc_hd__nand2_2 _35955_ (.A(_11830_),
    .B(_09870_),
    .Y(_14306_));
 sky130_fd_sc_hd__nand2_2 _35956_ (.A(_14304_),
    .B(_14306_),
    .Y(_14307_));
 sky130_fd_sc_hd__and3_2 _35957_ (.A(_14305_),
    .B(_14084_),
    .C(_14307_),
    .X(_14308_));
 sky130_vsdinv _35958_ (.A(_14308_),
    .Y(_14309_));
 sky130_fd_sc_hd__o2bb2ai_2 _35959_ (.A1_N(_14307_),
    .A2_N(_14305_),
    .B1(_16963_),
    .B2(_18811_),
    .Y(_14310_));
 sky130_fd_sc_hd__nor2_2 _35960_ (.A(_14081_),
    .B(_14082_),
    .Y(_14311_));
 sky130_fd_sc_hd__o21bai_2 _35961_ (.A1(_14088_),
    .A2(_14087_),
    .B1_N(_14311_),
    .Y(_14312_));
 sky130_fd_sc_hd__a21oi_2 _35962_ (.A1(_14309_),
    .A2(_14310_),
    .B1(_14312_),
    .Y(_14313_));
 sky130_fd_sc_hd__nand3_2 _35963_ (.A(_14309_),
    .B(_14312_),
    .C(_14310_),
    .Y(_14314_));
 sky130_vsdinv _35964_ (.A(_14314_),
    .Y(_14315_));
 sky130_fd_sc_hd__buf_1 _35965_ (.A(_13863_),
    .X(_14316_));
 sky130_fd_sc_hd__o21bai_2 _35966_ (.A1(_14313_),
    .A2(_14315_),
    .B1_N(_14316_),
    .Y(_14317_));
 sky130_fd_sc_hd__a21o_2 _35967_ (.A1(_14309_),
    .A2(_14310_),
    .B1(_14312_),
    .X(_14318_));
 sky130_fd_sc_hd__nand3_2 _35968_ (.A(_14318_),
    .B(_14316_),
    .C(_14314_),
    .Y(_14319_));
 sky130_fd_sc_hd__nand2_2 _35969_ (.A(_14317_),
    .B(_14319_),
    .Y(_14320_));
 sky130_fd_sc_hd__a21boi_2 _35970_ (.A1(_14302_),
    .A2(_14303_),
    .B1_N(_14320_),
    .Y(_14321_));
 sky130_fd_sc_hd__nand2_2 _35971_ (.A(_14302_),
    .B(_14303_),
    .Y(_14322_));
 sky130_fd_sc_hd__nor2_2 _35972_ (.A(_14320_),
    .B(_14322_),
    .Y(_14323_));
 sky130_fd_sc_hd__nand2_2 _35973_ (.A(_14048_),
    .B(_14044_),
    .Y(_14324_));
 sky130_fd_sc_hd__o21bai_2 _35974_ (.A1(_14321_),
    .A2(_14323_),
    .B1_N(_14324_),
    .Y(_14325_));
 sky130_fd_sc_hd__nand3b_2 _35975_ (.A_N(_14320_),
    .B(_14303_),
    .C(_14302_),
    .Y(_14326_));
 sky130_fd_sc_hd__nand3b_2 _35976_ (.A_N(_14321_),
    .B(_14324_),
    .C(_14326_),
    .Y(_14327_));
 sky130_fd_sc_hd__a21boi_2 _35977_ (.A1(_14097_),
    .A2(_14079_),
    .B1_N(_14080_),
    .Y(_14328_));
 sky130_vsdinv _35978_ (.A(_14328_),
    .Y(_14329_));
 sky130_fd_sc_hd__a21o_2 _35979_ (.A1(_14325_),
    .A2(_14327_),
    .B1(_14329_),
    .X(_14330_));
 sky130_fd_sc_hd__nand3_2 _35980_ (.A(_14325_),
    .B(_14327_),
    .C(_14329_),
    .Y(_14331_));
 sky130_fd_sc_hd__nand2_2 _35981_ (.A(_14330_),
    .B(_14331_),
    .Y(_14332_));
 sky130_fd_sc_hd__buf_1 _35982_ (.A(_14332_),
    .X(_14333_));
 sky130_fd_sc_hd__a21boi_2 _35983_ (.A1(_14281_),
    .A2(_14286_),
    .B1_N(_14333_),
    .Y(_14334_));
 sky130_fd_sc_hd__a21oi_2 _35984_ (.A1(_14283_),
    .A2(_14284_),
    .B1(_14280_),
    .Y(_14335_));
 sky130_fd_sc_hd__nor3b_2 _35985_ (.A(_14333_),
    .B(_14335_),
    .C_N(_14286_),
    .Y(_14336_));
 sky130_fd_sc_hd__a21oi_2 _35986_ (.A1(_14057_),
    .A2(_14058_),
    .B1(_14055_),
    .Y(_14337_));
 sky130_fd_sc_hd__o21ai_2 _35987_ (.A1(_14112_),
    .A2(_14337_),
    .B1(_14059_),
    .Y(_14338_));
 sky130_fd_sc_hd__o21bai_2 _35988_ (.A1(_14334_),
    .A2(_14336_),
    .B1_N(_14338_),
    .Y(_14339_));
 sky130_vsdinv _35989_ (.A(_14285_),
    .Y(_14340_));
 sky130_fd_sc_hd__o21ai_2 _35990_ (.A1(_14335_),
    .A2(_14340_),
    .B1(_14333_),
    .Y(_14341_));
 sky130_fd_sc_hd__nand3b_2 _35991_ (.A_N(_14332_),
    .B(_14281_),
    .C(_14286_),
    .Y(_14342_));
 sky130_fd_sc_hd__nand3_2 _35992_ (.A(_14341_),
    .B(_14338_),
    .C(_14342_),
    .Y(_14343_));
 sky130_fd_sc_hd__buf_1 _35993_ (.A(_14343_),
    .X(_14344_));
 sky130_fd_sc_hd__nand2_2 _35994_ (.A(_14095_),
    .B(_14093_),
    .Y(_14345_));
 sky130_fd_sc_hd__nand2_2 _35995_ (.A(_14345_),
    .B(_14128_),
    .Y(_14346_));
 sky130_fd_sc_hd__buf_1 _35996_ (.A(_14125_),
    .X(_14347_));
 sky130_fd_sc_hd__buf_1 _35997_ (.A(_14126_),
    .X(_14348_));
 sky130_fd_sc_hd__o211ai_2 _35998_ (.A1(_14347_),
    .A2(_14348_),
    .B1(_14093_),
    .C1(_14095_),
    .Y(_14349_));
 sky130_fd_sc_hd__a21boi_2 _35999_ (.A1(_14123_),
    .A2(_13419_),
    .B1_N(_14124_),
    .Y(_14350_));
 sky130_vsdinv _36000_ (.A(_14350_),
    .Y(_14351_));
 sky130_fd_sc_hd__buf_1 _36001_ (.A(_14351_),
    .X(_14352_));
 sky130_fd_sc_hd__a21oi_2 _36002_ (.A1(_14346_),
    .A2(_14349_),
    .B1(_14352_),
    .Y(_14353_));
 sky130_fd_sc_hd__buf_1 _36003_ (.A(_14351_),
    .X(_14354_));
 sky130_fd_sc_hd__nand3_2 _36004_ (.A(_14346_),
    .B(_14349_),
    .C(_14354_),
    .Y(_14355_));
 sky130_vsdinv _36005_ (.A(_14355_),
    .Y(_14356_));
 sky130_fd_sc_hd__nand2_2 _36006_ (.A(_14134_),
    .B(_14129_),
    .Y(_14357_));
 sky130_fd_sc_hd__o21bai_2 _36007_ (.A1(_14353_),
    .A2(_14356_),
    .B1_N(_14357_),
    .Y(_14358_));
 sky130_fd_sc_hd__nand3b_2 _36008_ (.A_N(_14353_),
    .B(_14355_),
    .C(_14357_),
    .Y(_14359_));
 sky130_fd_sc_hd__buf_1 _36009_ (.A(_12944_),
    .X(_14360_));
 sky130_fd_sc_hd__a21o_2 _36010_ (.A1(_14358_),
    .A2(_14359_),
    .B1(_14360_),
    .X(_14361_));
 sky130_fd_sc_hd__nand3_2 _36011_ (.A(_14358_),
    .B(_14360_),
    .C(_14359_),
    .Y(_14362_));
 sky130_fd_sc_hd__nand2_2 _36012_ (.A(_14361_),
    .B(_14362_),
    .Y(_14363_));
 sky130_fd_sc_hd__a21boi_2 _36013_ (.A1(_14103_),
    .A2(_14109_),
    .B1_N(_14104_),
    .Y(_14364_));
 sky130_fd_sc_hd__nand2_2 _36014_ (.A(_14363_),
    .B(_14364_),
    .Y(_14365_));
 sky130_fd_sc_hd__nand2_2 _36015_ (.A(_14110_),
    .B(_14104_),
    .Y(_14366_));
 sky130_fd_sc_hd__nand3_2 _36016_ (.A(_14366_),
    .B(_14362_),
    .C(_14361_),
    .Y(_14367_));
 sky130_fd_sc_hd__a21boi_2 _36017_ (.A1(_14136_),
    .A2(_13194_),
    .B1_N(_14138_),
    .Y(_14368_));
 sky130_vsdinv _36018_ (.A(_14368_),
    .Y(_14369_));
 sky130_fd_sc_hd__a21o_2 _36019_ (.A1(_14365_),
    .A2(_14367_),
    .B1(_14369_),
    .X(_14370_));
 sky130_fd_sc_hd__nand3_2 _36020_ (.A(_14365_),
    .B(_14367_),
    .C(_14369_),
    .Y(_14371_));
 sky130_fd_sc_hd__nand2_2 _36021_ (.A(_14370_),
    .B(_14371_),
    .Y(_14372_));
 sky130_fd_sc_hd__a21boi_2 _36022_ (.A1(_14339_),
    .A2(_14344_),
    .B1_N(_14372_),
    .Y(_14373_));
 sky130_fd_sc_hd__a21oi_2 _36023_ (.A1(_14341_),
    .A2(_14342_),
    .B1(_14338_),
    .Y(_14374_));
 sky130_vsdinv _36024_ (.A(_14344_),
    .Y(_14375_));
 sky130_fd_sc_hd__nor3_2 _36025_ (.A(_14372_),
    .B(_14374_),
    .C(_14375_),
    .Y(_14376_));
 sky130_fd_sc_hd__o21ai_2 _36026_ (.A1(_14155_),
    .A2(_14156_),
    .B1(_14120_),
    .Y(_14377_));
 sky130_fd_sc_hd__o21bai_2 _36027_ (.A1(_14373_),
    .A2(_14376_),
    .B1_N(_14377_),
    .Y(_14378_));
 sky130_fd_sc_hd__nand2_2 _36028_ (.A(_14339_),
    .B(_14343_),
    .Y(_14379_));
 sky130_fd_sc_hd__nand2_2 _36029_ (.A(_14379_),
    .B(_14372_),
    .Y(_14380_));
 sky130_fd_sc_hd__and2_2 _36030_ (.A(_14370_),
    .B(_14371_),
    .X(_14381_));
 sky130_fd_sc_hd__nand3_2 _36031_ (.A(_14381_),
    .B(_14344_),
    .C(_14339_),
    .Y(_14382_));
 sky130_fd_sc_hd__nand3_2 _36032_ (.A(_14380_),
    .B(_14377_),
    .C(_14382_),
    .Y(_14383_));
 sky130_fd_sc_hd__nand2_2 _36033_ (.A(_14150_),
    .B(_14146_),
    .Y(_14384_));
 sky130_fd_sc_hd__xor2_2 _36034_ (.A(_13693_),
    .B(_14384_),
    .X(_14385_));
 sky130_fd_sc_hd__a21oi_2 _36035_ (.A1(_14378_),
    .A2(_14383_),
    .B1(_14385_),
    .Y(_14386_));
 sky130_vsdinv _36036_ (.A(_14385_),
    .Y(_14387_));
 sky130_fd_sc_hd__a21oi_2 _36037_ (.A1(_14380_),
    .A2(_14382_),
    .B1(_14377_),
    .Y(_14388_));
 sky130_vsdinv _36038_ (.A(_14383_),
    .Y(_14389_));
 sky130_fd_sc_hd__nor3_2 _36039_ (.A(_14387_),
    .B(_14388_),
    .C(_14389_),
    .Y(_14390_));
 sky130_fd_sc_hd__o21ai_2 _36040_ (.A1(_14167_),
    .A2(_14178_),
    .B1(_14169_),
    .Y(_14391_));
 sky130_fd_sc_hd__o21bai_2 _36041_ (.A1(_14386_),
    .A2(_14390_),
    .B1_N(_14391_),
    .Y(_14392_));
 sky130_fd_sc_hd__o21bai_2 _36042_ (.A1(_14388_),
    .A2(_14389_),
    .B1_N(_14385_),
    .Y(_14393_));
 sky130_fd_sc_hd__nand3_2 _36043_ (.A(_14378_),
    .B(_14385_),
    .C(_14383_),
    .Y(_14394_));
 sky130_fd_sc_hd__nand3_2 _36044_ (.A(_14393_),
    .B(_14394_),
    .C(_14391_),
    .Y(_14395_));
 sky130_fd_sc_hd__nand2_2 _36045_ (.A(_14392_),
    .B(_14395_),
    .Y(_14396_));
 sky130_fd_sc_hd__a21oi_2 _36046_ (.A1(_13922_),
    .A2(_13918_),
    .B1(_13952_),
    .Y(_14397_));
 sky130_vsdinv _36047_ (.A(_14397_),
    .Y(_14398_));
 sky130_fd_sc_hd__nand2_2 _36048_ (.A(_14396_),
    .B(_14398_),
    .Y(_14399_));
 sky130_fd_sc_hd__nand3_2 _36049_ (.A(_14392_),
    .B(_14397_),
    .C(_14395_),
    .Y(_14400_));
 sky130_vsdinv _36050_ (.A(_14175_),
    .Y(_14401_));
 sky130_fd_sc_hd__o21ai_2 _36051_ (.A1(_14401_),
    .A2(_14172_),
    .B1(_14173_),
    .Y(_14402_));
 sky130_fd_sc_hd__a21o_2 _36052_ (.A1(_14399_),
    .A2(_14400_),
    .B1(_14402_),
    .X(_14403_));
 sky130_fd_sc_hd__nand3_2 _36053_ (.A(_14399_),
    .B(_14402_),
    .C(_14400_),
    .Y(_14404_));
 sky130_fd_sc_hd__nand2_2 _36054_ (.A(_14403_),
    .B(_14404_),
    .Y(_14405_));
 sky130_fd_sc_hd__a21oi_2 _36055_ (.A1(_14180_),
    .A2(_14173_),
    .B1(_14175_),
    .Y(_14406_));
 sky130_fd_sc_hd__nor3_2 _36056_ (.A(_14401_),
    .B(_14172_),
    .C(_14174_),
    .Y(_14407_));
 sky130_fd_sc_hd__o21bai_2 _36057_ (.A1(_14406_),
    .A2(_14407_),
    .B1_N(_14182_),
    .Y(_14408_));
 sky130_fd_sc_hd__a21oi_2 _36058_ (.A1(_14194_),
    .A2(_14408_),
    .B1(_14185_),
    .Y(_14409_));
 sky130_fd_sc_hd__xor2_2 _36059_ (.A(_14405_),
    .B(_14409_),
    .X(_02664_));
 sky130_fd_sc_hd__nand2_2 _36060_ (.A(_10481_),
    .B(_08262_),
    .Y(_14410_));
 sky130_fd_sc_hd__buf_1 _36061_ (.A(_11599_),
    .X(_14411_));
 sky130_fd_sc_hd__nand3b_2 _36062_ (.A_N(_14410_),
    .B(_14411_),
    .C(_19232_),
    .Y(_14412_));
 sky130_fd_sc_hd__o21ai_2 _36063_ (.A1(_10743_),
    .A2(_11332_),
    .B1(_14410_),
    .Y(_14413_));
 sky130_fd_sc_hd__and2_2 _36064_ (.A(_18704_),
    .B(_10150_),
    .X(_14414_));
 sky130_fd_sc_hd__a21o_2 _36065_ (.A1(_14412_),
    .A2(_14413_),
    .B1(_14414_),
    .X(_14415_));
 sky130_fd_sc_hd__nand3_2 _36066_ (.A(_14412_),
    .B(_14413_),
    .C(_14414_),
    .Y(_14416_));
 sky130_fd_sc_hd__nand2_2 _36067_ (.A(_14200_),
    .B(_14196_),
    .Y(_14417_));
 sky130_fd_sc_hd__a21o_2 _36068_ (.A1(_14415_),
    .A2(_14416_),
    .B1(_14417_),
    .X(_14418_));
 sky130_fd_sc_hd__nand3_2 _36069_ (.A(_14417_),
    .B(_14415_),
    .C(_14416_),
    .Y(_14419_));
 sky130_fd_sc_hd__and2_2 _36070_ (.A(_09606_),
    .B(_07966_),
    .X(_14420_));
 sky130_fd_sc_hd__buf_1 _36071_ (.A(_14420_),
    .X(_14421_));
 sky130_fd_sc_hd__nand2_2 _36072_ (.A(_18711_),
    .B(_07118_),
    .Y(_14422_));
 sky130_fd_sc_hd__nand2_2 _36073_ (.A(_18717_),
    .B(_07944_),
    .Y(_14423_));
 sky130_fd_sc_hd__xnor2_2 _36074_ (.A(_14422_),
    .B(_14423_),
    .Y(_14424_));
 sky130_fd_sc_hd__xnor2_2 _36075_ (.A(_14421_),
    .B(_14424_),
    .Y(_14425_));
 sky130_fd_sc_hd__a21oi_2 _36076_ (.A1(_14418_),
    .A2(_14419_),
    .B1(_14425_),
    .Y(_14426_));
 sky130_fd_sc_hd__nand3_2 _36077_ (.A(_14418_),
    .B(_14425_),
    .C(_14419_),
    .Y(_14427_));
 sky130_vsdinv _36078_ (.A(_14427_),
    .Y(_14428_));
 sky130_fd_sc_hd__a21oi_2 _36079_ (.A1(_14199_),
    .A2(_14200_),
    .B1(_14201_),
    .Y(_14429_));
 sky130_fd_sc_hd__xor2_2 _36080_ (.A(_14205_),
    .B(_14208_),
    .X(_14430_));
 sky130_fd_sc_hd__o21ai_2 _36081_ (.A1(_14429_),
    .A2(_14430_),
    .B1(_14203_),
    .Y(_14431_));
 sky130_fd_sc_hd__o21bai_2 _36082_ (.A1(_14426_),
    .A2(_14428_),
    .B1_N(_14431_),
    .Y(_14432_));
 sky130_fd_sc_hd__a21o_2 _36083_ (.A1(_14418_),
    .A2(_14419_),
    .B1(_14425_),
    .X(_14433_));
 sky130_fd_sc_hd__nand3_2 _36084_ (.A(_14433_),
    .B(_14427_),
    .C(_14431_),
    .Y(_14434_));
 sky130_fd_sc_hd__nand2_2 _36085_ (.A(_10452_),
    .B(_08549_),
    .Y(_14435_));
 sky130_fd_sc_hd__nand2_2 _36086_ (.A(_11636_),
    .B(_12004_),
    .Y(_14436_));
 sky130_fd_sc_hd__xor2_2 _36087_ (.A(_14435_),
    .B(_14436_),
    .X(_14437_));
 sky130_fd_sc_hd__nand3_2 _36088_ (.A(_14437_),
    .B(_13508_),
    .C(_09105_),
    .Y(_14438_));
 sky130_fd_sc_hd__xnor2_2 _36089_ (.A(_14435_),
    .B(_14436_),
    .Y(_14439_));
 sky130_fd_sc_hd__o21ai_2 _36090_ (.A1(_10246_),
    .A2(_19187_),
    .B1(_14439_),
    .Y(_14440_));
 sky130_fd_sc_hd__nand2_2 _36091_ (.A(_14206_),
    .B(_14207_),
    .Y(_14441_));
 sky130_fd_sc_hd__nor2_2 _36092_ (.A(_14206_),
    .B(_14207_),
    .Y(_14442_));
 sky130_fd_sc_hd__a21oi_2 _36093_ (.A1(_14441_),
    .A2(_14205_),
    .B1(_14442_),
    .Y(_14443_));
 sky130_fd_sc_hd__a21bo_2 _36094_ (.A1(_14438_),
    .A2(_14440_),
    .B1_N(_14443_),
    .X(_14444_));
 sky130_fd_sc_hd__nand3b_2 _36095_ (.A_N(_14443_),
    .B(_14438_),
    .C(_14440_),
    .Y(_14445_));
 sky130_fd_sc_hd__o21ai_2 _36096_ (.A1(_14219_),
    .A2(_14220_),
    .B1(_14222_),
    .Y(_14446_));
 sky130_fd_sc_hd__a21o_2 _36097_ (.A1(_14444_),
    .A2(_14445_),
    .B1(_14446_),
    .X(_14447_));
 sky130_fd_sc_hd__nand3_2 _36098_ (.A(_14444_),
    .B(_14446_),
    .C(_14445_),
    .Y(_14448_));
 sky130_fd_sc_hd__nand2_2 _36099_ (.A(_14447_),
    .B(_14448_),
    .Y(_14449_));
 sky130_fd_sc_hd__buf_1 _36100_ (.A(_14449_),
    .X(_14450_));
 sky130_fd_sc_hd__a21boi_2 _36101_ (.A1(_14432_),
    .A2(_14434_),
    .B1_N(_14450_),
    .Y(_14451_));
 sky130_fd_sc_hd__a21oi_2 _36102_ (.A1(_14433_),
    .A2(_14427_),
    .B1(_14431_),
    .Y(_14452_));
 sky130_vsdinv _36103_ (.A(_14434_),
    .Y(_14453_));
 sky130_fd_sc_hd__nor3_2 _36104_ (.A(_14450_),
    .B(_14452_),
    .C(_14453_),
    .Y(_14454_));
 sky130_fd_sc_hd__o21ai_2 _36105_ (.A1(_14234_),
    .A2(_14236_),
    .B1(_14218_),
    .Y(_14455_));
 sky130_fd_sc_hd__o21bai_2 _36106_ (.A1(_14451_),
    .A2(_14454_),
    .B1_N(_14455_),
    .Y(_14456_));
 sky130_fd_sc_hd__o21ai_2 _36107_ (.A1(_14452_),
    .A2(_14453_),
    .B1(_14450_),
    .Y(_14457_));
 sky130_fd_sc_hd__nand3b_2 _36108_ (.A_N(_14449_),
    .B(_14432_),
    .C(_14434_),
    .Y(_14458_));
 sky130_fd_sc_hd__nand3_2 _36109_ (.A(_14457_),
    .B(_14458_),
    .C(_14455_),
    .Y(_14459_));
 sky130_fd_sc_hd__buf_1 _36110_ (.A(_14459_),
    .X(_14460_));
 sky130_fd_sc_hd__nand2_2 _36111_ (.A(_10421_),
    .B(_09492_),
    .Y(_14461_));
 sky130_fd_sc_hd__nand2_2 _36112_ (.A(_08731_),
    .B(_09493_),
    .Y(_14462_));
 sky130_fd_sc_hd__xor2_2 _36113_ (.A(_14461_),
    .B(_14462_),
    .X(_14463_));
 sky130_fd_sc_hd__and2_2 _36114_ (.A(_08085_),
    .B(_12325_),
    .X(_14464_));
 sky130_fd_sc_hd__nand2_2 _36115_ (.A(_14463_),
    .B(_14464_),
    .Y(_14465_));
 sky130_fd_sc_hd__xnor2_2 _36116_ (.A(_14461_),
    .B(_14462_),
    .Y(_14466_));
 sky130_fd_sc_hd__o21ai_2 _36117_ (.A1(_08232_),
    .A2(_19169_),
    .B1(_14466_),
    .Y(_14467_));
 sky130_fd_sc_hd__a21oi_2 _36118_ (.A1(_14248_),
    .A2(_14252_),
    .B1(_14249_),
    .Y(_14468_));
 sky130_vsdinv _36119_ (.A(_14468_),
    .Y(_14469_));
 sky130_fd_sc_hd__a21o_2 _36120_ (.A1(_14465_),
    .A2(_14467_),
    .B1(_14469_),
    .X(_14470_));
 sky130_fd_sc_hd__nand3_2 _36121_ (.A(_14465_),
    .B(_14467_),
    .C(_14469_),
    .Y(_14471_));
 sky130_fd_sc_hd__and2_2 _36122_ (.A(_07162_),
    .B(_13113_),
    .X(_14472_));
 sky130_fd_sc_hd__nand2_2 _36123_ (.A(_12806_),
    .B(_11788_),
    .Y(_14473_));
 sky130_fd_sc_hd__nand3b_2 _36124_ (.A_N(_14473_),
    .B(_18766_),
    .C(_10043_),
    .Y(_14474_));
 sky130_fd_sc_hd__a22o_2 _36125_ (.A1(_12847_),
    .A2(_09809_),
    .B1(_10430_),
    .B2(_10052_),
    .X(_14475_));
 sky130_fd_sc_hd__nand2_2 _36126_ (.A(_14474_),
    .B(_14475_),
    .Y(_14476_));
 sky130_fd_sc_hd__xnor2_2 _36127_ (.A(_14472_),
    .B(_14476_),
    .Y(_14477_));
 sky130_fd_sc_hd__a21oi_2 _36128_ (.A1(_14470_),
    .A2(_14471_),
    .B1(_14477_),
    .Y(_14478_));
 sky130_fd_sc_hd__nand3_2 _36129_ (.A(_14470_),
    .B(_14477_),
    .C(_14471_),
    .Y(_14479_));
 sky130_vsdinv _36130_ (.A(_14479_),
    .Y(_14480_));
 sky130_fd_sc_hd__nand2_2 _36131_ (.A(_14232_),
    .B(_14229_),
    .Y(_14481_));
 sky130_fd_sc_hd__o21bai_2 _36132_ (.A1(_14478_),
    .A2(_14480_),
    .B1_N(_14481_),
    .Y(_14482_));
 sky130_fd_sc_hd__nand3b_2 _36133_ (.A_N(_14478_),
    .B(_14481_),
    .C(_14479_),
    .Y(_14483_));
 sky130_vsdinv _36134_ (.A(_14258_),
    .Y(_14484_));
 sky130_fd_sc_hd__a21oi_2 _36135_ (.A1(_14257_),
    .A2(_14264_),
    .B1(_14484_),
    .Y(_14485_));
 sky130_vsdinv _36136_ (.A(_14485_),
    .Y(_14486_));
 sky130_fd_sc_hd__a21oi_2 _36137_ (.A1(_14482_),
    .A2(_14483_),
    .B1(_14486_),
    .Y(_14487_));
 sky130_fd_sc_hd__nand3_2 _36138_ (.A(_14482_),
    .B(_14486_),
    .C(_14483_),
    .Y(_14488_));
 sky130_vsdinv _36139_ (.A(_14488_),
    .Y(_14489_));
 sky130_fd_sc_hd__nor2_2 _36140_ (.A(_14487_),
    .B(_14489_),
    .Y(_14490_));
 sky130_fd_sc_hd__a21oi_2 _36141_ (.A1(_14456_),
    .A2(_14460_),
    .B1(_14490_),
    .Y(_14491_));
 sky130_fd_sc_hd__nand2_2 _36142_ (.A(_14482_),
    .B(_14483_),
    .Y(_14492_));
 sky130_fd_sc_hd__nand2_2 _36143_ (.A(_14492_),
    .B(_14485_),
    .Y(_14493_));
 sky130_fd_sc_hd__nand2_2 _36144_ (.A(_14493_),
    .B(_14488_),
    .Y(_14494_));
 sky130_fd_sc_hd__a21oi_2 _36145_ (.A1(_14457_),
    .A2(_14458_),
    .B1(_14455_),
    .Y(_14495_));
 sky130_vsdinv _36146_ (.A(_14460_),
    .Y(_14496_));
 sky130_fd_sc_hd__nor3_2 _36147_ (.A(_14494_),
    .B(_14495_),
    .C(_14496_),
    .Y(_14497_));
 sky130_fd_sc_hd__o21ai_2 _36148_ (.A1(_14276_),
    .A2(_14278_),
    .B1(_14244_),
    .Y(_14498_));
 sky130_fd_sc_hd__o21bai_2 _36149_ (.A1(_14491_),
    .A2(_14497_),
    .B1_N(_14498_),
    .Y(_14499_));
 sky130_fd_sc_hd__o2bb2ai_2 _36150_ (.A1_N(_14460_),
    .A2_N(_14456_),
    .B1(_14489_),
    .B2(_14487_),
    .Y(_14500_));
 sky130_fd_sc_hd__nand3_2 _36151_ (.A(_14490_),
    .B(_14460_),
    .C(_14456_),
    .Y(_14501_));
 sky130_fd_sc_hd__nand3_2 _36152_ (.A(_14500_),
    .B(_14501_),
    .C(_14498_),
    .Y(_14502_));
 sky130_fd_sc_hd__buf_1 _36153_ (.A(_14502_),
    .X(_14503_));
 sky130_fd_sc_hd__nand2_2 _36154_ (.A(_10777_),
    .B(_19144_),
    .Y(_14504_));
 sky130_fd_sc_hd__nand2_2 _36155_ (.A(_12289_),
    .B(_19139_),
    .Y(_14505_));
 sky130_fd_sc_hd__xor2_2 _36156_ (.A(_14504_),
    .B(_14505_),
    .X(_14506_));
 sky130_fd_sc_hd__nand3_2 _36157_ (.A(_14506_),
    .B(_06668_),
    .C(_19134_),
    .Y(_14507_));
 sky130_fd_sc_hd__xnor2_2 _36158_ (.A(_14504_),
    .B(_14505_),
    .Y(_14508_));
 sky130_fd_sc_hd__o21ai_2 _36159_ (.A1(_18793_),
    .A2(_12389_),
    .B1(_14508_),
    .Y(_14509_));
 sky130_fd_sc_hd__a21boi_2 _36160_ (.A1(_14262_),
    .A2(_14259_),
    .B1_N(_14261_),
    .Y(_14510_));
 sky130_fd_sc_hd__a21boi_2 _36161_ (.A1(_14507_),
    .A2(_14509_),
    .B1_N(_14510_),
    .Y(_14511_));
 sky130_fd_sc_hd__nand3b_2 _36162_ (.A_N(_14510_),
    .B(_14507_),
    .C(_14509_),
    .Y(_14512_));
 sky130_vsdinv _36163_ (.A(_14512_),
    .Y(_14513_));
 sky130_fd_sc_hd__o21ai_2 _36164_ (.A1(_14287_),
    .A2(_14288_),
    .B1(_14290_),
    .Y(_14514_));
 sky130_fd_sc_hd__o21bai_2 _36165_ (.A1(_14511_),
    .A2(_14513_),
    .B1_N(_14514_),
    .Y(_14515_));
 sky130_fd_sc_hd__a21bo_2 _36166_ (.A1(_14507_),
    .A2(_14509_),
    .B1_N(_14510_),
    .X(_14516_));
 sky130_fd_sc_hd__nand3_2 _36167_ (.A(_14516_),
    .B(_14514_),
    .C(_14512_),
    .Y(_14517_));
 sky130_fd_sc_hd__nand2_2 _36168_ (.A(_14299_),
    .B(_14296_),
    .Y(_14518_));
 sky130_fd_sc_hd__a21o_2 _36169_ (.A1(_14515_),
    .A2(_14517_),
    .B1(_14518_),
    .X(_14519_));
 sky130_fd_sc_hd__nand3_2 _36170_ (.A(_14515_),
    .B(_14518_),
    .C(_14517_),
    .Y(_14520_));
 sky130_fd_sc_hd__a21boi_2 _36171_ (.A1(_14085_),
    .A2(_14307_),
    .B1_N(_14305_),
    .Y(_14521_));
 sky130_fd_sc_hd__buf_1 _36172_ (.A(_10881_),
    .X(_14522_));
 sky130_fd_sc_hd__nand2_2 _36173_ (.A(_14522_),
    .B(_06545_),
    .Y(_14523_));
 sky130_fd_sc_hd__nand2_2 _36174_ (.A(_14306_),
    .B(_14523_),
    .Y(_14524_));
 sky130_fd_sc_hd__nand3_2 _36175_ (.A(_11204_),
    .B(_06535_),
    .C(_08043_),
    .Y(_14525_));
 sky130_fd_sc_hd__a21boi_2 _36176_ (.A1(_14524_),
    .A2(_14525_),
    .B1_N(_14085_),
    .Y(_14526_));
 sky130_fd_sc_hd__o211a_2 _36177_ (.A1(_16962_),
    .A2(_18810_),
    .B1(_14525_),
    .C1(_14524_),
    .X(_14527_));
 sky130_fd_sc_hd__nor2_2 _36178_ (.A(_14526_),
    .B(_14527_),
    .Y(_14528_));
 sky130_fd_sc_hd__or2b_2 _36179_ (.A(_14521_),
    .B_N(_14528_),
    .X(_14529_));
 sky130_fd_sc_hd__o21ai_2 _36180_ (.A1(_14527_),
    .A2(_14526_),
    .B1(_14521_),
    .Y(_14530_));
 sky130_vsdinv _36181_ (.A(_13864_),
    .Y(_14531_));
 sky130_fd_sc_hd__a21oi_2 _36182_ (.A1(_14529_),
    .A2(_14530_),
    .B1(_14531_),
    .Y(_14532_));
 sky130_fd_sc_hd__o211a_2 _36183_ (.A1(_13860_),
    .A2(_13861_),
    .B1(_14530_),
    .C1(_14529_),
    .X(_14533_));
 sky130_fd_sc_hd__nor2_2 _36184_ (.A(_14532_),
    .B(_14533_),
    .Y(_14534_));
 sky130_fd_sc_hd__a21oi_2 _36185_ (.A1(_14519_),
    .A2(_14520_),
    .B1(_14534_),
    .Y(_14535_));
 sky130_fd_sc_hd__nand3_2 _36186_ (.A(_14519_),
    .B(_14534_),
    .C(_14520_),
    .Y(_14536_));
 sky130_vsdinv _36187_ (.A(_14536_),
    .Y(_14537_));
 sky130_fd_sc_hd__a21boi_2 _36188_ (.A1(_14269_),
    .A2(_14272_),
    .B1_N(_14270_),
    .Y(_14538_));
 sky130_fd_sc_hd__o21ai_2 _36189_ (.A1(_14535_),
    .A2(_14537_),
    .B1(_14538_),
    .Y(_14539_));
 sky130_fd_sc_hd__o2bb2ai_2 _36190_ (.A1_N(_14520_),
    .A2_N(_14519_),
    .B1(_14532_),
    .B2(_14533_),
    .Y(_14540_));
 sky130_fd_sc_hd__nand3b_2 _36191_ (.A_N(_14538_),
    .B(_14536_),
    .C(_14540_),
    .Y(_14541_));
 sky130_fd_sc_hd__o21a_2 _36192_ (.A1(_14320_),
    .A2(_14322_),
    .B1(_14303_),
    .X(_14542_));
 sky130_vsdinv _36193_ (.A(_14542_),
    .Y(_14543_));
 sky130_fd_sc_hd__a21oi_2 _36194_ (.A1(_14539_),
    .A2(_14541_),
    .B1(_14543_),
    .Y(_14544_));
 sky130_fd_sc_hd__nand3_2 _36195_ (.A(_14539_),
    .B(_14543_),
    .C(_14541_),
    .Y(_14545_));
 sky130_vsdinv _36196_ (.A(_14545_),
    .Y(_14546_));
 sky130_fd_sc_hd__nor2_2 _36197_ (.A(_14544_),
    .B(_14546_),
    .Y(_14547_));
 sky130_fd_sc_hd__a21oi_2 _36198_ (.A1(_14499_),
    .A2(_14503_),
    .B1(_14547_),
    .Y(_14548_));
 sky130_fd_sc_hd__a21boi_2 _36199_ (.A1(_14540_),
    .A2(_14536_),
    .B1_N(_14538_),
    .Y(_14549_));
 sky130_fd_sc_hd__nor3_2 _36200_ (.A(_14538_),
    .B(_14535_),
    .C(_14537_),
    .Y(_14550_));
 sky130_fd_sc_hd__o21bai_2 _36201_ (.A1(_14549_),
    .A2(_14550_),
    .B1_N(_14543_),
    .Y(_14551_));
 sky130_fd_sc_hd__nand2_2 _36202_ (.A(_14551_),
    .B(_14545_),
    .Y(_14552_));
 sky130_fd_sc_hd__a21oi_2 _36203_ (.A1(_14500_),
    .A2(_14501_),
    .B1(_14498_),
    .Y(_14553_));
 sky130_vsdinv _36204_ (.A(_14503_),
    .Y(_14554_));
 sky130_fd_sc_hd__nor3_2 _36205_ (.A(_14552_),
    .B(_14553_),
    .C(_14554_),
    .Y(_14555_));
 sky130_fd_sc_hd__o21ai_2 _36206_ (.A1(_14333_),
    .A2(_14335_),
    .B1(_14286_),
    .Y(_14556_));
 sky130_fd_sc_hd__o21bai_2 _36207_ (.A1(_14548_),
    .A2(_14555_),
    .B1_N(_14556_),
    .Y(_14557_));
 sky130_fd_sc_hd__nand2_2 _36208_ (.A(_14499_),
    .B(_14502_),
    .Y(_14558_));
 sky130_fd_sc_hd__nand2_2 _36209_ (.A(_14558_),
    .B(_14552_),
    .Y(_14559_));
 sky130_fd_sc_hd__nand3_2 _36210_ (.A(_14547_),
    .B(_14499_),
    .C(_14503_),
    .Y(_14560_));
 sky130_fd_sc_hd__nand3_2 _36211_ (.A(_14559_),
    .B(_14560_),
    .C(_14556_),
    .Y(_14561_));
 sky130_fd_sc_hd__buf_1 _36212_ (.A(_14561_),
    .X(_14562_));
 sky130_fd_sc_hd__o211ai_2 _36213_ (.A1(_14347_),
    .A2(_14348_),
    .B1(_14314_),
    .C1(_14319_),
    .Y(_14563_));
 sky130_fd_sc_hd__o21ai_2 _36214_ (.A1(_14531_),
    .A2(_14313_),
    .B1(_14314_),
    .Y(_14564_));
 sky130_fd_sc_hd__nand2_2 _36215_ (.A(_14128_),
    .B(_14564_),
    .Y(_14565_));
 sky130_fd_sc_hd__nand3_2 _36216_ (.A(_14563_),
    .B(_14565_),
    .C(_14354_),
    .Y(_14566_));
 sky130_vsdinv _36217_ (.A(_14566_),
    .Y(_14567_));
 sky130_fd_sc_hd__a21oi_2 _36218_ (.A1(_14563_),
    .A2(_14565_),
    .B1(_14352_),
    .Y(_14568_));
 sky130_fd_sc_hd__nand2_2 _36219_ (.A(_14355_),
    .B(_14346_),
    .Y(_14569_));
 sky130_fd_sc_hd__o21bai_2 _36220_ (.A1(_14567_),
    .A2(_14568_),
    .B1_N(_14569_),
    .Y(_14570_));
 sky130_fd_sc_hd__nand3b_2 _36221_ (.A_N(_14568_),
    .B(_14566_),
    .C(_14569_),
    .Y(_14571_));
 sky130_fd_sc_hd__a21o_2 _36222_ (.A1(_14570_),
    .A2(_14571_),
    .B1(_13193_),
    .X(_14572_));
 sky130_fd_sc_hd__nand3_2 _36223_ (.A(_14570_),
    .B(_14360_),
    .C(_14571_),
    .Y(_14573_));
 sky130_fd_sc_hd__nand2_2 _36224_ (.A(_14331_),
    .B(_14327_),
    .Y(_14574_));
 sky130_fd_sc_hd__a21o_2 _36225_ (.A1(_14572_),
    .A2(_14573_),
    .B1(_14574_),
    .X(_14575_));
 sky130_fd_sc_hd__nand3_2 _36226_ (.A(_14574_),
    .B(_14572_),
    .C(_14573_),
    .Y(_14576_));
 sky130_fd_sc_hd__buf_1 _36227_ (.A(_14576_),
    .X(_14577_));
 sky130_fd_sc_hd__a21boi_2 _36228_ (.A1(_14358_),
    .A2(_13440_),
    .B1_N(_14359_),
    .Y(_14578_));
 sky130_vsdinv _36229_ (.A(_14578_),
    .Y(_14579_));
 sky130_fd_sc_hd__a21oi_2 _36230_ (.A1(_14575_),
    .A2(_14577_),
    .B1(_14579_),
    .Y(_14580_));
 sky130_fd_sc_hd__nand3_2 _36231_ (.A(_14575_),
    .B(_14579_),
    .C(_14576_),
    .Y(_14581_));
 sky130_vsdinv _36232_ (.A(_14581_),
    .Y(_14582_));
 sky130_fd_sc_hd__nor2_2 _36233_ (.A(_14580_),
    .B(_14582_),
    .Y(_14583_));
 sky130_fd_sc_hd__a21oi_2 _36234_ (.A1(_14557_),
    .A2(_14562_),
    .B1(_14583_),
    .Y(_14584_));
 sky130_fd_sc_hd__nand2_2 _36235_ (.A(_14575_),
    .B(_14577_),
    .Y(_14585_));
 sky130_fd_sc_hd__nand2_2 _36236_ (.A(_14585_),
    .B(_14578_),
    .Y(_14586_));
 sky130_fd_sc_hd__nand2_2 _36237_ (.A(_14586_),
    .B(_14581_),
    .Y(_14587_));
 sky130_fd_sc_hd__a21oi_2 _36238_ (.A1(_14559_),
    .A2(_14560_),
    .B1(_14556_),
    .Y(_14588_));
 sky130_vsdinv _36239_ (.A(_14562_),
    .Y(_14589_));
 sky130_fd_sc_hd__nor3_2 _36240_ (.A(_14587_),
    .B(_14588_),
    .C(_14589_),
    .Y(_14590_));
 sky130_fd_sc_hd__o21ai_2 _36241_ (.A1(_14372_),
    .A2(_14374_),
    .B1(_14344_),
    .Y(_14591_));
 sky130_fd_sc_hd__o21bai_2 _36242_ (.A1(_14584_),
    .A2(_14590_),
    .B1_N(_14591_),
    .Y(_14592_));
 sky130_fd_sc_hd__nand2_2 _36243_ (.A(_14557_),
    .B(_14561_),
    .Y(_14593_));
 sky130_fd_sc_hd__nand2_2 _36244_ (.A(_14593_),
    .B(_14587_),
    .Y(_14594_));
 sky130_fd_sc_hd__nand3_2 _36245_ (.A(_14583_),
    .B(_14557_),
    .C(_14562_),
    .Y(_14595_));
 sky130_fd_sc_hd__nand3_2 _36246_ (.A(_14594_),
    .B(_14595_),
    .C(_14591_),
    .Y(_14596_));
 sky130_fd_sc_hd__buf_1 _36247_ (.A(_14596_),
    .X(_14597_));
 sky130_fd_sc_hd__nand2_2 _36248_ (.A(_14371_),
    .B(_14367_),
    .Y(_14598_));
 sky130_fd_sc_hd__xor2_2 _36249_ (.A(_13693_),
    .B(_14598_),
    .X(_14599_));
 sky130_fd_sc_hd__a21oi_2 _36250_ (.A1(_14592_),
    .A2(_14597_),
    .B1(_14599_),
    .Y(_14600_));
 sky130_vsdinv _36251_ (.A(_14599_),
    .Y(_14601_));
 sky130_fd_sc_hd__a21oi_2 _36252_ (.A1(_14594_),
    .A2(_14595_),
    .B1(_14591_),
    .Y(_14602_));
 sky130_vsdinv _36253_ (.A(_14597_),
    .Y(_14603_));
 sky130_fd_sc_hd__nor3_2 _36254_ (.A(_14601_),
    .B(_14602_),
    .C(_14603_),
    .Y(_14604_));
 sky130_fd_sc_hd__o21ai_2 _36255_ (.A1(_14387_),
    .A2(_14388_),
    .B1(_14383_),
    .Y(_14605_));
 sky130_fd_sc_hd__o21bai_2 _36256_ (.A1(_14600_),
    .A2(_14604_),
    .B1_N(_14605_),
    .Y(_14606_));
 sky130_fd_sc_hd__nand2_2 _36257_ (.A(_14592_),
    .B(_14596_),
    .Y(_14607_));
 sky130_fd_sc_hd__nand2_2 _36258_ (.A(_14607_),
    .B(_14601_),
    .Y(_14608_));
 sky130_fd_sc_hd__nand3_2 _36259_ (.A(_14592_),
    .B(_14599_),
    .C(_14597_),
    .Y(_14609_));
 sky130_fd_sc_hd__nand3_2 _36260_ (.A(_14608_),
    .B(_14609_),
    .C(_14605_),
    .Y(_14610_));
 sky130_fd_sc_hd__a21oi_2 _36261_ (.A1(_14150_),
    .A2(_14146_),
    .B1(_13952_),
    .Y(_14611_));
 sky130_fd_sc_hd__a21oi_2 _36262_ (.A1(_14606_),
    .A2(_14610_),
    .B1(_14611_),
    .Y(_14612_));
 sky130_vsdinv _36263_ (.A(_14611_),
    .Y(_14613_));
 sky130_fd_sc_hd__a21oi_2 _36264_ (.A1(_14608_),
    .A2(_14609_),
    .B1(_14605_),
    .Y(_14614_));
 sky130_vsdinv _36265_ (.A(_14610_),
    .Y(_14615_));
 sky130_fd_sc_hd__nor3_2 _36266_ (.A(_14613_),
    .B(_14614_),
    .C(_14615_),
    .Y(_14616_));
 sky130_fd_sc_hd__a21oi_2 _36267_ (.A1(_14393_),
    .A2(_14394_),
    .B1(_14391_),
    .Y(_14617_));
 sky130_fd_sc_hd__o21ai_2 _36268_ (.A1(_14398_),
    .A2(_14617_),
    .B1(_14395_),
    .Y(_14618_));
 sky130_fd_sc_hd__o21bai_2 _36269_ (.A1(_14612_),
    .A2(_14616_),
    .B1_N(_14618_),
    .Y(_14619_));
 sky130_fd_sc_hd__o21bai_2 _36270_ (.A1(_14614_),
    .A2(_14615_),
    .B1_N(_14611_),
    .Y(_14620_));
 sky130_fd_sc_hd__nand3_2 _36271_ (.A(_14606_),
    .B(_14611_),
    .C(_14610_),
    .Y(_14621_));
 sky130_fd_sc_hd__nand3_2 _36272_ (.A(_14620_),
    .B(_14618_),
    .C(_14621_),
    .Y(_14622_));
 sky130_fd_sc_hd__nand2_2 _36273_ (.A(_14619_),
    .B(_14622_),
    .Y(_14623_));
 sky130_fd_sc_hd__nand2_2 _36274_ (.A(_14408_),
    .B(_14184_),
    .Y(_14624_));
 sky130_fd_sc_hd__nor2_2 _36275_ (.A(_14624_),
    .B(_14405_),
    .Y(_14625_));
 sky130_fd_sc_hd__a21oi_2 _36276_ (.A1(_14399_),
    .A2(_14400_),
    .B1(_14402_),
    .Y(_14626_));
 sky130_fd_sc_hd__a21oi_2 _36277_ (.A1(_14184_),
    .A2(_14404_),
    .B1(_14626_),
    .Y(_14627_));
 sky130_fd_sc_hd__a21oi_2 _36278_ (.A1(_14194_),
    .A2(_14625_),
    .B1(_14627_),
    .Y(_14628_));
 sky130_fd_sc_hd__xor2_2 _36279_ (.A(_14623_),
    .B(_14628_),
    .X(_02665_));
 sky130_fd_sc_hd__nand2_2 _36280_ (.A(_10777_),
    .B(_19139_),
    .Y(_14629_));
 sky130_fd_sc_hd__nand2_2 _36281_ (.A(_18786_),
    .B(_19133_),
    .Y(_14630_));
 sky130_fd_sc_hd__xnor2_2 _36282_ (.A(_14629_),
    .B(_14630_),
    .Y(_14631_));
 sky130_fd_sc_hd__and2_2 _36283_ (.A(_11830_),
    .B(_06666_),
    .X(_14632_));
 sky130_fd_sc_hd__buf_1 _36284_ (.A(_14632_),
    .X(_14633_));
 sky130_vsdinv _36285_ (.A(_14633_),
    .Y(_14634_));
 sky130_fd_sc_hd__nand2_2 _36286_ (.A(_14631_),
    .B(_14634_),
    .Y(_14635_));
 sky130_fd_sc_hd__xor2_2 _36287_ (.A(_14629_),
    .B(_14630_),
    .X(_14636_));
 sky130_fd_sc_hd__nand2_2 _36288_ (.A(_14636_),
    .B(_14633_),
    .Y(_14637_));
 sky130_fd_sc_hd__a21boi_2 _36289_ (.A1(_14475_),
    .A2(_14472_),
    .B1_N(_14474_),
    .Y(_14638_));
 sky130_fd_sc_hd__a21bo_2 _36290_ (.A1(_14635_),
    .A2(_14637_),
    .B1_N(_14638_),
    .X(_14639_));
 sky130_fd_sc_hd__nand3b_2 _36291_ (.A_N(_14638_),
    .B(_14635_),
    .C(_14637_),
    .Y(_14640_));
 sky130_fd_sc_hd__o21a_2 _36292_ (.A1(_14504_),
    .A2(_14505_),
    .B1(_14507_),
    .X(_14641_));
 sky130_fd_sc_hd__a21bo_2 _36293_ (.A1(_14639_),
    .A2(_14640_),
    .B1_N(_14641_),
    .X(_14642_));
 sky130_fd_sc_hd__nand3b_2 _36294_ (.A_N(_14641_),
    .B(_14639_),
    .C(_14640_),
    .Y(_14643_));
 sky130_fd_sc_hd__a21o_2 _36295_ (.A1(_14516_),
    .A2(_14514_),
    .B1(_14513_),
    .X(_14644_));
 sky130_fd_sc_hd__a21o_2 _36296_ (.A1(_14642_),
    .A2(_14643_),
    .B1(_14644_),
    .X(_14645_));
 sky130_fd_sc_hd__nand3_2 _36297_ (.A(_14642_),
    .B(_14644_),
    .C(_14643_),
    .Y(_14646_));
 sky130_fd_sc_hd__nand2_2 _36298_ (.A(_14645_),
    .B(_14646_),
    .Y(_14647_));
 sky130_fd_sc_hd__buf_1 _36299_ (.A(_12099_),
    .X(_14648_));
 sky130_fd_sc_hd__and4_2 _36300_ (.A(_14648_),
    .B(_18799_),
    .C(_06538_),
    .D(_06276_),
    .X(_14649_));
 sky130_fd_sc_hd__o21ba_2 _36301_ (.A1(_14085_),
    .A2(_14524_),
    .B1_N(_14649_),
    .X(_14650_));
 sky130_fd_sc_hd__xor2_2 _36302_ (.A(_14650_),
    .B(_13864_),
    .X(_14651_));
 sky130_vsdinv _36303_ (.A(_14651_),
    .Y(_14652_));
 sky130_fd_sc_hd__buf_1 _36304_ (.A(_14652_),
    .X(_14653_));
 sky130_fd_sc_hd__nand2_2 _36305_ (.A(_14647_),
    .B(_14653_),
    .Y(_14654_));
 sky130_fd_sc_hd__buf_1 _36306_ (.A(_14651_),
    .X(_14655_));
 sky130_fd_sc_hd__buf_1 _36307_ (.A(_14655_),
    .X(_14656_));
 sky130_fd_sc_hd__nand3_2 _36308_ (.A(_14645_),
    .B(_14656_),
    .C(_14646_),
    .Y(_14657_));
 sky130_fd_sc_hd__nand2_2 _36309_ (.A(_14488_),
    .B(_14483_),
    .Y(_14658_));
 sky130_fd_sc_hd__a21o_2 _36310_ (.A1(_14654_),
    .A2(_14657_),
    .B1(_14658_),
    .X(_14659_));
 sky130_vsdinv _36311_ (.A(_14520_),
    .Y(_14660_));
 sky130_fd_sc_hd__a21oi_2 _36312_ (.A1(_14519_),
    .A2(_14534_),
    .B1(_14660_),
    .Y(_14661_));
 sky130_vsdinv _36313_ (.A(_14661_),
    .Y(_14662_));
 sky130_fd_sc_hd__nand3_2 _36314_ (.A(_14658_),
    .B(_14654_),
    .C(_14657_),
    .Y(_14663_));
 sky130_fd_sc_hd__nand3_2 _36315_ (.A(_14659_),
    .B(_14662_),
    .C(_14663_),
    .Y(_14664_));
 sky130_fd_sc_hd__a21o_2 _36316_ (.A1(_14659_),
    .A2(_14663_),
    .B1(_14662_),
    .X(_14665_));
 sky130_fd_sc_hd__buf_1 _36317_ (.A(_10043_),
    .X(_14666_));
 sky130_fd_sc_hd__nand2_2 _36318_ (.A(_08730_),
    .B(_11433_),
    .Y(_14667_));
 sky130_fd_sc_hd__nand2_2 _36319_ (.A(_10415_),
    .B(_19167_),
    .Y(_14668_));
 sky130_fd_sc_hd__xor2_2 _36320_ (.A(_14667_),
    .B(_14668_),
    .X(_14669_));
 sky130_fd_sc_hd__a21o_2 _36321_ (.A1(_08086_),
    .A2(_14666_),
    .B1(_14669_),
    .X(_14670_));
 sky130_fd_sc_hd__and2_2 _36322_ (.A(_07846_),
    .B(_09809_),
    .X(_14671_));
 sky130_fd_sc_hd__nand2_2 _36323_ (.A(_14669_),
    .B(_14671_),
    .Y(_14672_));
 sky130_fd_sc_hd__o21ai_2 _36324_ (.A1(_14461_),
    .A2(_14462_),
    .B1(_14465_),
    .Y(_14673_));
 sky130_fd_sc_hd__a21o_2 _36325_ (.A1(_14670_),
    .A2(_14672_),
    .B1(_14673_),
    .X(_14674_));
 sky130_fd_sc_hd__nand3_2 _36326_ (.A(_14673_),
    .B(_14670_),
    .C(_14672_),
    .Y(_14675_));
 sky130_fd_sc_hd__and2_2 _36327_ (.A(_07162_),
    .B(_10895_),
    .X(_14676_));
 sky130_fd_sc_hd__a22oi_2 _36328_ (.A1(_18766_),
    .A2(_13580_),
    .B1(_18772_),
    .B2(_13113_),
    .Y(_14677_));
 sky130_fd_sc_hd__and4_2 _36329_ (.A(_10429_),
    .B(_12806_),
    .C(_13830_),
    .D(_11788_),
    .X(_14678_));
 sky130_fd_sc_hd__nor2_2 _36330_ (.A(_14677_),
    .B(_14678_),
    .Y(_14679_));
 sky130_fd_sc_hd__xor2_2 _36331_ (.A(_14676_),
    .B(_14679_),
    .X(_14680_));
 sky130_fd_sc_hd__a21oi_2 _36332_ (.A1(_14674_),
    .A2(_14675_),
    .B1(_14680_),
    .Y(_14681_));
 sky130_fd_sc_hd__nand3_2 _36333_ (.A(_14674_),
    .B(_14680_),
    .C(_14675_),
    .Y(_14682_));
 sky130_vsdinv _36334_ (.A(_14682_),
    .Y(_14683_));
 sky130_fd_sc_hd__nand2_2 _36335_ (.A(_14448_),
    .B(_14445_),
    .Y(_14684_));
 sky130_fd_sc_hd__o21bai_2 _36336_ (.A1(_14681_),
    .A2(_14683_),
    .B1_N(_14684_),
    .Y(_14685_));
 sky130_fd_sc_hd__nand3b_2 _36337_ (.A_N(_14681_),
    .B(_14684_),
    .C(_14682_),
    .Y(_14686_));
 sky130_fd_sc_hd__a21boi_2 _36338_ (.A1(_14470_),
    .A2(_14477_),
    .B1_N(_14471_),
    .Y(_14687_));
 sky130_vsdinv _36339_ (.A(_14687_),
    .Y(_14688_));
 sky130_fd_sc_hd__nand3_2 _36340_ (.A(_14685_),
    .B(_14686_),
    .C(_14688_),
    .Y(_14689_));
 sky130_vsdinv _36341_ (.A(_14689_),
    .Y(_14690_));
 sky130_fd_sc_hd__a21oi_2 _36342_ (.A1(_14685_),
    .A2(_14686_),
    .B1(_14688_),
    .Y(_14691_));
 sky130_fd_sc_hd__nand2_2 _36343_ (.A(_10487_),
    .B(_08255_),
    .Y(_14692_));
 sky130_fd_sc_hd__nand3b_2 _36344_ (.A_N(_14692_),
    .B(_10673_),
    .C(_19227_),
    .Y(_14693_));
 sky130_fd_sc_hd__o21ai_2 _36345_ (.A1(_06746_),
    .A2(_11332_),
    .B1(_14692_),
    .Y(_14694_));
 sky130_fd_sc_hd__and2_2 _36346_ (.A(_10268_),
    .B(_07606_),
    .X(_14695_));
 sky130_fd_sc_hd__a21o_2 _36347_ (.A1(_14693_),
    .A2(_14694_),
    .B1(_14695_),
    .X(_14696_));
 sky130_fd_sc_hd__nand3_2 _36348_ (.A(_14693_),
    .B(_14694_),
    .C(_14695_),
    .Y(_14697_));
 sky130_fd_sc_hd__nand2_2 _36349_ (.A(_14416_),
    .B(_14412_),
    .Y(_14698_));
 sky130_fd_sc_hd__a21o_2 _36350_ (.A1(_14696_),
    .A2(_14697_),
    .B1(_14698_),
    .X(_14699_));
 sky130_fd_sc_hd__nand3_2 _36351_ (.A(_14698_),
    .B(_14696_),
    .C(_14697_),
    .Y(_14700_));
 sky130_fd_sc_hd__buf_1 _36352_ (.A(_09320_),
    .X(_14701_));
 sky130_fd_sc_hd__nand2_2 _36353_ (.A(_14701_),
    .B(_13997_),
    .Y(_14702_));
 sky130_fd_sc_hd__nand2_2 _36354_ (.A(_18711_),
    .B(_10376_),
    .Y(_14703_));
 sky130_fd_sc_hd__nand2_2 _36355_ (.A(_10687_),
    .B(_10383_),
    .Y(_14704_));
 sky130_fd_sc_hd__xnor2_2 _36356_ (.A(_14703_),
    .B(_14704_),
    .Y(_14705_));
 sky130_fd_sc_hd__xor2_2 _36357_ (.A(_14702_),
    .B(_14705_),
    .X(_14706_));
 sky130_fd_sc_hd__a21oi_2 _36358_ (.A1(_14699_),
    .A2(_14700_),
    .B1(_14706_),
    .Y(_14707_));
 sky130_fd_sc_hd__nand3_2 _36359_ (.A(_14699_),
    .B(_14706_),
    .C(_14700_),
    .Y(_14708_));
 sky130_vsdinv _36360_ (.A(_14708_),
    .Y(_14709_));
 sky130_fd_sc_hd__a21oi_2 _36361_ (.A1(_14415_),
    .A2(_14416_),
    .B1(_14417_),
    .Y(_14710_));
 sky130_fd_sc_hd__xor2_2 _36362_ (.A(_14421_),
    .B(_14424_),
    .X(_14711_));
 sky130_fd_sc_hd__o21ai_2 _36363_ (.A1(_14710_),
    .A2(_14711_),
    .B1(_14419_),
    .Y(_14712_));
 sky130_fd_sc_hd__o21bai_2 _36364_ (.A1(_14707_),
    .A2(_14709_),
    .B1_N(_14712_),
    .Y(_14713_));
 sky130_fd_sc_hd__nand3b_2 _36365_ (.A_N(_14707_),
    .B(_14708_),
    .C(_14712_),
    .Y(_14714_));
 sky130_fd_sc_hd__nand2_2 _36366_ (.A(_14713_),
    .B(_14714_),
    .Y(_14715_));
 sky130_fd_sc_hd__buf_1 _36367_ (.A(_18736_),
    .X(_14716_));
 sky130_fd_sc_hd__nand3b_2 _36368_ (.A_N(_14435_),
    .B(_14716_),
    .C(_13787_),
    .Y(_14717_));
 sky130_fd_sc_hd__o31a_2 _36369_ (.A1(_18742_),
    .A2(_19188_),
    .A3(_14439_),
    .B1(_14717_),
    .X(_14718_));
 sky130_vsdinv _36370_ (.A(_14718_),
    .Y(_14719_));
 sky130_fd_sc_hd__nand2_2 _36371_ (.A(_12500_),
    .B(_09078_),
    .Y(_14720_));
 sky130_fd_sc_hd__nand2_2 _36372_ (.A(_08756_),
    .B(_09079_),
    .Y(_14721_));
 sky130_fd_sc_hd__xor2_2 _36373_ (.A(_14720_),
    .B(_14721_),
    .X(_14722_));
 sky130_fd_sc_hd__nand3_2 _36374_ (.A(_14722_),
    .B(_08459_),
    .C(_12329_),
    .Y(_14723_));
 sky130_fd_sc_hd__xnor2_2 _36375_ (.A(_14720_),
    .B(_14721_),
    .Y(_14724_));
 sky130_fd_sc_hd__o21ai_2 _36376_ (.A1(_18742_),
    .A2(_19182_),
    .B1(_14724_),
    .Y(_14725_));
 sky130_fd_sc_hd__nand2_2 _36377_ (.A(_14422_),
    .B(_14423_),
    .Y(_14726_));
 sky130_fd_sc_hd__nor2_2 _36378_ (.A(_14422_),
    .B(_14423_),
    .Y(_14727_));
 sky130_fd_sc_hd__a21oi_2 _36379_ (.A1(_14726_),
    .A2(_14421_),
    .B1(_14727_),
    .Y(_14728_));
 sky130_vsdinv _36380_ (.A(_14728_),
    .Y(_14729_));
 sky130_fd_sc_hd__a21o_2 _36381_ (.A1(_14723_),
    .A2(_14725_),
    .B1(_14729_),
    .X(_14730_));
 sky130_fd_sc_hd__nand3_2 _36382_ (.A(_14723_),
    .B(_14725_),
    .C(_14729_),
    .Y(_14731_));
 sky130_fd_sc_hd__nand2_2 _36383_ (.A(_14730_),
    .B(_14731_),
    .Y(_14732_));
 sky130_fd_sc_hd__xor2_2 _36384_ (.A(_14719_),
    .B(_14732_),
    .X(_14733_));
 sky130_fd_sc_hd__nand2_2 _36385_ (.A(_14715_),
    .B(_14733_),
    .Y(_14734_));
 sky130_fd_sc_hd__xor2_2 _36386_ (.A(_14718_),
    .B(_14732_),
    .X(_14735_));
 sky130_fd_sc_hd__nand3_2 _36387_ (.A(_14735_),
    .B(_14714_),
    .C(_14713_),
    .Y(_14736_));
 sky130_fd_sc_hd__o21ai_2 _36388_ (.A1(_14450_),
    .A2(_14452_),
    .B1(_14434_),
    .Y(_14737_));
 sky130_fd_sc_hd__a21oi_2 _36389_ (.A1(_14734_),
    .A2(_14736_),
    .B1(_14737_),
    .Y(_14738_));
 sky130_fd_sc_hd__nand3_2 _36390_ (.A(_14734_),
    .B(_14736_),
    .C(_14737_),
    .Y(_14739_));
 sky130_vsdinv _36391_ (.A(_14739_),
    .Y(_14740_));
 sky130_fd_sc_hd__o22ai_2 _36392_ (.A1(_14690_),
    .A2(_14691_),
    .B1(_14738_),
    .B2(_14740_),
    .Y(_14741_));
 sky130_fd_sc_hd__nor2_2 _36393_ (.A(_14691_),
    .B(_14690_),
    .Y(_14742_));
 sky130_fd_sc_hd__a21o_2 _36394_ (.A1(_14734_),
    .A2(_14736_),
    .B1(_14737_),
    .X(_14743_));
 sky130_fd_sc_hd__nand3_2 _36395_ (.A(_14742_),
    .B(_14739_),
    .C(_14743_),
    .Y(_14744_));
 sky130_fd_sc_hd__nand2_2 _36396_ (.A(_14741_),
    .B(_14744_),
    .Y(_14745_));
 sky130_fd_sc_hd__o21ai_2 _36397_ (.A1(_14494_),
    .A2(_14495_),
    .B1(_14459_),
    .Y(_14746_));
 sky130_vsdinv _36398_ (.A(_14746_),
    .Y(_14747_));
 sky130_fd_sc_hd__nand2_2 _36399_ (.A(_14745_),
    .B(_14747_),
    .Y(_14748_));
 sky130_fd_sc_hd__nand3_2 _36400_ (.A(_14741_),
    .B(_14744_),
    .C(_14746_),
    .Y(_14749_));
 sky130_fd_sc_hd__a22oi_2 _36401_ (.A1(_14664_),
    .A2(_14665_),
    .B1(_14748_),
    .B2(_14749_),
    .Y(_14750_));
 sky130_fd_sc_hd__nand2_2 _36402_ (.A(_14665_),
    .B(_14664_),
    .Y(_14751_));
 sky130_fd_sc_hd__nand2_2 _36403_ (.A(_14748_),
    .B(_14749_),
    .Y(_14752_));
 sky130_fd_sc_hd__nor2_2 _36404_ (.A(_14751_),
    .B(_14752_),
    .Y(_14753_));
 sky130_fd_sc_hd__o21ai_2 _36405_ (.A1(_14552_),
    .A2(_14553_),
    .B1(_14503_),
    .Y(_14754_));
 sky130_fd_sc_hd__o21bai_2 _36406_ (.A1(_14750_),
    .A2(_14753_),
    .B1_N(_14754_),
    .Y(_14755_));
 sky130_fd_sc_hd__nand2_2 _36407_ (.A(_14752_),
    .B(_14751_),
    .Y(_14756_));
 sky130_fd_sc_hd__a21oi_2 _36408_ (.A1(_14659_),
    .A2(_14663_),
    .B1(_14662_),
    .Y(_14757_));
 sky130_vsdinv _36409_ (.A(_14664_),
    .Y(_14758_));
 sky130_fd_sc_hd__nor2_2 _36410_ (.A(_14757_),
    .B(_14758_),
    .Y(_14759_));
 sky130_fd_sc_hd__nand3_2 _36411_ (.A(_14759_),
    .B(_14748_),
    .C(_14749_),
    .Y(_14760_));
 sky130_fd_sc_hd__nand3_2 _36412_ (.A(_14756_),
    .B(_14760_),
    .C(_14754_),
    .Y(_14761_));
 sky130_fd_sc_hd__o21ai_2 _36413_ (.A1(_14649_),
    .A2(_14532_),
    .B1(_14127_),
    .Y(_14762_));
 sky130_vsdinv _36414_ (.A(_14649_),
    .Y(_14763_));
 sky130_fd_sc_hd__nand2_2 _36415_ (.A(_14529_),
    .B(_14530_),
    .Y(_14764_));
 sky130_fd_sc_hd__nand2_2 _36416_ (.A(_14764_),
    .B(_14316_),
    .Y(_14765_));
 sky130_fd_sc_hd__o211ai_2 _36417_ (.A1(_14125_),
    .A2(_14126_),
    .B1(_14763_),
    .C1(_14765_),
    .Y(_14766_));
 sky130_fd_sc_hd__a21oi_2 _36418_ (.A1(_14762_),
    .A2(_14766_),
    .B1(_14354_),
    .Y(_14767_));
 sky130_fd_sc_hd__a21boi_2 _36419_ (.A1(_14563_),
    .A2(_14354_),
    .B1_N(_14565_),
    .Y(_14768_));
 sky130_vsdinv _36420_ (.A(_14768_),
    .Y(_14769_));
 sky130_fd_sc_hd__nand3_2 _36421_ (.A(_14762_),
    .B(_14766_),
    .C(_14351_),
    .Y(_14770_));
 sky130_fd_sc_hd__nand3b_2 _36422_ (.A_N(_14767_),
    .B(_14769_),
    .C(_14770_),
    .Y(_14771_));
 sky130_vsdinv _36423_ (.A(_14770_),
    .Y(_14772_));
 sky130_fd_sc_hd__o21ai_2 _36424_ (.A1(_14767_),
    .A2(_14772_),
    .B1(_14768_),
    .Y(_14773_));
 sky130_fd_sc_hd__a21oi_2 _36425_ (.A1(_14771_),
    .A2(_14773_),
    .B1(_13193_),
    .Y(_14774_));
 sky130_fd_sc_hd__and3_2 _36426_ (.A(_14771_),
    .B(_14773_),
    .C(_12944_),
    .X(_14775_));
 sky130_vsdinv _36427_ (.A(_14775_),
    .Y(_14776_));
 sky130_fd_sc_hd__o21ai_2 _36428_ (.A1(_14542_),
    .A2(_14549_),
    .B1(_14541_),
    .Y(_14777_));
 sky130_fd_sc_hd__nand3b_2 _36429_ (.A_N(_14774_),
    .B(_14776_),
    .C(_14777_),
    .Y(_14778_));
 sky130_fd_sc_hd__buf_1 _36430_ (.A(_14778_),
    .X(_14779_));
 sky130_fd_sc_hd__o21bai_2 _36431_ (.A1(_14774_),
    .A2(_14775_),
    .B1_N(_14777_),
    .Y(_14780_));
 sky130_fd_sc_hd__a21boi_2 _36432_ (.A1(_14570_),
    .A2(_13440_),
    .B1_N(_14571_),
    .Y(_14781_));
 sky130_vsdinv _36433_ (.A(_14781_),
    .Y(_14782_));
 sky130_fd_sc_hd__a21oi_2 _36434_ (.A1(_14779_),
    .A2(_14780_),
    .B1(_14782_),
    .Y(_14783_));
 sky130_fd_sc_hd__nand3_2 _36435_ (.A(_14778_),
    .B(_14782_),
    .C(_14780_),
    .Y(_14784_));
 sky130_vsdinv _36436_ (.A(_14784_),
    .Y(_14785_));
 sky130_fd_sc_hd__nor2_2 _36437_ (.A(_14783_),
    .B(_14785_),
    .Y(_14786_));
 sky130_fd_sc_hd__a21oi_2 _36438_ (.A1(_14755_),
    .A2(_14761_),
    .B1(_14786_),
    .Y(_14787_));
 sky130_fd_sc_hd__nand2_2 _36439_ (.A(_14779_),
    .B(_14780_),
    .Y(_14788_));
 sky130_fd_sc_hd__nand2_2 _36440_ (.A(_14788_),
    .B(_14781_),
    .Y(_14789_));
 sky130_fd_sc_hd__nand2_2 _36441_ (.A(_14789_),
    .B(_14784_),
    .Y(_14790_));
 sky130_fd_sc_hd__a21oi_2 _36442_ (.A1(_14756_),
    .A2(_14760_),
    .B1(_14754_),
    .Y(_14791_));
 sky130_vsdinv _36443_ (.A(_14761_),
    .Y(_14792_));
 sky130_fd_sc_hd__nor3_2 _36444_ (.A(_14790_),
    .B(_14791_),
    .C(_14792_),
    .Y(_14793_));
 sky130_fd_sc_hd__o21ai_2 _36445_ (.A1(_14587_),
    .A2(_14588_),
    .B1(_14562_),
    .Y(_14794_));
 sky130_fd_sc_hd__o21bai_2 _36446_ (.A1(_14787_),
    .A2(_14793_),
    .B1_N(_14794_),
    .Y(_14795_));
 sky130_fd_sc_hd__o22ai_2 _36447_ (.A1(_14785_),
    .A2(_14783_),
    .B1(_14791_),
    .B2(_14792_),
    .Y(_14796_));
 sky130_fd_sc_hd__nand3_2 _36448_ (.A(_14786_),
    .B(_14755_),
    .C(_14761_),
    .Y(_14797_));
 sky130_fd_sc_hd__nand3_2 _36449_ (.A(_14796_),
    .B(_14797_),
    .C(_14794_),
    .Y(_14798_));
 sky130_fd_sc_hd__buf_1 _36450_ (.A(_14798_),
    .X(_14799_));
 sky130_fd_sc_hd__nand2_2 _36451_ (.A(_14581_),
    .B(_14577_),
    .Y(_14800_));
 sky130_fd_sc_hd__xor2_2 _36452_ (.A(_13693_),
    .B(_14800_),
    .X(_14801_));
 sky130_fd_sc_hd__a21oi_2 _36453_ (.A1(_14795_),
    .A2(_14799_),
    .B1(_14801_),
    .Y(_14802_));
 sky130_vsdinv _36454_ (.A(_14801_),
    .Y(_14803_));
 sky130_fd_sc_hd__a21oi_2 _36455_ (.A1(_14796_),
    .A2(_14797_),
    .B1(_14794_),
    .Y(_14804_));
 sky130_fd_sc_hd__nor3b_2 _36456_ (.A(_14803_),
    .B(_14804_),
    .C_N(_14799_),
    .Y(_14805_));
 sky130_fd_sc_hd__o21ai_2 _36457_ (.A1(_14601_),
    .A2(_14602_),
    .B1(_14597_),
    .Y(_14806_));
 sky130_fd_sc_hd__o21bai_2 _36458_ (.A1(_14802_),
    .A2(_14805_),
    .B1_N(_14806_),
    .Y(_14807_));
 sky130_fd_sc_hd__nand2_2 _36459_ (.A(_14795_),
    .B(_14798_),
    .Y(_14808_));
 sky130_fd_sc_hd__nand2_2 _36460_ (.A(_14808_),
    .B(_14803_),
    .Y(_14809_));
 sky130_fd_sc_hd__nand3_2 _36461_ (.A(_14795_),
    .B(_14801_),
    .C(_14799_),
    .Y(_14810_));
 sky130_fd_sc_hd__nand3_2 _36462_ (.A(_14809_),
    .B(_14810_),
    .C(_14806_),
    .Y(_14811_));
 sky130_fd_sc_hd__buf_1 _36463_ (.A(_13468_),
    .X(_14812_));
 sky130_fd_sc_hd__a21oi_2 _36464_ (.A1(_14371_),
    .A2(_14367_),
    .B1(_14812_),
    .Y(_14813_));
 sky130_fd_sc_hd__a21oi_2 _36465_ (.A1(_14807_),
    .A2(_14811_),
    .B1(_14813_),
    .Y(_14814_));
 sky130_vsdinv _36466_ (.A(_14813_),
    .Y(_14815_));
 sky130_fd_sc_hd__a21oi_2 _36467_ (.A1(_14809_),
    .A2(_14810_),
    .B1(_14806_),
    .Y(_14816_));
 sky130_vsdinv _36468_ (.A(_14811_),
    .Y(_14817_));
 sky130_fd_sc_hd__nor3_2 _36469_ (.A(_14815_),
    .B(_14816_),
    .C(_14817_),
    .Y(_14818_));
 sky130_fd_sc_hd__o21ai_2 _36470_ (.A1(_14613_),
    .A2(_14614_),
    .B1(_14610_),
    .Y(_14819_));
 sky130_fd_sc_hd__o21bai_2 _36471_ (.A1(_14814_),
    .A2(_14818_),
    .B1_N(_14819_),
    .Y(_14820_));
 sky130_fd_sc_hd__o21bai_2 _36472_ (.A1(_14816_),
    .A2(_14817_),
    .B1_N(_14813_),
    .Y(_14821_));
 sky130_fd_sc_hd__nand3_2 _36473_ (.A(_14807_),
    .B(_14813_),
    .C(_14811_),
    .Y(_14822_));
 sky130_fd_sc_hd__nand3_2 _36474_ (.A(_14821_),
    .B(_14819_),
    .C(_14822_),
    .Y(_14823_));
 sky130_fd_sc_hd__and2_2 _36475_ (.A(_14820_),
    .B(_14823_),
    .X(_14824_));
 sky130_fd_sc_hd__o21ai_2 _36476_ (.A1(_14623_),
    .A2(_14628_),
    .B1(_14622_),
    .Y(_14825_));
 sky130_fd_sc_hd__xor2_2 _36477_ (.A(_14824_),
    .B(_14825_),
    .X(_02666_));
 sky130_fd_sc_hd__nand2_2 _36478_ (.A(_08011_),
    .B(_12097_),
    .Y(_14826_));
 sky130_fd_sc_hd__nand2_2 _36479_ (.A(_12099_),
    .B(_07474_),
    .Y(_14827_));
 sky130_fd_sc_hd__xor2_2 _36480_ (.A(_14826_),
    .B(_14827_),
    .X(_14828_));
 sky130_fd_sc_hd__nand2_2 _36481_ (.A(_14828_),
    .B(_14633_),
    .Y(_14829_));
 sky130_fd_sc_hd__buf_1 _36482_ (.A(_14522_),
    .X(_14830_));
 sky130_fd_sc_hd__buf_1 _36483_ (.A(_14830_),
    .X(_14831_));
 sky130_fd_sc_hd__a21o_2 _36484_ (.A1(_14831_),
    .A2(_06668_),
    .B1(_14828_),
    .X(_14832_));
 sky130_fd_sc_hd__a21oi_2 _36485_ (.A1(_14679_),
    .A2(_14676_),
    .B1(_14678_),
    .Y(_14833_));
 sky130_fd_sc_hd__a21bo_2 _36486_ (.A1(_14829_),
    .A2(_14832_),
    .B1_N(_14833_),
    .X(_14834_));
 sky130_fd_sc_hd__nand3b_2 _36487_ (.A_N(_14833_),
    .B(_14829_),
    .C(_14832_),
    .Y(_14835_));
 sky130_fd_sc_hd__o21a_2 _36488_ (.A1(_14629_),
    .A2(_14630_),
    .B1(_14637_),
    .X(_14836_));
 sky130_vsdinv _36489_ (.A(_14836_),
    .Y(_14837_));
 sky130_fd_sc_hd__a21o_2 _36490_ (.A1(_14834_),
    .A2(_14835_),
    .B1(_14837_),
    .X(_14838_));
 sky130_fd_sc_hd__nand3_2 _36491_ (.A(_14834_),
    .B(_14835_),
    .C(_14837_),
    .Y(_14839_));
 sky130_fd_sc_hd__nand2_2 _36492_ (.A(_14643_),
    .B(_14640_),
    .Y(_14840_));
 sky130_fd_sc_hd__a21o_2 _36493_ (.A1(_14838_),
    .A2(_14839_),
    .B1(_14840_),
    .X(_14841_));
 sky130_fd_sc_hd__nand3_2 _36494_ (.A(_14838_),
    .B(_14839_),
    .C(_14840_),
    .Y(_14842_));
 sky130_fd_sc_hd__buf_1 _36495_ (.A(_14655_),
    .X(_14843_));
 sky130_fd_sc_hd__a21o_2 _36496_ (.A1(_14841_),
    .A2(_14842_),
    .B1(_14843_),
    .X(_14844_));
 sky130_fd_sc_hd__nand3_2 _36497_ (.A(_14841_),
    .B(_14843_),
    .C(_14842_),
    .Y(_14845_));
 sky130_fd_sc_hd__nand2_2 _36498_ (.A(_14689_),
    .B(_14686_),
    .Y(_14846_));
 sky130_fd_sc_hd__a21o_2 _36499_ (.A1(_14844_),
    .A2(_14845_),
    .B1(_14846_),
    .X(_14847_));
 sky130_fd_sc_hd__nand3_2 _36500_ (.A(_14844_),
    .B(_14846_),
    .C(_14845_),
    .Y(_14848_));
 sky130_fd_sc_hd__buf_1 _36501_ (.A(_14656_),
    .X(_14849_));
 sky130_fd_sc_hd__a21boi_2 _36502_ (.A1(_14645_),
    .A2(_14849_),
    .B1_N(_14646_),
    .Y(_14850_));
 sky130_fd_sc_hd__a21bo_2 _36503_ (.A1(_14847_),
    .A2(_14848_),
    .B1_N(_14850_),
    .X(_14851_));
 sky130_fd_sc_hd__nand3b_2 _36504_ (.A_N(_14850_),
    .B(_14847_),
    .C(_14848_),
    .Y(_14852_));
 sky130_fd_sc_hd__nand2_2 _36505_ (.A(_14851_),
    .B(_14852_),
    .Y(_14853_));
 sky130_fd_sc_hd__nand3b_2 _36506_ (.A_N(_14703_),
    .B(_18719_),
    .C(_08304_),
    .Y(_14854_));
 sky130_fd_sc_hd__nand3b_2 _36507_ (.A_N(_14705_),
    .B(_14701_),
    .C(_13997_),
    .Y(_14855_));
 sky130_fd_sc_hd__and2_2 _36508_ (.A(_08458_),
    .B(_09785_),
    .X(_14856_));
 sky130_fd_sc_hd__buf_1 _36509_ (.A(_09006_),
    .X(_14857_));
 sky130_fd_sc_hd__nand2_2 _36510_ (.A(_14857_),
    .B(_10070_),
    .Y(_14858_));
 sky130_fd_sc_hd__nand2_2 _36511_ (.A(_18735_),
    .B(_09089_),
    .Y(_14859_));
 sky130_fd_sc_hd__xnor2_2 _36512_ (.A(_14858_),
    .B(_14859_),
    .Y(_14860_));
 sky130_fd_sc_hd__xor2_2 _36513_ (.A(_14856_),
    .B(_14860_),
    .X(_14861_));
 sky130_fd_sc_hd__a21o_2 _36514_ (.A1(_14854_),
    .A2(_14855_),
    .B1(_14861_),
    .X(_14862_));
 sky130_fd_sc_hd__buf_1 _36515_ (.A(_11036_),
    .X(_14863_));
 sky130_fd_sc_hd__nand3b_2 _36516_ (.A_N(_14720_),
    .B(_14716_),
    .C(_09105_),
    .Y(_14864_));
 sky130_fd_sc_hd__o31a_2 _36517_ (.A1(_14863_),
    .A2(_19182_),
    .A3(_14724_),
    .B1(_14864_),
    .X(_14865_));
 sky130_vsdinv _36518_ (.A(_14865_),
    .Y(_14866_));
 sky130_fd_sc_hd__nand3_2 _36519_ (.A(_14861_),
    .B(_14854_),
    .C(_14855_),
    .Y(_14867_));
 sky130_fd_sc_hd__nand3_2 _36520_ (.A(_14862_),
    .B(_14866_),
    .C(_14867_),
    .Y(_14868_));
 sky130_fd_sc_hd__a21o_2 _36521_ (.A1(_14862_),
    .A2(_14867_),
    .B1(_14866_),
    .X(_14869_));
 sky130_fd_sc_hd__and2_2 _36522_ (.A(_10268_),
    .B(_08300_),
    .X(_14870_));
 sky130_fd_sc_hd__buf_1 _36523_ (.A(_10994_),
    .X(_14871_));
 sky130_fd_sc_hd__a22oi_2 _36524_ (.A1(_14871_),
    .A2(_06937_),
    .B1(_19217_),
    .B2(_11322_),
    .Y(_14872_));
 sky130_fd_sc_hd__nand2_2 _36525_ (.A(_18695_),
    .B(_07737_),
    .Y(_14873_));
 sky130_fd_sc_hd__nor3_2 _36526_ (.A(_07329_),
    .B(_11005_),
    .C(_14873_),
    .Y(_14874_));
 sky130_fd_sc_hd__nor2_2 _36527_ (.A(_14872_),
    .B(_14874_),
    .Y(_14875_));
 sky130_fd_sc_hd__xnor2_2 _36528_ (.A(_14870_),
    .B(_14875_),
    .Y(_14876_));
 sky130_fd_sc_hd__a21boi_2 _36529_ (.A1(_14694_),
    .A2(_14695_),
    .B1_N(_14693_),
    .Y(_14877_));
 sky130_fd_sc_hd__nand2_2 _36530_ (.A(_14876_),
    .B(_14877_),
    .Y(_14878_));
 sky130_fd_sc_hd__o21bai_2 _36531_ (.A1(_14872_),
    .A2(_14874_),
    .B1_N(_14870_),
    .Y(_14879_));
 sky130_vsdinv _36532_ (.A(_14872_),
    .Y(_14880_));
 sky130_fd_sc_hd__nand3b_2 _36533_ (.A_N(_14874_),
    .B(_14880_),
    .C(_14870_),
    .Y(_14881_));
 sky130_fd_sc_hd__nand3b_2 _36534_ (.A_N(_14877_),
    .B(_14879_),
    .C(_14881_),
    .Y(_14882_));
 sky130_fd_sc_hd__and2_2 _36535_ (.A(_09321_),
    .B(_12292_),
    .X(_14883_));
 sky130_fd_sc_hd__buf_1 _36536_ (.A(_11338_),
    .X(_14884_));
 sky130_fd_sc_hd__a22oi_2 _36537_ (.A1(_14884_),
    .A2(_11714_),
    .B1(_18718_),
    .B2(_12288_),
    .Y(_14885_));
 sky130_fd_sc_hd__and4_2 _36538_ (.A(_10261_),
    .B(_10687_),
    .C(_08553_),
    .D(_10383_),
    .X(_14886_));
 sky130_fd_sc_hd__nor2_2 _36539_ (.A(_14885_),
    .B(_14886_),
    .Y(_14887_));
 sky130_fd_sc_hd__xor2_2 _36540_ (.A(_14883_),
    .B(_14887_),
    .X(_14888_));
 sky130_fd_sc_hd__a21oi_2 _36541_ (.A1(_14878_),
    .A2(_14882_),
    .B1(_14888_),
    .Y(_14889_));
 sky130_fd_sc_hd__nand3_2 _36542_ (.A(_14878_),
    .B(_14882_),
    .C(_14888_),
    .Y(_14890_));
 sky130_vsdinv _36543_ (.A(_14890_),
    .Y(_14891_));
 sky130_fd_sc_hd__nand2_2 _36544_ (.A(_14708_),
    .B(_14700_),
    .Y(_14892_));
 sky130_fd_sc_hd__o21bai_2 _36545_ (.A1(_14889_),
    .A2(_14891_),
    .B1_N(_14892_),
    .Y(_14893_));
 sky130_fd_sc_hd__nand3b_2 _36546_ (.A_N(_14889_),
    .B(_14890_),
    .C(_14892_),
    .Y(_14894_));
 sky130_fd_sc_hd__a22o_2 _36547_ (.A1(_14868_),
    .A2(_14869_),
    .B1(_14893_),
    .B2(_14894_),
    .X(_14895_));
 sky130_fd_sc_hd__nand2_2 _36548_ (.A(_14869_),
    .B(_14868_),
    .Y(_14896_));
 sky130_fd_sc_hd__nand3b_2 _36549_ (.A_N(_14896_),
    .B(_14893_),
    .C(_14894_),
    .Y(_14897_));
 sky130_fd_sc_hd__nand2_2 _36550_ (.A(_14736_),
    .B(_14714_),
    .Y(_14898_));
 sky130_fd_sc_hd__a21oi_2 _36551_ (.A1(_14895_),
    .A2(_14897_),
    .B1(_14898_),
    .Y(_14899_));
 sky130_fd_sc_hd__nand3_2 _36552_ (.A(_14895_),
    .B(_14897_),
    .C(_14898_),
    .Y(_14900_));
 sky130_vsdinv _36553_ (.A(_14900_),
    .Y(_14901_));
 sky130_fd_sc_hd__and2_2 _36554_ (.A(_12538_),
    .B(_11199_),
    .X(_14902_));
 sky130_fd_sc_hd__a22oi_2 _36555_ (.A1(_12805_),
    .A2(_12316_),
    .B1(_08220_),
    .B2(_12069_),
    .Y(_14903_));
 sky130_fd_sc_hd__and4_2 _36556_ (.A(_18765_),
    .B(_12254_),
    .C(_11791_),
    .D(_09805_),
    .X(_14904_));
 sky130_fd_sc_hd__nor2_2 _36557_ (.A(_14903_),
    .B(_14904_),
    .Y(_14905_));
 sky130_fd_sc_hd__xor2_2 _36558_ (.A(_14902_),
    .B(_14905_),
    .X(_14906_));
 sky130_vsdinv _36559_ (.A(_14906_),
    .Y(_14907_));
 sky130_fd_sc_hd__a22o_2 _36560_ (.A1(_14245_),
    .A2(_11224_),
    .B1(_11968_),
    .B2(_19162_),
    .X(_14908_));
 sky130_fd_sc_hd__nand2_2 _36561_ (.A(_08730_),
    .B(_09790_),
    .Y(_14909_));
 sky130_fd_sc_hd__nand3b_2 _36562_ (.A_N(_14909_),
    .B(_11074_),
    .C(_10849_),
    .Y(_14910_));
 sky130_fd_sc_hd__o2bb2ai_2 _36563_ (.A1_N(_14908_),
    .A2_N(_14910_),
    .B1(_13050_),
    .B2(_19158_),
    .Y(_14911_));
 sky130_fd_sc_hd__and2_2 _36564_ (.A(_12531_),
    .B(_12035_),
    .X(_14912_));
 sky130_fd_sc_hd__nand3_2 _36565_ (.A(_14910_),
    .B(_14908_),
    .C(_14912_),
    .Y(_14913_));
 sky130_fd_sc_hd__nand2_2 _36566_ (.A(_14911_),
    .B(_14913_),
    .Y(_14914_));
 sky130_fd_sc_hd__o21ai_2 _36567_ (.A1(_14667_),
    .A2(_14668_),
    .B1(_14672_),
    .Y(_14915_));
 sky130_fd_sc_hd__xor2_2 _36568_ (.A(_14914_),
    .B(_14915_),
    .X(_14916_));
 sky130_fd_sc_hd__nor2_2 _36569_ (.A(_14907_),
    .B(_14916_),
    .Y(_14917_));
 sky130_fd_sc_hd__and2_2 _36570_ (.A(_14916_),
    .B(_14907_),
    .X(_14918_));
 sky130_fd_sc_hd__a21boi_2 _36571_ (.A1(_14719_),
    .A2(_14730_),
    .B1_N(_14731_),
    .Y(_14919_));
 sky130_vsdinv _36572_ (.A(_14919_),
    .Y(_14920_));
 sky130_fd_sc_hd__o21bai_2 _36573_ (.A1(_14917_),
    .A2(_14918_),
    .B1_N(_14920_),
    .Y(_14921_));
 sky130_fd_sc_hd__nand2_2 _36574_ (.A(_14916_),
    .B(_14907_),
    .Y(_14922_));
 sky130_fd_sc_hd__nand3b_2 _36575_ (.A_N(_14917_),
    .B(_14920_),
    .C(_14922_),
    .Y(_14923_));
 sky130_fd_sc_hd__a21boi_2 _36576_ (.A1(_14674_),
    .A2(_14680_),
    .B1_N(_14675_),
    .Y(_14924_));
 sky130_fd_sc_hd__a21bo_2 _36577_ (.A1(_14921_),
    .A2(_14923_),
    .B1_N(_14924_),
    .X(_14925_));
 sky130_fd_sc_hd__nand3b_2 _36578_ (.A_N(_14924_),
    .B(_14921_),
    .C(_14923_),
    .Y(_14926_));
 sky130_fd_sc_hd__nand2_2 _36579_ (.A(_14925_),
    .B(_14926_),
    .Y(_14927_));
 sky130_fd_sc_hd__o21ai_2 _36580_ (.A1(_14899_),
    .A2(_14901_),
    .B1(_14927_),
    .Y(_14928_));
 sky130_fd_sc_hd__a21o_2 _36581_ (.A1(_14895_),
    .A2(_14897_),
    .B1(_14898_),
    .X(_14929_));
 sky130_fd_sc_hd__nand3b_2 _36582_ (.A_N(_14927_),
    .B(_14929_),
    .C(_14900_),
    .Y(_14930_));
 sky130_fd_sc_hd__o31ai_2 _36583_ (.A1(_14691_),
    .A2(_14690_),
    .A3(_14738_),
    .B1(_14739_),
    .Y(_14931_));
 sky130_fd_sc_hd__a21o_2 _36584_ (.A1(_14928_),
    .A2(_14930_),
    .B1(_14931_),
    .X(_14932_));
 sky130_fd_sc_hd__nand3_2 _36585_ (.A(_14928_),
    .B(_14930_),
    .C(_14931_),
    .Y(_14933_));
 sky130_fd_sc_hd__nand3b_2 _36586_ (.A_N(_14853_),
    .B(_14932_),
    .C(_14933_),
    .Y(_14934_));
 sky130_fd_sc_hd__a21oi_2 _36587_ (.A1(_14928_),
    .A2(_14930_),
    .B1(_14931_),
    .Y(_14935_));
 sky130_vsdinv _36588_ (.A(_14933_),
    .Y(_14936_));
 sky130_fd_sc_hd__o21ai_2 _36589_ (.A1(_14935_),
    .A2(_14936_),
    .B1(_14853_),
    .Y(_14937_));
 sky130_fd_sc_hd__o21ai_2 _36590_ (.A1(_14751_),
    .A2(_14752_),
    .B1(_14749_),
    .Y(_14938_));
 sky130_fd_sc_hd__a21oi_2 _36591_ (.A1(_14934_),
    .A2(_14937_),
    .B1(_14938_),
    .Y(_14939_));
 sky130_fd_sc_hd__nand3_2 _36592_ (.A(_14934_),
    .B(_14937_),
    .C(_14938_),
    .Y(_14940_));
 sky130_vsdinv _36593_ (.A(_14940_),
    .Y(_14941_));
 sky130_fd_sc_hd__a21oi_2 _36594_ (.A1(_14316_),
    .A2(_14650_),
    .B1(_14649_),
    .Y(_14942_));
 sky130_fd_sc_hd__or2b_2 _36595_ (.A(_14942_),
    .B_N(_14128_),
    .X(_14943_));
 sky130_fd_sc_hd__o21ai_2 _36596_ (.A1(_14347_),
    .A2(_14348_),
    .B1(_14942_),
    .Y(_14944_));
 sky130_fd_sc_hd__a21oi_2 _36597_ (.A1(_14943_),
    .A2(_14944_),
    .B1(_14352_),
    .Y(_14945_));
 sky130_fd_sc_hd__and3_2 _36598_ (.A(_14943_),
    .B(_14352_),
    .C(_14944_),
    .X(_14946_));
 sky130_fd_sc_hd__a211o_2 _36599_ (.A1(_14762_),
    .A2(_14770_),
    .B1(_14945_),
    .C1(_14946_),
    .X(_14947_));
 sky130_fd_sc_hd__o211ai_2 _36600_ (.A1(_14945_),
    .A2(_14946_),
    .B1(_14762_),
    .C1(_14770_),
    .Y(_14948_));
 sky130_fd_sc_hd__a21o_2 _36601_ (.A1(_14947_),
    .A2(_14948_),
    .B1(_13194_),
    .X(_14949_));
 sky130_fd_sc_hd__nand3_2 _36602_ (.A(_14947_),
    .B(_13194_),
    .C(_14948_),
    .Y(_14950_));
 sky130_fd_sc_hd__a21boi_2 _36603_ (.A1(_14659_),
    .A2(_14662_),
    .B1_N(_14663_),
    .Y(_14951_));
 sky130_fd_sc_hd__a21bo_2 _36604_ (.A1(_14949_),
    .A2(_14950_),
    .B1_N(_14951_),
    .X(_14952_));
 sky130_fd_sc_hd__nand3b_2 _36605_ (.A_N(_14951_),
    .B(_14949_),
    .C(_14950_),
    .Y(_14953_));
 sky130_fd_sc_hd__nand2_2 _36606_ (.A(_14952_),
    .B(_14953_),
    .Y(_14954_));
 sky130_fd_sc_hd__buf_1 _36607_ (.A(_14360_),
    .X(_14955_));
 sky130_fd_sc_hd__a21boi_2 _36608_ (.A1(_14955_),
    .A2(_14773_),
    .B1_N(_14771_),
    .Y(_14956_));
 sky130_fd_sc_hd__nand2_2 _36609_ (.A(_14954_),
    .B(_14956_),
    .Y(_14957_));
 sky130_fd_sc_hd__nand3b_2 _36610_ (.A_N(_14956_),
    .B(_14952_),
    .C(_14953_),
    .Y(_14958_));
 sky130_fd_sc_hd__nand2_2 _36611_ (.A(_14957_),
    .B(_14958_),
    .Y(_14959_));
 sky130_fd_sc_hd__o21ai_2 _36612_ (.A1(_14939_),
    .A2(_14941_),
    .B1(_14959_),
    .Y(_14960_));
 sky130_fd_sc_hd__a21o_2 _36613_ (.A1(_14934_),
    .A2(_14937_),
    .B1(_14938_),
    .X(_14961_));
 sky130_fd_sc_hd__nand3b_2 _36614_ (.A_N(_14959_),
    .B(_14961_),
    .C(_14940_),
    .Y(_14962_));
 sky130_fd_sc_hd__o21ai_2 _36615_ (.A1(_14790_),
    .A2(_14791_),
    .B1(_14761_),
    .Y(_14963_));
 sky130_fd_sc_hd__a21oi_2 _36616_ (.A1(_14960_),
    .A2(_14962_),
    .B1(_14963_),
    .Y(_14964_));
 sky130_fd_sc_hd__nand3_2 _36617_ (.A(_14960_),
    .B(_14962_),
    .C(_14963_),
    .Y(_14965_));
 sky130_vsdinv _36618_ (.A(_14965_),
    .Y(_14966_));
 sky130_fd_sc_hd__a21boi_2 _36619_ (.A1(_14782_),
    .A2(_14780_),
    .B1_N(_14779_),
    .Y(_14967_));
 sky130_fd_sc_hd__xor2_2 _36620_ (.A(_13456_),
    .B(_14967_),
    .X(_14968_));
 sky130_fd_sc_hd__o21bai_2 _36621_ (.A1(_14964_),
    .A2(_14966_),
    .B1_N(_14968_),
    .Y(_14969_));
 sky130_fd_sc_hd__a21o_2 _36622_ (.A1(_14960_),
    .A2(_14962_),
    .B1(_14963_),
    .X(_14970_));
 sky130_fd_sc_hd__nand3_2 _36623_ (.A(_14970_),
    .B(_14968_),
    .C(_14965_),
    .Y(_14971_));
 sky130_fd_sc_hd__o21ai_2 _36624_ (.A1(_14803_),
    .A2(_14804_),
    .B1(_14799_),
    .Y(_14972_));
 sky130_fd_sc_hd__a21oi_2 _36625_ (.A1(_14969_),
    .A2(_14971_),
    .B1(_14972_),
    .Y(_14973_));
 sky130_fd_sc_hd__and3_2 _36626_ (.A(_14969_),
    .B(_14971_),
    .C(_14972_),
    .X(_14974_));
 sky130_fd_sc_hd__buf_1 _36627_ (.A(_13468_),
    .X(_14975_));
 sky130_fd_sc_hd__buf_1 _36628_ (.A(_14975_),
    .X(_14976_));
 sky130_fd_sc_hd__a21oi_2 _36629_ (.A1(_14581_),
    .A2(_14577_),
    .B1(_14976_),
    .Y(_14977_));
 sky130_fd_sc_hd__o21bai_2 _36630_ (.A1(_14973_),
    .A2(_14974_),
    .B1_N(_14977_),
    .Y(_14978_));
 sky130_fd_sc_hd__a21o_2 _36631_ (.A1(_14969_),
    .A2(_14971_),
    .B1(_14972_),
    .X(_14979_));
 sky130_fd_sc_hd__nand3_2 _36632_ (.A(_14969_),
    .B(_14971_),
    .C(_14972_),
    .Y(_14980_));
 sky130_fd_sc_hd__nand3_2 _36633_ (.A(_14979_),
    .B(_14977_),
    .C(_14980_),
    .Y(_14981_));
 sky130_fd_sc_hd__o21ai_2 _36634_ (.A1(_14815_),
    .A2(_14816_),
    .B1(_14811_),
    .Y(_14982_));
 sky130_fd_sc_hd__a21oi_2 _36635_ (.A1(_14978_),
    .A2(_14981_),
    .B1(_14982_),
    .Y(_14983_));
 sky130_fd_sc_hd__nand3_2 _36636_ (.A(_14978_),
    .B(_14981_),
    .C(_14982_),
    .Y(_14984_));
 sky130_vsdinv _36637_ (.A(_14984_),
    .Y(_14985_));
 sky130_fd_sc_hd__nor2_2 _36638_ (.A(_14983_),
    .B(_14985_),
    .Y(_14986_));
 sky130_fd_sc_hd__nand2_2 _36639_ (.A(_14820_),
    .B(_14823_),
    .Y(_14987_));
 sky130_fd_sc_hd__nor2_2 _36640_ (.A(_14623_),
    .B(_14987_),
    .Y(_14988_));
 sky130_fd_sc_hd__nand2_2 _36641_ (.A(_14625_),
    .B(_14988_),
    .Y(_14989_));
 sky130_fd_sc_hd__nor2_2 _36642_ (.A(_14190_),
    .B(_14989_),
    .Y(_14990_));
 sky130_fd_sc_hd__nand3_2 _36643_ (.A(_10992_),
    .B(_13243_),
    .C(_14990_),
    .Y(_14991_));
 sky130_fd_sc_hd__o21ai_2 _36644_ (.A1(_13246_),
    .A2(_13244_),
    .B1(_14990_),
    .Y(_14992_));
 sky130_vsdinv _36645_ (.A(_14404_),
    .Y(_14993_));
 sky130_fd_sc_hd__nor2_2 _36646_ (.A(_14626_),
    .B(_14993_),
    .Y(_14994_));
 sky130_fd_sc_hd__nand2_2 _36647_ (.A(_14186_),
    .B(_14994_),
    .Y(_14995_));
 sky130_fd_sc_hd__and2_2 _36648_ (.A(_14619_),
    .B(_14622_),
    .X(_14996_));
 sky130_fd_sc_hd__nand2_2 _36649_ (.A(_14824_),
    .B(_14996_),
    .Y(_14997_));
 sky130_fd_sc_hd__nor2_2 _36650_ (.A(_14995_),
    .B(_14997_),
    .Y(_14998_));
 sky130_fd_sc_hd__nand3_2 _36651_ (.A(_14824_),
    .B(_14996_),
    .C(_14627_),
    .Y(_14999_));
 sky130_fd_sc_hd__or2b_2 _36652_ (.A(_14622_),
    .B_N(_14820_),
    .X(_15000_));
 sky130_fd_sc_hd__nand3_2 _36653_ (.A(_14999_),
    .B(_14823_),
    .C(_15000_),
    .Y(_15001_));
 sky130_fd_sc_hd__a21oi_2 _36654_ (.A1(_14998_),
    .A2(_14193_),
    .B1(_15001_),
    .Y(_15002_));
 sky130_fd_sc_hd__nand3_2 _36655_ (.A(_14991_),
    .B(_14992_),
    .C(_15002_),
    .Y(_15003_));
 sky130_fd_sc_hd__buf_1 _36656_ (.A(_15003_),
    .X(_15004_));
 sky130_fd_sc_hd__xor2_2 _36657_ (.A(_14986_),
    .B(_15004_),
    .X(_02667_));
 sky130_fd_sc_hd__and2_2 _36658_ (.A(_10268_),
    .B(_07967_),
    .X(_15005_));
 sky130_fd_sc_hd__a22oi_2 _36659_ (.A1(_10482_),
    .A2(_08300_),
    .B1(_19212_),
    .B2(_14411_),
    .Y(_15006_));
 sky130_fd_sc_hd__nand2_2 _36660_ (.A(_10482_),
    .B(_07942_),
    .Y(_15007_));
 sky130_fd_sc_hd__nor3_2 _36661_ (.A(_07948_),
    .B(_16970_),
    .C(_15007_),
    .Y(_15008_));
 sky130_fd_sc_hd__nor2_2 _36662_ (.A(_15006_),
    .B(_15008_),
    .Y(_15009_));
 sky130_fd_sc_hd__xnor2_2 _36663_ (.A(_15005_),
    .B(_15009_),
    .Y(_15010_));
 sky130_fd_sc_hd__a21oi_2 _36664_ (.A1(_14880_),
    .A2(_14870_),
    .B1(_14874_),
    .Y(_15011_));
 sky130_fd_sc_hd__nand2_2 _36665_ (.A(_15010_),
    .B(_15011_),
    .Y(_15012_));
 sky130_fd_sc_hd__o21bai_2 _36666_ (.A1(_15006_),
    .A2(_15008_),
    .B1_N(_15005_),
    .Y(_15013_));
 sky130_vsdinv _36667_ (.A(_15006_),
    .Y(_15014_));
 sky130_fd_sc_hd__nand3b_2 _36668_ (.A_N(_15008_),
    .B(_15014_),
    .C(_15005_),
    .Y(_15015_));
 sky130_fd_sc_hd__nand3b_2 _36669_ (.A_N(_15011_),
    .B(_15013_),
    .C(_15015_),
    .Y(_15016_));
 sky130_fd_sc_hd__buf_1 _36670_ (.A(_09320_),
    .X(_15017_));
 sky130_fd_sc_hd__and2_2 _36671_ (.A(_15017_),
    .B(_09105_),
    .X(_15018_));
 sky130_fd_sc_hd__buf_1 _36672_ (.A(_14884_),
    .X(_15019_));
 sky130_fd_sc_hd__buf_1 _36673_ (.A(_10262_),
    .X(_15020_));
 sky130_fd_sc_hd__buf_1 _36674_ (.A(_15020_),
    .X(_15021_));
 sky130_fd_sc_hd__a22oi_2 _36675_ (.A1(_15019_),
    .A2(_13997_),
    .B1(_15021_),
    .B2(_13787_),
    .Y(_15022_));
 sky130_fd_sc_hd__buf_1 _36676_ (.A(_10683_),
    .X(_15023_));
 sky130_fd_sc_hd__and4_2 _36677_ (.A(_15023_),
    .B(_18718_),
    .C(_11441_),
    .D(_12288_),
    .X(_15024_));
 sky130_fd_sc_hd__nor2_2 _36678_ (.A(_15022_),
    .B(_15024_),
    .Y(_15025_));
 sky130_fd_sc_hd__xor2_2 _36679_ (.A(_15018_),
    .B(_15025_),
    .X(_15026_));
 sky130_fd_sc_hd__a21o_2 _36680_ (.A1(_15012_),
    .A2(_15016_),
    .B1(_15026_),
    .X(_15027_));
 sky130_fd_sc_hd__nand3_2 _36681_ (.A(_15012_),
    .B(_15016_),
    .C(_15026_),
    .Y(_15028_));
 sky130_fd_sc_hd__nand2_2 _36682_ (.A(_14890_),
    .B(_14882_),
    .Y(_15029_));
 sky130_fd_sc_hd__a21oi_2 _36683_ (.A1(_15027_),
    .A2(_15028_),
    .B1(_15029_),
    .Y(_15030_));
 sky130_fd_sc_hd__nand3_2 _36684_ (.A(_15029_),
    .B(_15027_),
    .C(_15028_),
    .Y(_15031_));
 sky130_vsdinv _36685_ (.A(_15031_),
    .Y(_15032_));
 sky130_fd_sc_hd__and2_2 _36686_ (.A(_08458_),
    .B(_10844_),
    .X(_15033_));
 sky130_fd_sc_hd__nand2_2 _36687_ (.A(_14857_),
    .B(_08830_),
    .Y(_15034_));
 sky130_fd_sc_hd__nand2_2 _36688_ (.A(_18735_),
    .B(_12842_),
    .Y(_15035_));
 sky130_fd_sc_hd__xnor2_2 _36689_ (.A(_15034_),
    .B(_15035_),
    .Y(_15036_));
 sky130_fd_sc_hd__xor2_2 _36690_ (.A(_15033_),
    .B(_15036_),
    .X(_15037_));
 sky130_fd_sc_hd__a21o_2 _36691_ (.A1(_14887_),
    .A2(_14883_),
    .B1(_14886_),
    .X(_15038_));
 sky130_fd_sc_hd__or2b_2 _36692_ (.A(_15037_),
    .B_N(_15038_),
    .X(_15039_));
 sky130_fd_sc_hd__or2b_2 _36693_ (.A(_15038_),
    .B_N(_15037_),
    .X(_15040_));
 sky130_fd_sc_hd__nand3b_2 _36694_ (.A_N(_14858_),
    .B(_14716_),
    .C(_12329_),
    .Y(_15041_));
 sky130_fd_sc_hd__o31a_2 _36695_ (.A1(_14863_),
    .A2(_19175_),
    .A3(_14860_),
    .B1(_15041_),
    .X(_15042_));
 sky130_vsdinv _36696_ (.A(_15042_),
    .Y(_15043_));
 sky130_fd_sc_hd__a21o_2 _36697_ (.A1(_15039_),
    .A2(_15040_),
    .B1(_15043_),
    .X(_15044_));
 sky130_fd_sc_hd__nand3_2 _36698_ (.A(_15039_),
    .B(_15040_),
    .C(_15043_),
    .Y(_15045_));
 sky130_fd_sc_hd__nand2_2 _36699_ (.A(_15044_),
    .B(_15045_),
    .Y(_15046_));
 sky130_fd_sc_hd__o21ai_2 _36700_ (.A1(_15030_),
    .A2(_15032_),
    .B1(_15046_),
    .Y(_15047_));
 sky130_fd_sc_hd__a21o_2 _36701_ (.A1(_15027_),
    .A2(_15028_),
    .B1(_15029_),
    .X(_15048_));
 sky130_fd_sc_hd__nand3b_2 _36702_ (.A_N(_15046_),
    .B(_15048_),
    .C(_15031_),
    .Y(_15049_));
 sky130_fd_sc_hd__o21ba_2 _36703_ (.A1(_14889_),
    .A2(_14891_),
    .B1_N(_14892_),
    .X(_15050_));
 sky130_fd_sc_hd__o21ai_2 _36704_ (.A1(_14896_),
    .A2(_15050_),
    .B1(_14894_),
    .Y(_15051_));
 sky130_fd_sc_hd__a21oi_2 _36705_ (.A1(_15047_),
    .A2(_15049_),
    .B1(_15051_),
    .Y(_15052_));
 sky130_fd_sc_hd__nand3_2 _36706_ (.A(_15047_),
    .B(_15049_),
    .C(_15051_),
    .Y(_15053_));
 sky130_vsdinv _36707_ (.A(_15053_),
    .Y(_15054_));
 sky130_fd_sc_hd__a21boi_2 _36708_ (.A1(_14866_),
    .A2(_14867_),
    .B1_N(_14862_),
    .Y(_15055_));
 sky130_fd_sc_hd__and2_2 _36709_ (.A(_07162_),
    .B(_10900_),
    .X(_15056_));
 sky130_fd_sc_hd__buf_1 _36710_ (.A(_10555_),
    .X(_15057_));
 sky130_fd_sc_hd__a22oi_2 _36711_ (.A1(_08219_),
    .A2(_15057_),
    .B1(_18772_),
    .B2(_10897_),
    .Y(_15058_));
 sky130_fd_sc_hd__and4_2 _36712_ (.A(_12540_),
    .B(_10433_),
    .C(_12871_),
    .D(_19144_),
    .X(_15059_));
 sky130_fd_sc_hd__nor2_2 _36713_ (.A(_15058_),
    .B(_15059_),
    .Y(_15060_));
 sky130_fd_sc_hd__xor2_2 _36714_ (.A(_15056_),
    .B(_15060_),
    .X(_15061_));
 sky130_vsdinv _36715_ (.A(_15061_),
    .Y(_15062_));
 sky130_fd_sc_hd__nand2_2 _36716_ (.A(_14913_),
    .B(_14910_),
    .Y(_15063_));
 sky130_fd_sc_hd__nand2_2 _36717_ (.A(_18748_),
    .B(_10537_),
    .Y(_15064_));
 sky130_fd_sc_hd__nand2_2 _36718_ (.A(_08473_),
    .B(_19156_),
    .Y(_15065_));
 sky130_fd_sc_hd__xor2_2 _36719_ (.A(_15064_),
    .B(_15065_),
    .X(_15066_));
 sky130_fd_sc_hd__and2_2 _36720_ (.A(_12531_),
    .B(_12316_),
    .X(_15067_));
 sky130_fd_sc_hd__nand2_2 _36721_ (.A(_15066_),
    .B(_15067_),
    .Y(_15068_));
 sky130_fd_sc_hd__xnor2_2 _36722_ (.A(_15064_),
    .B(_15065_),
    .Y(_15069_));
 sky130_fd_sc_hd__o21ai_2 _36723_ (.A1(_10736_),
    .A2(_19151_),
    .B1(_15069_),
    .Y(_15070_));
 sky130_fd_sc_hd__nand2_2 _36724_ (.A(_15068_),
    .B(_15070_),
    .Y(_15071_));
 sky130_fd_sc_hd__xor2_2 _36725_ (.A(_15063_),
    .B(_15071_),
    .X(_15072_));
 sky130_fd_sc_hd__nor2_2 _36726_ (.A(_15062_),
    .B(_15072_),
    .Y(_15073_));
 sky130_vsdinv _36727_ (.A(_15073_),
    .Y(_15074_));
 sky130_fd_sc_hd__nand2_2 _36728_ (.A(_15072_),
    .B(_15062_),
    .Y(_15075_));
 sky130_fd_sc_hd__nand3b_2 _36729_ (.A_N(_15055_),
    .B(_15074_),
    .C(_15075_),
    .Y(_15076_));
 sky130_vsdinv _36730_ (.A(_15075_),
    .Y(_15077_));
 sky130_fd_sc_hd__o21ai_2 _36731_ (.A1(_15073_),
    .A2(_15077_),
    .B1(_15055_),
    .Y(_15078_));
 sky130_fd_sc_hd__nand3_2 _36732_ (.A(_14915_),
    .B(_14911_),
    .C(_14913_),
    .Y(_15079_));
 sky130_fd_sc_hd__o21a_2 _36733_ (.A1(_14907_),
    .A2(_14916_),
    .B1(_15079_),
    .X(_15080_));
 sky130_vsdinv _36734_ (.A(_15080_),
    .Y(_15081_));
 sky130_fd_sc_hd__a21o_2 _36735_ (.A1(_15076_),
    .A2(_15078_),
    .B1(_15081_),
    .X(_15082_));
 sky130_fd_sc_hd__nand3_2 _36736_ (.A(_15076_),
    .B(_15078_),
    .C(_15081_),
    .Y(_15083_));
 sky130_fd_sc_hd__nand2_2 _36737_ (.A(_15082_),
    .B(_15083_),
    .Y(_15084_));
 sky130_fd_sc_hd__o21ai_2 _36738_ (.A1(_15052_),
    .A2(_15054_),
    .B1(_15084_),
    .Y(_15085_));
 sky130_fd_sc_hd__a21o_2 _36739_ (.A1(_15047_),
    .A2(_15049_),
    .B1(_15051_),
    .X(_15086_));
 sky130_fd_sc_hd__nand3b_2 _36740_ (.A_N(_15084_),
    .B(_15086_),
    .C(_15053_),
    .Y(_15087_));
 sky130_fd_sc_hd__o21ai_2 _36741_ (.A1(_14927_),
    .A2(_14899_),
    .B1(_14900_),
    .Y(_15088_));
 sky130_fd_sc_hd__a21o_2 _36742_ (.A1(_15085_),
    .A2(_15087_),
    .B1(_15088_),
    .X(_15089_));
 sky130_fd_sc_hd__nand3_2 _36743_ (.A(_15085_),
    .B(_15087_),
    .C(_15088_),
    .Y(_15090_));
 sky130_fd_sc_hd__a21oi_2 _36744_ (.A1(_14905_),
    .A2(_14902_),
    .B1(_14904_),
    .Y(_15091_));
 sky130_fd_sc_hd__o21a_2 _36745_ (.A1(_07392_),
    .A2(_07395_),
    .B1(_11203_),
    .X(_15092_));
 sky130_fd_sc_hd__nand3_2 _36746_ (.A(_14522_),
    .B(_11108_),
    .C(_08013_),
    .Y(_15093_));
 sky130_fd_sc_hd__and3_2 _36747_ (.A(_15092_),
    .B(_14632_),
    .C(_15093_),
    .X(_15094_));
 sky130_vsdinv _36748_ (.A(_15094_),
    .Y(_15095_));
 sky130_fd_sc_hd__a21oi_2 _36749_ (.A1(_15092_),
    .A2(_15093_),
    .B1(_14632_),
    .Y(_15096_));
 sky130_vsdinv _36750_ (.A(_15096_),
    .Y(_15097_));
 sky130_fd_sc_hd__nand3b_2 _36751_ (.A_N(_15091_),
    .B(_15095_),
    .C(_15097_),
    .Y(_15098_));
 sky130_fd_sc_hd__buf_1 _36752_ (.A(_15094_),
    .X(_15099_));
 sky130_fd_sc_hd__buf_1 _36753_ (.A(_15096_),
    .X(_15100_));
 sky130_fd_sc_hd__o21ai_2 _36754_ (.A1(_15099_),
    .A2(_15100_),
    .B1(_15091_),
    .Y(_15101_));
 sky130_fd_sc_hd__o21a_2 _36755_ (.A1(_14826_),
    .A2(_14827_),
    .B1(_14829_),
    .X(_15102_));
 sky130_vsdinv _36756_ (.A(_15102_),
    .Y(_15103_));
 sky130_fd_sc_hd__a21o_2 _36757_ (.A1(_15098_),
    .A2(_15101_),
    .B1(_15103_),
    .X(_15104_));
 sky130_fd_sc_hd__nand3_2 _36758_ (.A(_15103_),
    .B(_15098_),
    .C(_15101_),
    .Y(_15105_));
 sky130_fd_sc_hd__nand2_2 _36759_ (.A(_14839_),
    .B(_14835_),
    .Y(_15106_));
 sky130_fd_sc_hd__a21o_2 _36760_ (.A1(_15104_),
    .A2(_15105_),
    .B1(_15106_),
    .X(_15107_));
 sky130_fd_sc_hd__nand3_2 _36761_ (.A(_15106_),
    .B(_15104_),
    .C(_15105_),
    .Y(_15108_));
 sky130_fd_sc_hd__nand3_2 _36762_ (.A(_15107_),
    .B(_15108_),
    .C(_14656_),
    .Y(_15109_));
 sky130_fd_sc_hd__a21o_2 _36763_ (.A1(_15107_),
    .A2(_15108_),
    .B1(_14655_),
    .X(_15110_));
 sky130_fd_sc_hd__nand2_2 _36764_ (.A(_14926_),
    .B(_14923_),
    .Y(_15111_));
 sky130_fd_sc_hd__a21o_2 _36765_ (.A1(_15109_),
    .A2(_15110_),
    .B1(_15111_),
    .X(_15112_));
 sky130_fd_sc_hd__nand3_2 _36766_ (.A(_15111_),
    .B(_15110_),
    .C(_15109_),
    .Y(_15113_));
 sky130_fd_sc_hd__buf_1 _36767_ (.A(_14655_),
    .X(_15114_));
 sky130_vsdinv _36768_ (.A(_14842_),
    .Y(_15115_));
 sky130_fd_sc_hd__a21oi_2 _36769_ (.A1(_14841_),
    .A2(_15114_),
    .B1(_15115_),
    .Y(_15116_));
 sky130_vsdinv _36770_ (.A(_15116_),
    .Y(_15117_));
 sky130_fd_sc_hd__a21o_2 _36771_ (.A1(_15112_),
    .A2(_15113_),
    .B1(_15117_),
    .X(_15118_));
 sky130_fd_sc_hd__nand3_2 _36772_ (.A(_15112_),
    .B(_15117_),
    .C(_15113_),
    .Y(_15119_));
 sky130_fd_sc_hd__nand2_2 _36773_ (.A(_15118_),
    .B(_15119_),
    .Y(_15120_));
 sky130_fd_sc_hd__buf_1 _36774_ (.A(_15120_),
    .X(_15121_));
 sky130_fd_sc_hd__a21boi_2 _36775_ (.A1(_15089_),
    .A2(_15090_),
    .B1_N(_15121_),
    .Y(_15122_));
 sky130_fd_sc_hd__a21oi_2 _36776_ (.A1(_15085_),
    .A2(_15087_),
    .B1(_15088_),
    .Y(_15123_));
 sky130_vsdinv _36777_ (.A(_15090_),
    .Y(_15124_));
 sky130_fd_sc_hd__nor3_2 _36778_ (.A(_15121_),
    .B(_15123_),
    .C(_15124_),
    .Y(_15125_));
 sky130_fd_sc_hd__o21ai_2 _36779_ (.A1(_14935_),
    .A2(_14853_),
    .B1(_14933_),
    .Y(_15126_));
 sky130_fd_sc_hd__o21bai_2 _36780_ (.A1(_15122_),
    .A2(_15125_),
    .B1_N(_15126_),
    .Y(_15127_));
 sky130_fd_sc_hd__o21ai_2 _36781_ (.A1(_15123_),
    .A2(_15124_),
    .B1(_15121_),
    .Y(_15128_));
 sky130_fd_sc_hd__nand3b_2 _36782_ (.A_N(_15120_),
    .B(_15090_),
    .C(_15089_),
    .Y(_15129_));
 sky130_fd_sc_hd__nand3_2 _36783_ (.A(_15128_),
    .B(_15129_),
    .C(_15126_),
    .Y(_15130_));
 sky130_fd_sc_hd__buf_1 _36784_ (.A(_15130_),
    .X(_15131_));
 sky130_fd_sc_hd__nor3b_2 _36785_ (.A(_14350_),
    .B(_14942_),
    .C_N(_14127_),
    .Y(_15132_));
 sky130_vsdinv _36786_ (.A(_12943_),
    .Y(_15133_));
 sky130_fd_sc_hd__o211ai_2 _36787_ (.A1(_14347_),
    .A2(_14348_),
    .B1(_14350_),
    .C1(_14942_),
    .Y(_15134_));
 sky130_fd_sc_hd__nor3b_2 _36788_ (.A(_15132_),
    .B(_15133_),
    .C_N(_15134_),
    .Y(_15135_));
 sky130_vsdinv _36789_ (.A(_15132_),
    .Y(_15136_));
 sky130_fd_sc_hd__a21oi_2 _36790_ (.A1(_15136_),
    .A2(_15134_),
    .B1(_12943_),
    .Y(_15137_));
 sky130_fd_sc_hd__nor2_2 _36791_ (.A(_15135_),
    .B(_15137_),
    .Y(_15138_));
 sky130_vsdinv _36792_ (.A(_15138_),
    .Y(_15139_));
 sky130_fd_sc_hd__buf_1 _36793_ (.A(_15139_),
    .X(_15140_));
 sky130_fd_sc_hd__a21o_2 _36794_ (.A1(_14852_),
    .A2(_14848_),
    .B1(_15140_),
    .X(_15141_));
 sky130_fd_sc_hd__buf_1 _36795_ (.A(_15139_),
    .X(_15142_));
 sky130_fd_sc_hd__nand3_2 _36796_ (.A(_14852_),
    .B(_14848_),
    .C(_15142_),
    .Y(_15143_));
 sky130_fd_sc_hd__a31oi_2 _36797_ (.A1(_14947_),
    .A2(_14948_),
    .A3(_14955_),
    .B1(_15132_),
    .Y(_15144_));
 sky130_vsdinv _36798_ (.A(_15144_),
    .Y(_15145_));
 sky130_fd_sc_hd__a21o_2 _36799_ (.A1(_15141_),
    .A2(_15143_),
    .B1(_15145_),
    .X(_15146_));
 sky130_fd_sc_hd__nand3b_2 _36800_ (.A_N(_15144_),
    .B(_15141_),
    .C(_15143_),
    .Y(_15147_));
 sky130_fd_sc_hd__nand2_2 _36801_ (.A(_15146_),
    .B(_15147_),
    .Y(_15148_));
 sky130_fd_sc_hd__buf_1 _36802_ (.A(_15148_),
    .X(_15149_));
 sky130_fd_sc_hd__a21boi_2 _36803_ (.A1(_15127_),
    .A2(_15131_),
    .B1_N(_15149_),
    .Y(_15150_));
 sky130_fd_sc_hd__a21oi_2 _36804_ (.A1(_15128_),
    .A2(_15129_),
    .B1(_15126_),
    .Y(_15151_));
 sky130_fd_sc_hd__nor3b_2 _36805_ (.A(_15149_),
    .B(_15151_),
    .C_N(_15131_),
    .Y(_15152_));
 sky130_fd_sc_hd__o21ai_2 _36806_ (.A1(_14959_),
    .A2(_14939_),
    .B1(_14940_),
    .Y(_15153_));
 sky130_fd_sc_hd__o21bai_2 _36807_ (.A1(_15150_),
    .A2(_15152_),
    .B1_N(_15153_),
    .Y(_15154_));
 sky130_vsdinv _36808_ (.A(_15130_),
    .Y(_15155_));
 sky130_fd_sc_hd__o21ai_2 _36809_ (.A1(_15151_),
    .A2(_15155_),
    .B1(_15149_),
    .Y(_15156_));
 sky130_fd_sc_hd__nand3b_2 _36810_ (.A_N(_15148_),
    .B(_15127_),
    .C(_15131_),
    .Y(_15157_));
 sky130_fd_sc_hd__nand3_2 _36811_ (.A(_15156_),
    .B(_15153_),
    .C(_15157_),
    .Y(_15158_));
 sky130_fd_sc_hd__buf_1 _36812_ (.A(_15158_),
    .X(_15159_));
 sky130_fd_sc_hd__buf_1 _36813_ (.A(_13213_),
    .X(_15160_));
 sky130_fd_sc_hd__nand2_2 _36814_ (.A(_14958_),
    .B(_14953_),
    .Y(_15161_));
 sky130_fd_sc_hd__xor2_2 _36815_ (.A(_15160_),
    .B(_15161_),
    .X(_15162_));
 sky130_fd_sc_hd__buf_1 _36816_ (.A(_15162_),
    .X(_15163_));
 sky130_fd_sc_hd__a21oi_2 _36817_ (.A1(_15154_),
    .A2(_15159_),
    .B1(_15163_),
    .Y(_15164_));
 sky130_vsdinv _36818_ (.A(_15162_),
    .Y(_15165_));
 sky130_fd_sc_hd__a21oi_2 _36819_ (.A1(_15156_),
    .A2(_15157_),
    .B1(_15153_),
    .Y(_15166_));
 sky130_fd_sc_hd__nor3b_2 _36820_ (.A(_15165_),
    .B(_15166_),
    .C_N(_15158_),
    .Y(_15167_));
 sky130_vsdinv _36821_ (.A(_14968_),
    .Y(_15168_));
 sky130_fd_sc_hd__o21ai_2 _36822_ (.A1(_15168_),
    .A2(_14964_),
    .B1(_14965_),
    .Y(_15169_));
 sky130_fd_sc_hd__o21bai_2 _36823_ (.A1(_15164_),
    .A2(_15167_),
    .B1_N(_15169_),
    .Y(_15170_));
 sky130_fd_sc_hd__a21o_2 _36824_ (.A1(_15154_),
    .A2(_15158_),
    .B1(_15163_),
    .X(_15171_));
 sky130_fd_sc_hd__nand3_2 _36825_ (.A(_15154_),
    .B(_15163_),
    .C(_15159_),
    .Y(_15172_));
 sky130_fd_sc_hd__nand3_2 _36826_ (.A(_15171_),
    .B(_15169_),
    .C(_15172_),
    .Y(_15173_));
 sky130_fd_sc_hd__a21oi_2 _36827_ (.A1(_14784_),
    .A2(_14779_),
    .B1(_14812_),
    .Y(_15174_));
 sky130_fd_sc_hd__a21oi_2 _36828_ (.A1(_15170_),
    .A2(_15173_),
    .B1(_15174_),
    .Y(_15175_));
 sky130_fd_sc_hd__nand3_2 _36829_ (.A(_15170_),
    .B(_15174_),
    .C(_15173_),
    .Y(_15176_));
 sky130_vsdinv _36830_ (.A(_15176_),
    .Y(_15177_));
 sky130_vsdinv _36831_ (.A(_14977_),
    .Y(_15178_));
 sky130_fd_sc_hd__o21ai_2 _36832_ (.A1(_15178_),
    .A2(_14973_),
    .B1(_14980_),
    .Y(_15179_));
 sky130_fd_sc_hd__o21bai_2 _36833_ (.A1(_15175_),
    .A2(_15177_),
    .B1_N(_15179_),
    .Y(_15180_));
 sky130_fd_sc_hd__buf_1 _36834_ (.A(_14975_),
    .X(_15181_));
 sky130_fd_sc_hd__buf_1 _36835_ (.A(_15181_),
    .X(_15182_));
 sky130_fd_sc_hd__o2bb2ai_2 _36836_ (.A1_N(_15173_),
    .A2_N(_15170_),
    .B1(_15182_),
    .B2(_14967_),
    .Y(_15183_));
 sky130_fd_sc_hd__nand3_2 _36837_ (.A(_15183_),
    .B(_15179_),
    .C(_15176_),
    .Y(_15184_));
 sky130_fd_sc_hd__nand2_2 _36838_ (.A(_15180_),
    .B(_15184_),
    .Y(_15185_));
 sky130_fd_sc_hd__a21oi_2 _36839_ (.A1(_15004_),
    .A2(_14986_),
    .B1(_14985_),
    .Y(_15186_));
 sky130_fd_sc_hd__xor2_2 _36840_ (.A(_15185_),
    .B(_15186_),
    .X(_02668_));
 sky130_fd_sc_hd__a21oi_2 _36841_ (.A1(_15014_),
    .A2(_15005_),
    .B1(_15008_),
    .Y(_15187_));
 sky130_vsdinv _36842_ (.A(_15187_),
    .Y(_15188_));
 sky130_fd_sc_hd__and2_2 _36843_ (.A(_10484_),
    .B(_08553_),
    .X(_15189_));
 sky130_fd_sc_hd__a22oi_2 _36844_ (.A1(_18695_),
    .A2(_07751_),
    .B1(_19208_),
    .B2(_10997_),
    .Y(_15190_));
 sky130_fd_sc_hd__nand2_2 _36845_ (.A(_14871_),
    .B(_10383_),
    .Y(_15191_));
 sky130_fd_sc_hd__nor3_2 _36846_ (.A(_08300_),
    .B(_11332_),
    .C(_15191_),
    .Y(_15192_));
 sky130_fd_sc_hd__nor2_2 _36847_ (.A(_15190_),
    .B(_15192_),
    .Y(_15193_));
 sky130_fd_sc_hd__xor2_2 _36848_ (.A(_15189_),
    .B(_15193_),
    .X(_15194_));
 sky130_fd_sc_hd__nor2_2 _36849_ (.A(_15188_),
    .B(_15194_),
    .Y(_15195_));
 sky130_fd_sc_hd__nand2_2 _36850_ (.A(_15194_),
    .B(_15188_),
    .Y(_15196_));
 sky130_vsdinv _36851_ (.A(_15196_),
    .Y(_15197_));
 sky130_fd_sc_hd__and2_2 _36852_ (.A(_09321_),
    .B(_12839_),
    .X(_15198_));
 sky130_fd_sc_hd__buf_1 _36853_ (.A(_18717_),
    .X(_15199_));
 sky130_fd_sc_hd__a22oi_2 _36854_ (.A1(_15023_),
    .A2(_11441_),
    .B1(_15199_),
    .B2(_09104_),
    .Y(_15200_));
 sky130_fd_sc_hd__and4_2 _36855_ (.A(_10261_),
    .B(_10687_),
    .C(_09079_),
    .D(_09078_),
    .X(_15201_));
 sky130_fd_sc_hd__nor2_2 _36856_ (.A(_15200_),
    .B(_15201_),
    .Y(_15202_));
 sky130_fd_sc_hd__xor2_2 _36857_ (.A(_15198_),
    .B(_15202_),
    .X(_15203_));
 sky130_fd_sc_hd__o21bai_2 _36858_ (.A1(_15195_),
    .A2(_15197_),
    .B1_N(_15203_),
    .Y(_15204_));
 sky130_fd_sc_hd__nand3b_2 _36859_ (.A_N(_15195_),
    .B(_15196_),
    .C(_15203_),
    .Y(_15205_));
 sky130_fd_sc_hd__nand2_2 _36860_ (.A(_15028_),
    .B(_15016_),
    .Y(_15206_));
 sky130_fd_sc_hd__a21oi_2 _36861_ (.A1(_15204_),
    .A2(_15205_),
    .B1(_15206_),
    .Y(_15207_));
 sky130_fd_sc_hd__nand3_2 _36862_ (.A(_15204_),
    .B(_15206_),
    .C(_15205_),
    .Y(_15208_));
 sky130_vsdinv _36863_ (.A(_15208_),
    .Y(_15209_));
 sky130_fd_sc_hd__nand3b_2 _36864_ (.A_N(_15034_),
    .B(_18737_),
    .C(_12330_),
    .Y(_15210_));
 sky130_fd_sc_hd__o31a_2 _36865_ (.A1(_14863_),
    .A2(_19169_),
    .A3(_15036_),
    .B1(_15210_),
    .X(_15211_));
 sky130_fd_sc_hd__a21o_2 _36866_ (.A1(_15025_),
    .A2(_15018_),
    .B1(_15024_),
    .X(_15212_));
 sky130_fd_sc_hd__nand2_2 _36867_ (.A(_18728_),
    .B(_09497_),
    .Y(_15213_));
 sky130_fd_sc_hd__nand2_2 _36868_ (.A(_09313_),
    .B(_19167_),
    .Y(_15214_));
 sky130_fd_sc_hd__xor2_2 _36869_ (.A(_15213_),
    .B(_15214_),
    .X(_15215_));
 sky130_fd_sc_hd__nand3_2 _36870_ (.A(_15215_),
    .B(_08459_),
    .C(_14666_),
    .Y(_15216_));
 sky130_fd_sc_hd__xnor2_2 _36871_ (.A(_15213_),
    .B(_15214_),
    .Y(_15217_));
 sky130_fd_sc_hd__o21ai_2 _36872_ (.A1(_18742_),
    .A2(_19164_),
    .B1(_15217_),
    .Y(_15218_));
 sky130_fd_sc_hd__nand2_2 _36873_ (.A(_15216_),
    .B(_15218_),
    .Y(_15219_));
 sky130_fd_sc_hd__xor2_2 _36874_ (.A(_15212_),
    .B(_15219_),
    .X(_15220_));
 sky130_fd_sc_hd__xor2_2 _36875_ (.A(_15211_),
    .B(_15220_),
    .X(_15221_));
 sky130_fd_sc_hd__o21bai_2 _36876_ (.A1(_15207_),
    .A2(_15209_),
    .B1_N(_15221_),
    .Y(_15222_));
 sky130_fd_sc_hd__a21o_2 _36877_ (.A1(_15204_),
    .A2(_15205_),
    .B1(_15206_),
    .X(_15223_));
 sky130_fd_sc_hd__nand3_2 _36878_ (.A(_15223_),
    .B(_15221_),
    .C(_15208_),
    .Y(_15224_));
 sky130_fd_sc_hd__o21ai_2 _36879_ (.A1(_15030_),
    .A2(_15046_),
    .B1(_15031_),
    .Y(_15225_));
 sky130_fd_sc_hd__a21oi_2 _36880_ (.A1(_15222_),
    .A2(_15224_),
    .B1(_15225_),
    .Y(_15226_));
 sky130_fd_sc_hd__nand3_2 _36881_ (.A(_15222_),
    .B(_15224_),
    .C(_15225_),
    .Y(_15227_));
 sky130_vsdinv _36882_ (.A(_15227_),
    .Y(_15228_));
 sky130_fd_sc_hd__nand2_2 _36883_ (.A(_12527_),
    .B(_09802_),
    .Y(_15229_));
 sky130_fd_sc_hd__nand2_2 _36884_ (.A(_12794_),
    .B(_10877_),
    .Y(_15230_));
 sky130_fd_sc_hd__xor2_2 _36885_ (.A(_15229_),
    .B(_15230_),
    .X(_15231_));
 sky130_fd_sc_hd__and2_2 _36886_ (.A(_07846_),
    .B(_15057_),
    .X(_15232_));
 sky130_fd_sc_hd__nand2_2 _36887_ (.A(_15231_),
    .B(_15232_),
    .Y(_15233_));
 sky130_fd_sc_hd__xnor2_2 _36888_ (.A(_15229_),
    .B(_15230_),
    .Y(_15234_));
 sky130_fd_sc_hd__o21ai_2 _36889_ (.A1(_18761_),
    .A2(_19146_),
    .B1(_15234_),
    .Y(_15235_));
 sky130_fd_sc_hd__nand2_2 _36890_ (.A(_15233_),
    .B(_15235_),
    .Y(_15236_));
 sky130_fd_sc_hd__o211ai_2 _36891_ (.A1(_15064_),
    .A2(_15065_),
    .B1(_15068_),
    .C1(_15236_),
    .Y(_15237_));
 sky130_fd_sc_hd__o21ai_2 _36892_ (.A1(_15064_),
    .A2(_15065_),
    .B1(_15068_),
    .Y(_15238_));
 sky130_fd_sc_hd__nand3_2 _36893_ (.A(_15238_),
    .B(_15235_),
    .C(_15233_),
    .Y(_15239_));
 sky130_fd_sc_hd__nand2_2 _36894_ (.A(_15237_),
    .B(_15239_),
    .Y(_15240_));
 sky130_fd_sc_hd__and2_2 _36895_ (.A(_14522_),
    .B(_11064_),
    .X(_15241_));
 sky130_fd_sc_hd__buf_1 _36896_ (.A(_15241_),
    .X(_15242_));
 sky130_fd_sc_hd__nand2_2 _36897_ (.A(_12540_),
    .B(_12871_),
    .Y(_15243_));
 sky130_fd_sc_hd__nand2_2 _36898_ (.A(_12806_),
    .B(_12905_),
    .Y(_15244_));
 sky130_fd_sc_hd__xnor2_2 _36899_ (.A(_15243_),
    .B(_15244_),
    .Y(_15245_));
 sky130_fd_sc_hd__xor2_2 _36900_ (.A(_15242_),
    .B(_15245_),
    .X(_15246_));
 sky130_fd_sc_hd__nand2_2 _36901_ (.A(_15240_),
    .B(_15246_),
    .Y(_15247_));
 sky130_fd_sc_hd__nand3b_2 _36902_ (.A_N(_15246_),
    .B(_15237_),
    .C(_15239_),
    .Y(_15248_));
 sky130_vsdinv _36903_ (.A(_15039_),
    .Y(_15249_));
 sky130_fd_sc_hd__a221o_2 _36904_ (.A1(_15043_),
    .A2(_15040_),
    .B1(_15247_),
    .B2(_15248_),
    .C1(_15249_),
    .X(_15250_));
 sky130_fd_sc_hd__a21boi_2 _36905_ (.A1(_15043_),
    .A2(_15040_),
    .B1_N(_15039_),
    .Y(_15251_));
 sky130_fd_sc_hd__nand3b_2 _36906_ (.A_N(_15251_),
    .B(_15248_),
    .C(_15247_),
    .Y(_15252_));
 sky130_fd_sc_hd__nand2_2 _36907_ (.A(_15250_),
    .B(_15252_),
    .Y(_15253_));
 sky130_fd_sc_hd__nand3_2 _36908_ (.A(_15068_),
    .B(_15070_),
    .C(_15063_),
    .Y(_15254_));
 sky130_fd_sc_hd__o21a_2 _36909_ (.A1(_15062_),
    .A2(_15072_),
    .B1(_15254_),
    .X(_15255_));
 sky130_fd_sc_hd__nand2_2 _36910_ (.A(_15253_),
    .B(_15255_),
    .Y(_15256_));
 sky130_fd_sc_hd__nand3b_2 _36911_ (.A_N(_15255_),
    .B(_15250_),
    .C(_15252_),
    .Y(_15257_));
 sky130_fd_sc_hd__nand2_2 _36912_ (.A(_15256_),
    .B(_15257_),
    .Y(_15258_));
 sky130_fd_sc_hd__o21ai_2 _36913_ (.A1(_15226_),
    .A2(_15228_),
    .B1(_15258_),
    .Y(_15259_));
 sky130_fd_sc_hd__a21o_2 _36914_ (.A1(_15222_),
    .A2(_15224_),
    .B1(_15225_),
    .X(_15260_));
 sky130_fd_sc_hd__nand3b_2 _36915_ (.A_N(_15258_),
    .B(_15260_),
    .C(_15227_),
    .Y(_15261_));
 sky130_fd_sc_hd__o21ai_2 _36916_ (.A1(_15084_),
    .A2(_15052_),
    .B1(_15053_),
    .Y(_15262_));
 sky130_fd_sc_hd__a21o_2 _36917_ (.A1(_15259_),
    .A2(_15261_),
    .B1(_15262_),
    .X(_15263_));
 sky130_fd_sc_hd__nand3_2 _36918_ (.A(_15259_),
    .B(_15261_),
    .C(_15262_),
    .Y(_15264_));
 sky130_fd_sc_hd__buf_1 _36919_ (.A(_15094_),
    .X(_15265_));
 sky130_fd_sc_hd__buf_1 _36920_ (.A(_15096_),
    .X(_15266_));
 sky130_fd_sc_hd__a21oi_2 _36921_ (.A1(_15060_),
    .A2(_15056_),
    .B1(_15059_),
    .Y(_15267_));
 sky130_fd_sc_hd__o21a_2 _36922_ (.A1(_15265_),
    .A2(_15266_),
    .B1(_15267_),
    .X(_15268_));
 sky130_fd_sc_hd__nor3_2 _36923_ (.A(_15099_),
    .B(_15100_),
    .C(_15267_),
    .Y(_15269_));
 sky130_vsdinv _36924_ (.A(_15093_),
    .Y(_15270_));
 sky130_fd_sc_hd__a21oi_2 _36925_ (.A1(_15092_),
    .A2(_14633_),
    .B1(_15270_),
    .Y(_15271_));
 sky130_vsdinv _36926_ (.A(_15271_),
    .Y(_15272_));
 sky130_fd_sc_hd__o21bai_2 _36927_ (.A1(_15268_),
    .A2(_15269_),
    .B1_N(_15272_),
    .Y(_15273_));
 sky130_fd_sc_hd__nand3b_2 _36928_ (.A_N(_15267_),
    .B(_15095_),
    .C(_15097_),
    .Y(_15274_));
 sky130_fd_sc_hd__buf_1 _36929_ (.A(_15272_),
    .X(_15275_));
 sky130_fd_sc_hd__nand3b_2 _36930_ (.A_N(_15268_),
    .B(_15274_),
    .C(_15275_),
    .Y(_15276_));
 sky130_fd_sc_hd__nand2_2 _36931_ (.A(_15105_),
    .B(_15098_),
    .Y(_15277_));
 sky130_fd_sc_hd__a21oi_2 _36932_ (.A1(_15273_),
    .A2(_15276_),
    .B1(_15277_),
    .Y(_15278_));
 sky130_fd_sc_hd__nand3_2 _36933_ (.A(_15277_),
    .B(_15273_),
    .C(_15276_),
    .Y(_15279_));
 sky130_fd_sc_hd__nor3b_2 _36934_ (.A(_14652_),
    .B(_15278_),
    .C_N(_15279_),
    .Y(_15280_));
 sky130_vsdinv _36935_ (.A(_15279_),
    .Y(_15281_));
 sky130_fd_sc_hd__o21a_2 _36936_ (.A1(_15278_),
    .A2(_15281_),
    .B1(_14652_),
    .X(_15282_));
 sky130_fd_sc_hd__o211ai_2 _36937_ (.A1(_15280_),
    .A2(_15282_),
    .B1(_15076_),
    .C1(_15083_),
    .Y(_15283_));
 sky130_fd_sc_hd__nand2_2 _36938_ (.A(_15083_),
    .B(_15076_),
    .Y(_15284_));
 sky130_vsdinv _36939_ (.A(_15280_),
    .Y(_15285_));
 sky130_fd_sc_hd__nand3b_2 _36940_ (.A_N(_15282_),
    .B(_15284_),
    .C(_15285_),
    .Y(_15286_));
 sky130_fd_sc_hd__a21boi_2 _36941_ (.A1(_15107_),
    .A2(_14843_),
    .B1_N(_15108_),
    .Y(_15287_));
 sky130_vsdinv _36942_ (.A(_15287_),
    .Y(_15288_));
 sky130_fd_sc_hd__a21o_2 _36943_ (.A1(_15283_),
    .A2(_15286_),
    .B1(_15288_),
    .X(_15289_));
 sky130_fd_sc_hd__nand3_2 _36944_ (.A(_15283_),
    .B(_15286_),
    .C(_15288_),
    .Y(_15290_));
 sky130_fd_sc_hd__nand2_2 _36945_ (.A(_15289_),
    .B(_15290_),
    .Y(_15291_));
 sky130_fd_sc_hd__buf_1 _36946_ (.A(_15291_),
    .X(_15292_));
 sky130_fd_sc_hd__a21boi_2 _36947_ (.A1(_15263_),
    .A2(_15264_),
    .B1_N(_15292_),
    .Y(_15293_));
 sky130_fd_sc_hd__a21oi_2 _36948_ (.A1(_15259_),
    .A2(_15261_),
    .B1(_15262_),
    .Y(_15294_));
 sky130_fd_sc_hd__nor3b_2 _36949_ (.A(_15292_),
    .B(_15294_),
    .C_N(_15264_),
    .Y(_15295_));
 sky130_fd_sc_hd__o21ai_2 _36950_ (.A1(_15121_),
    .A2(_15123_),
    .B1(_15090_),
    .Y(_15296_));
 sky130_fd_sc_hd__o21bai_2 _36951_ (.A1(_15293_),
    .A2(_15295_),
    .B1_N(_15296_),
    .Y(_15297_));
 sky130_fd_sc_hd__and3_2 _36952_ (.A(_15259_),
    .B(_15261_),
    .C(_15262_),
    .X(_15298_));
 sky130_fd_sc_hd__o21ai_2 _36953_ (.A1(_15294_),
    .A2(_15298_),
    .B1(_15292_),
    .Y(_15299_));
 sky130_fd_sc_hd__nand3b_2 _36954_ (.A_N(_15292_),
    .B(_15263_),
    .C(_15264_),
    .Y(_15300_));
 sky130_fd_sc_hd__nand3_2 _36955_ (.A(_15299_),
    .B(_15300_),
    .C(_15296_),
    .Y(_15301_));
 sky130_fd_sc_hd__a21o_2 _36956_ (.A1(_15119_),
    .A2(_15113_),
    .B1(_15142_),
    .X(_15302_));
 sky130_fd_sc_hd__buf_1 _36957_ (.A(_15139_),
    .X(_15303_));
 sky130_fd_sc_hd__nand3_2 _36958_ (.A(_15119_),
    .B(_15303_),
    .C(_15113_),
    .Y(_15304_));
 sky130_fd_sc_hd__a21oi_2 _36959_ (.A1(_13184_),
    .A2(_15134_),
    .B1(_15132_),
    .Y(_15305_));
 sky130_vsdinv _36960_ (.A(_15305_),
    .Y(_15306_));
 sky130_fd_sc_hd__buf_1 _36961_ (.A(_15306_),
    .X(_15307_));
 sky130_fd_sc_hd__a21o_2 _36962_ (.A1(_15302_),
    .A2(_15304_),
    .B1(_15307_),
    .X(_15308_));
 sky130_fd_sc_hd__buf_1 _36963_ (.A(_15306_),
    .X(_15309_));
 sky130_fd_sc_hd__nand3_2 _36964_ (.A(_15302_),
    .B(_15309_),
    .C(_15304_),
    .Y(_15310_));
 sky130_fd_sc_hd__nand2_2 _36965_ (.A(_15308_),
    .B(_15310_),
    .Y(_15311_));
 sky130_vsdinv _36966_ (.A(_15311_),
    .Y(_15312_));
 sky130_fd_sc_hd__a21oi_2 _36967_ (.A1(_15297_),
    .A2(_15301_),
    .B1(_15312_),
    .Y(_15313_));
 sky130_fd_sc_hd__a21oi_2 _36968_ (.A1(_15299_),
    .A2(_15300_),
    .B1(_15296_),
    .Y(_15314_));
 sky130_vsdinv _36969_ (.A(_15301_),
    .Y(_15315_));
 sky130_fd_sc_hd__nor3_2 _36970_ (.A(_15311_),
    .B(_15314_),
    .C(_15315_),
    .Y(_15316_));
 sky130_fd_sc_hd__o21ai_2 _36971_ (.A1(_15149_),
    .A2(_15151_),
    .B1(_15131_),
    .Y(_15317_));
 sky130_fd_sc_hd__o21bai_2 _36972_ (.A1(_15313_),
    .A2(_15316_),
    .B1_N(_15317_),
    .Y(_15318_));
 sky130_fd_sc_hd__o21ai_2 _36973_ (.A1(_15314_),
    .A2(_15315_),
    .B1(_15311_),
    .Y(_15319_));
 sky130_fd_sc_hd__nand3_2 _36974_ (.A(_15297_),
    .B(_15312_),
    .C(_15301_),
    .Y(_15320_));
 sky130_fd_sc_hd__nand3_2 _36975_ (.A(_15319_),
    .B(_15320_),
    .C(_15317_),
    .Y(_15321_));
 sky130_fd_sc_hd__nand2_2 _36976_ (.A(_15147_),
    .B(_15141_),
    .Y(_15322_));
 sky130_fd_sc_hd__xor2_2 _36977_ (.A(_15160_),
    .B(_15322_),
    .X(_15323_));
 sky130_fd_sc_hd__a21oi_2 _36978_ (.A1(_15318_),
    .A2(_15321_),
    .B1(_15323_),
    .Y(_15324_));
 sky130_fd_sc_hd__nand3_2 _36979_ (.A(_15318_),
    .B(_15323_),
    .C(_15321_),
    .Y(_15325_));
 sky130_vsdinv _36980_ (.A(_15325_),
    .Y(_15326_));
 sky130_fd_sc_hd__o21ai_2 _36981_ (.A1(_15165_),
    .A2(_15166_),
    .B1(_15159_),
    .Y(_15327_));
 sky130_fd_sc_hd__o21bai_2 _36982_ (.A1(_15324_),
    .A2(_15326_),
    .B1_N(_15327_),
    .Y(_15328_));
 sky130_fd_sc_hd__nand3b_2 _36983_ (.A_N(_15324_),
    .B(_15325_),
    .C(_15327_),
    .Y(_15329_));
 sky130_fd_sc_hd__a21oi_2 _36984_ (.A1(_14958_),
    .A2(_14953_),
    .B1(_15181_),
    .Y(_15330_));
 sky130_fd_sc_hd__a21o_2 _36985_ (.A1(_15328_),
    .A2(_15329_),
    .B1(_15330_),
    .X(_15331_));
 sky130_fd_sc_hd__nand3_2 _36986_ (.A(_15328_),
    .B(_15329_),
    .C(_15330_),
    .Y(_15332_));
 sky130_fd_sc_hd__nand2_2 _36987_ (.A(_15176_),
    .B(_15173_),
    .Y(_15333_));
 sky130_fd_sc_hd__a21oi_2 _36988_ (.A1(_15331_),
    .A2(_15332_),
    .B1(_15333_),
    .Y(_15334_));
 sky130_fd_sc_hd__nand3_2 _36989_ (.A(_15331_),
    .B(_15333_),
    .C(_15332_),
    .Y(_15335_));
 sky130_vsdinv _36990_ (.A(_15335_),
    .Y(_15336_));
 sky130_fd_sc_hd__nor2_2 _36991_ (.A(_15334_),
    .B(_15336_),
    .Y(_15337_));
 sky130_fd_sc_hd__nor3_2 _36992_ (.A(_14985_),
    .B(_14983_),
    .C(_15185_),
    .Y(_15338_));
 sky130_fd_sc_hd__a21oi_2 _36993_ (.A1(_15183_),
    .A2(_15176_),
    .B1(_15179_),
    .Y(_15339_));
 sky130_fd_sc_hd__a21oi_2 _36994_ (.A1(_14984_),
    .A2(_15184_),
    .B1(_15339_),
    .Y(_15340_));
 sky130_fd_sc_hd__a21oi_2 _36995_ (.A1(_15004_),
    .A2(_15338_),
    .B1(_15340_),
    .Y(_15341_));
 sky130_fd_sc_hd__xnor2_2 _36996_ (.A(_15337_),
    .B(_15341_),
    .Y(_02669_));
 sky130_fd_sc_hd__and2_2 _36997_ (.A(_09321_),
    .B(_10583_),
    .X(_15342_));
 sky130_fd_sc_hd__a22oi_2 _36998_ (.A1(_18712_),
    .A2(_08827_),
    .B1(_15199_),
    .B2(_12839_),
    .Y(_15343_));
 sky130_fd_sc_hd__and4_2 _36999_ (.A(_14884_),
    .B(_15020_),
    .C(_12836_),
    .D(_12295_),
    .X(_15344_));
 sky130_fd_sc_hd__nor2_2 _37000_ (.A(_15343_),
    .B(_15344_),
    .Y(_15345_));
 sky130_fd_sc_hd__xor2_2 _37001_ (.A(_15342_),
    .B(_15345_),
    .X(_15346_));
 sky130_vsdinv _37002_ (.A(_15346_),
    .Y(_15347_));
 sky130_vsdinv _37003_ (.A(_15190_),
    .Y(_15348_));
 sky130_fd_sc_hd__a21oi_2 _37004_ (.A1(_15348_),
    .A2(_15189_),
    .B1(_15192_),
    .Y(_15349_));
 sky130_vsdinv _37005_ (.A(_15349_),
    .Y(_15350_));
 sky130_fd_sc_hd__and2_2 _37006_ (.A(_10484_),
    .B(_08310_),
    .X(_15351_));
 sky130_fd_sc_hd__a22oi_2 _37007_ (.A1(_18695_),
    .A2(_07961_),
    .B1(_19204_),
    .B2(_10997_),
    .Y(_15352_));
 sky130_fd_sc_hd__nand2_2 _37008_ (.A(_10481_),
    .B(_08812_),
    .Y(_15353_));
 sky130_fd_sc_hd__nor3_2 _37009_ (.A(_07751_),
    .B(_11005_),
    .C(_15353_),
    .Y(_15354_));
 sky130_fd_sc_hd__nor2_2 _37010_ (.A(_15352_),
    .B(_15354_),
    .Y(_15355_));
 sky130_fd_sc_hd__xor2_2 _37011_ (.A(_15351_),
    .B(_15355_),
    .X(_15356_));
 sky130_fd_sc_hd__nor2_2 _37012_ (.A(_15350_),
    .B(_15356_),
    .Y(_15357_));
 sky130_fd_sc_hd__nand2_2 _37013_ (.A(_15356_),
    .B(_15350_),
    .Y(_15358_));
 sky130_fd_sc_hd__buf_1 _37014_ (.A(_15358_),
    .X(_15359_));
 sky130_fd_sc_hd__nor3b_2 _37015_ (.A(_15347_),
    .B(_15357_),
    .C_N(_15359_),
    .Y(_15360_));
 sky130_fd_sc_hd__or2b_2 _37016_ (.A(_15356_),
    .B_N(_15349_),
    .X(_15361_));
 sky130_fd_sc_hd__a21oi_2 _37017_ (.A1(_15361_),
    .A2(_15359_),
    .B1(_15346_),
    .Y(_15362_));
 sky130_vsdinv _37018_ (.A(_15203_),
    .Y(_15363_));
 sky130_fd_sc_hd__o21ai_2 _37019_ (.A1(_15363_),
    .A2(_15195_),
    .B1(_15196_),
    .Y(_15364_));
 sky130_fd_sc_hd__o21bai_2 _37020_ (.A1(_15360_),
    .A2(_15362_),
    .B1_N(_15364_),
    .Y(_15365_));
 sky130_vsdinv _37021_ (.A(_15358_),
    .Y(_15366_));
 sky130_fd_sc_hd__o21bai_2 _37022_ (.A1(_15357_),
    .A2(_15366_),
    .B1_N(_15346_),
    .Y(_15367_));
 sky130_fd_sc_hd__nand3_2 _37023_ (.A(_15361_),
    .B(_15359_),
    .C(_15346_),
    .Y(_15368_));
 sky130_fd_sc_hd__nand3_2 _37024_ (.A(_15367_),
    .B(_15368_),
    .C(_15364_),
    .Y(_15369_));
 sky130_fd_sc_hd__nand2_2 _37025_ (.A(_15365_),
    .B(_15369_),
    .Y(_15370_));
 sky130_fd_sc_hd__o21a_2 _37026_ (.A1(_15213_),
    .A2(_15214_),
    .B1(_15216_),
    .X(_15371_));
 sky130_vsdinv _37027_ (.A(_15371_),
    .Y(_15372_));
 sky130_fd_sc_hd__nand2_2 _37028_ (.A(_14857_),
    .B(_19167_),
    .Y(_15373_));
 sky130_fd_sc_hd__nand2_2 _37029_ (.A(_09313_),
    .B(_10042_),
    .Y(_15374_));
 sky130_fd_sc_hd__xnor2_2 _37030_ (.A(_15373_),
    .B(_15374_),
    .Y(_15375_));
 sky130_fd_sc_hd__buf_1 _37031_ (.A(_13026_),
    .X(_15376_));
 sky130_fd_sc_hd__nand3b_2 _37032_ (.A_N(_15375_),
    .B(_15376_),
    .C(_13369_),
    .Y(_15377_));
 sky130_fd_sc_hd__o21ai_2 _37033_ (.A1(_14863_),
    .A2(_19159_),
    .B1(_15375_),
    .Y(_15378_));
 sky130_fd_sc_hd__a21o_2 _37034_ (.A1(_15202_),
    .A2(_15198_),
    .B1(_15201_),
    .X(_15379_));
 sky130_fd_sc_hd__a21o_2 _37035_ (.A1(_15377_),
    .A2(_15378_),
    .B1(_15379_),
    .X(_15380_));
 sky130_fd_sc_hd__nand3_2 _37036_ (.A(_15379_),
    .B(_15377_),
    .C(_15378_),
    .Y(_15381_));
 sky130_fd_sc_hd__nand2_2 _37037_ (.A(_15380_),
    .B(_15381_),
    .Y(_15382_));
 sky130_fd_sc_hd__xor2_2 _37038_ (.A(_15372_),
    .B(_15382_),
    .X(_15383_));
 sky130_fd_sc_hd__nand2_2 _37039_ (.A(_15370_),
    .B(_15383_),
    .Y(_15384_));
 sky130_fd_sc_hd__nand3b_2 _37040_ (.A_N(_15383_),
    .B(_15365_),
    .C(_15369_),
    .Y(_15385_));
 sky130_vsdinv _37041_ (.A(_15211_),
    .Y(_15386_));
 sky130_fd_sc_hd__xor2_2 _37042_ (.A(_15386_),
    .B(_15220_),
    .X(_15387_));
 sky130_fd_sc_hd__o21ai_2 _37043_ (.A1(_15207_),
    .A2(_15387_),
    .B1(_15208_),
    .Y(_15388_));
 sky130_fd_sc_hd__a21o_2 _37044_ (.A1(_15384_),
    .A2(_15385_),
    .B1(_15388_),
    .X(_15389_));
 sky130_fd_sc_hd__nand3_2 _37045_ (.A(_15388_),
    .B(_15384_),
    .C(_15385_),
    .Y(_15390_));
 sky130_fd_sc_hd__buf_1 _37046_ (.A(_15390_),
    .X(_15391_));
 sky130_fd_sc_hd__a21oi_2 _37047_ (.A1(_15218_),
    .A2(_15216_),
    .B1(_15212_),
    .Y(_15392_));
 sky130_fd_sc_hd__nand3_2 _37048_ (.A(_15212_),
    .B(_15218_),
    .C(_15216_),
    .Y(_15393_));
 sky130_fd_sc_hd__nand3b_2 _37049_ (.A_N(_15392_),
    .B(_15386_),
    .C(_15393_),
    .Y(_15394_));
 sky130_fd_sc_hd__nand2_2 _37050_ (.A(_14245_),
    .B(_12316_),
    .Y(_15395_));
 sky130_fd_sc_hd__nand2_2 _37051_ (.A(_18754_),
    .B(_19144_),
    .Y(_15396_));
 sky130_fd_sc_hd__xor2_2 _37052_ (.A(_15395_),
    .B(_15396_),
    .X(_15397_));
 sky130_fd_sc_hd__and2_2 _37053_ (.A(_07846_),
    .B(_11199_),
    .X(_15398_));
 sky130_fd_sc_hd__nand2_2 _37054_ (.A(_15397_),
    .B(_15398_),
    .Y(_15399_));
 sky130_fd_sc_hd__xnor2_2 _37055_ (.A(_15395_),
    .B(_15396_),
    .Y(_15400_));
 sky130_fd_sc_hd__o21ai_2 _37056_ (.A1(_18761_),
    .A2(_19141_),
    .B1(_15400_),
    .Y(_15401_));
 sky130_fd_sc_hd__nand2_2 _37057_ (.A(_15399_),
    .B(_15401_),
    .Y(_15402_));
 sky130_fd_sc_hd__o211ai_2 _37058_ (.A1(_15229_),
    .A2(_15230_),
    .B1(_15233_),
    .C1(_15402_),
    .Y(_15403_));
 sky130_fd_sc_hd__o21ai_2 _37059_ (.A1(_15229_),
    .A2(_15230_),
    .B1(_15233_),
    .Y(_15404_));
 sky130_fd_sc_hd__nand3_2 _37060_ (.A(_15404_),
    .B(_15401_),
    .C(_15399_),
    .Y(_15405_));
 sky130_fd_sc_hd__nand2_2 _37061_ (.A(_12847_),
    .B(_10900_),
    .Y(_15406_));
 sky130_fd_sc_hd__nand2_2 _37062_ (.A(_14648_),
    .B(_18772_),
    .Y(_15407_));
 sky130_fd_sc_hd__xnor2_2 _37063_ (.A(_15406_),
    .B(_15407_),
    .Y(_15408_));
 sky130_fd_sc_hd__xor2_2 _37064_ (.A(_15242_),
    .B(_15408_),
    .X(_15409_));
 sky130_fd_sc_hd__a21boi_2 _37065_ (.A1(_15403_),
    .A2(_15405_),
    .B1_N(_15409_),
    .Y(_15410_));
 sky130_fd_sc_hd__nand2_2 _37066_ (.A(_15403_),
    .B(_15405_),
    .Y(_15411_));
 sky130_fd_sc_hd__nor2_2 _37067_ (.A(_15409_),
    .B(_15411_),
    .Y(_15412_));
 sky130_fd_sc_hd__a211o_2 _37068_ (.A1(_15394_),
    .A2(_15393_),
    .B1(_15410_),
    .C1(_15412_),
    .X(_15413_));
 sky130_fd_sc_hd__o211ai_2 _37069_ (.A1(_15410_),
    .A2(_15412_),
    .B1(_15393_),
    .C1(_15394_),
    .Y(_15414_));
 sky130_fd_sc_hd__o21a_2 _37070_ (.A1(_15246_),
    .A2(_15240_),
    .B1(_15239_),
    .X(_15415_));
 sky130_vsdinv _37071_ (.A(_15415_),
    .Y(_15416_));
 sky130_fd_sc_hd__a21o_2 _37072_ (.A1(_15413_),
    .A2(_15414_),
    .B1(_15416_),
    .X(_15417_));
 sky130_fd_sc_hd__nand3_2 _37073_ (.A(_15413_),
    .B(_15416_),
    .C(_15414_),
    .Y(_15418_));
 sky130_fd_sc_hd__nand2_2 _37074_ (.A(_15417_),
    .B(_15418_),
    .Y(_15419_));
 sky130_fd_sc_hd__buf_1 _37075_ (.A(_15419_),
    .X(_15420_));
 sky130_fd_sc_hd__a21boi_2 _37076_ (.A1(_15389_),
    .A2(_15391_),
    .B1_N(_15420_),
    .Y(_15421_));
 sky130_fd_sc_hd__a21oi_2 _37077_ (.A1(_15384_),
    .A2(_15385_),
    .B1(_15388_),
    .Y(_15422_));
 sky130_fd_sc_hd__nor3b_2 _37078_ (.A(_15420_),
    .B(_15422_),
    .C_N(_15391_),
    .Y(_15423_));
 sky130_fd_sc_hd__o21ai_2 _37079_ (.A1(_15258_),
    .A2(_15226_),
    .B1(_15227_),
    .Y(_15424_));
 sky130_fd_sc_hd__o21bai_2 _37080_ (.A1(_15421_),
    .A2(_15423_),
    .B1_N(_15424_),
    .Y(_15425_));
 sky130_vsdinv _37081_ (.A(_15390_),
    .Y(_15426_));
 sky130_fd_sc_hd__o21ai_2 _37082_ (.A1(_15422_),
    .A2(_15426_),
    .B1(_15420_),
    .Y(_15427_));
 sky130_fd_sc_hd__nand3b_2 _37083_ (.A_N(_15419_),
    .B(_15389_),
    .C(_15391_),
    .Y(_15428_));
 sky130_fd_sc_hd__nand3_2 _37084_ (.A(_15427_),
    .B(_15428_),
    .C(_15424_),
    .Y(_15429_));
 sky130_vsdinv _37085_ (.A(_15241_),
    .Y(_15430_));
 sky130_fd_sc_hd__nor2_2 _37086_ (.A(_15243_),
    .B(_15244_),
    .Y(_15431_));
 sky130_fd_sc_hd__o21ba_2 _37087_ (.A1(_15430_),
    .A2(_15245_),
    .B1_N(_15431_),
    .X(_15432_));
 sky130_fd_sc_hd__nand3b_2 _37088_ (.A_N(_15432_),
    .B(_15095_),
    .C(_15097_),
    .Y(_15433_));
 sky130_fd_sc_hd__o21ai_2 _37089_ (.A1(_15099_),
    .A2(_15100_),
    .B1(_15432_),
    .Y(_15434_));
 sky130_fd_sc_hd__buf_1 _37090_ (.A(_15272_),
    .X(_15435_));
 sky130_fd_sc_hd__a21o_2 _37091_ (.A1(_15433_),
    .A2(_15434_),
    .B1(_15435_),
    .X(_15436_));
 sky130_fd_sc_hd__nand3_2 _37092_ (.A(_15433_),
    .B(_15275_),
    .C(_15434_),
    .Y(_15437_));
 sky130_fd_sc_hd__o21ai_2 _37093_ (.A1(_15271_),
    .A2(_15268_),
    .B1(_15274_),
    .Y(_15438_));
 sky130_fd_sc_hd__a21oi_2 _37094_ (.A1(_15436_),
    .A2(_15437_),
    .B1(_15438_),
    .Y(_15439_));
 sky130_fd_sc_hd__and3_2 _37095_ (.A(_15436_),
    .B(_15437_),
    .C(_15438_),
    .X(_15440_));
 sky130_fd_sc_hd__o21a_2 _37096_ (.A1(_15439_),
    .A2(_15440_),
    .B1(_14653_),
    .X(_15441_));
 sky130_fd_sc_hd__nand2_2 _37097_ (.A(_15257_),
    .B(_15252_),
    .Y(_15442_));
 sky130_fd_sc_hd__nand3_2 _37098_ (.A(_15436_),
    .B(_15437_),
    .C(_15438_),
    .Y(_15443_));
 sky130_fd_sc_hd__nor3b_2 _37099_ (.A(_14652_),
    .B(_15439_),
    .C_N(_15443_),
    .Y(_15444_));
 sky130_vsdinv _37100_ (.A(_15444_),
    .Y(_15445_));
 sky130_fd_sc_hd__nand3b_2 _37101_ (.A_N(_15441_),
    .B(_15442_),
    .C(_15445_),
    .Y(_15446_));
 sky130_fd_sc_hd__o211ai_2 _37102_ (.A1(_15444_),
    .A2(_15441_),
    .B1(_15252_),
    .C1(_15257_),
    .Y(_15447_));
 sky130_fd_sc_hd__nand2_2 _37103_ (.A(_15446_),
    .B(_15447_),
    .Y(_15448_));
 sky130_fd_sc_hd__o21a_2 _37104_ (.A1(_14653_),
    .A2(_15278_),
    .B1(_15279_),
    .X(_15449_));
 sky130_fd_sc_hd__nand2_2 _37105_ (.A(_15448_),
    .B(_15449_),
    .Y(_15450_));
 sky130_fd_sc_hd__nand3b_2 _37106_ (.A_N(_15449_),
    .B(_15446_),
    .C(_15447_),
    .Y(_15451_));
 sky130_fd_sc_hd__nand2_2 _37107_ (.A(_15450_),
    .B(_15451_),
    .Y(_15452_));
 sky130_fd_sc_hd__buf_1 _37108_ (.A(_15452_),
    .X(_15453_));
 sky130_fd_sc_hd__a21boi_2 _37109_ (.A1(_15425_),
    .A2(_15429_),
    .B1_N(_15453_),
    .Y(_15454_));
 sky130_fd_sc_hd__a21oi_2 _37110_ (.A1(_15427_),
    .A2(_15428_),
    .B1(_15424_),
    .Y(_15455_));
 sky130_vsdinv _37111_ (.A(_15429_),
    .Y(_15456_));
 sky130_fd_sc_hd__nor3_2 _37112_ (.A(_15453_),
    .B(_15455_),
    .C(_15456_),
    .Y(_15457_));
 sky130_fd_sc_hd__o21ai_2 _37113_ (.A1(_15291_),
    .A2(_15294_),
    .B1(_15264_),
    .Y(_15458_));
 sky130_fd_sc_hd__o21bai_2 _37114_ (.A1(_15454_),
    .A2(_15457_),
    .B1_N(_15458_),
    .Y(_15459_));
 sky130_fd_sc_hd__o21ai_2 _37115_ (.A1(_15455_),
    .A2(_15456_),
    .B1(_15453_),
    .Y(_15460_));
 sky130_fd_sc_hd__nand3b_2 _37116_ (.A_N(_15452_),
    .B(_15425_),
    .C(_15429_),
    .Y(_15461_));
 sky130_fd_sc_hd__nand3_2 _37117_ (.A(_15460_),
    .B(_15458_),
    .C(_15461_),
    .Y(_15462_));
 sky130_fd_sc_hd__buf_1 _37118_ (.A(_15462_),
    .X(_15463_));
 sky130_fd_sc_hd__a21o_2 _37119_ (.A1(_15290_),
    .A2(_15286_),
    .B1(_15140_),
    .X(_15464_));
 sky130_fd_sc_hd__nand3_2 _37120_ (.A(_15290_),
    .B(_15140_),
    .C(_15286_),
    .Y(_15465_));
 sky130_fd_sc_hd__a21oi_2 _37121_ (.A1(_15464_),
    .A2(_15465_),
    .B1(_15309_),
    .Y(_15466_));
 sky130_vsdinv _37122_ (.A(_15466_),
    .Y(_15467_));
 sky130_fd_sc_hd__nand3_2 _37123_ (.A(_15464_),
    .B(_15307_),
    .C(_15465_),
    .Y(_15468_));
 sky130_fd_sc_hd__nand2_2 _37124_ (.A(_15467_),
    .B(_15468_),
    .Y(_15469_));
 sky130_fd_sc_hd__a21boi_2 _37125_ (.A1(_15459_),
    .A2(_15463_),
    .B1_N(_15469_),
    .Y(_15470_));
 sky130_fd_sc_hd__a21oi_2 _37126_ (.A1(_15460_),
    .A2(_15461_),
    .B1(_15458_),
    .Y(_15471_));
 sky130_fd_sc_hd__nor3b_2 _37127_ (.A(_15469_),
    .B(_15471_),
    .C_N(_15463_),
    .Y(_15472_));
 sky130_fd_sc_hd__o21ai_2 _37128_ (.A1(_15311_),
    .A2(_15314_),
    .B1(_15301_),
    .Y(_15473_));
 sky130_fd_sc_hd__o21bai_2 _37129_ (.A1(_15470_),
    .A2(_15472_),
    .B1_N(_15473_),
    .Y(_15474_));
 sky130_vsdinv _37130_ (.A(_15468_),
    .Y(_15475_));
 sky130_fd_sc_hd__o2bb2ai_2 _37131_ (.A1_N(_15463_),
    .A2_N(_15459_),
    .B1(_15475_),
    .B2(_15466_),
    .Y(_15476_));
 sky130_fd_sc_hd__nand3b_2 _37132_ (.A_N(_15469_),
    .B(_15462_),
    .C(_15459_),
    .Y(_15477_));
 sky130_fd_sc_hd__nand3_2 _37133_ (.A(_15476_),
    .B(_15477_),
    .C(_15473_),
    .Y(_15478_));
 sky130_fd_sc_hd__nand2_2 _37134_ (.A(_15310_),
    .B(_15302_),
    .Y(_15479_));
 sky130_fd_sc_hd__xor2_2 _37135_ (.A(_15160_),
    .B(_15479_),
    .X(_15480_));
 sky130_fd_sc_hd__a21oi_2 _37136_ (.A1(_15474_),
    .A2(_15478_),
    .B1(_15480_),
    .Y(_15481_));
 sky130_vsdinv _37137_ (.A(_15480_),
    .Y(_15482_));
 sky130_fd_sc_hd__a21oi_2 _37138_ (.A1(_15476_),
    .A2(_15477_),
    .B1(_15473_),
    .Y(_15483_));
 sky130_vsdinv _37139_ (.A(_15478_),
    .Y(_15484_));
 sky130_fd_sc_hd__nor3_2 _37140_ (.A(_15482_),
    .B(_15483_),
    .C(_15484_),
    .Y(_15485_));
 sky130_vsdinv _37141_ (.A(_15323_),
    .Y(_15486_));
 sky130_fd_sc_hd__a21oi_2 _37142_ (.A1(_15319_),
    .A2(_15320_),
    .B1(_15317_),
    .Y(_15487_));
 sky130_fd_sc_hd__o21ai_2 _37143_ (.A1(_15486_),
    .A2(_15487_),
    .B1(_15321_),
    .Y(_15488_));
 sky130_fd_sc_hd__o21bai_2 _37144_ (.A1(_15481_),
    .A2(_15485_),
    .B1_N(_15488_),
    .Y(_15489_));
 sky130_fd_sc_hd__o21bai_2 _37145_ (.A1(_15483_),
    .A2(_15484_),
    .B1_N(_15480_),
    .Y(_15490_));
 sky130_fd_sc_hd__nand3_2 _37146_ (.A(_15474_),
    .B(_15480_),
    .C(_15478_),
    .Y(_15491_));
 sky130_fd_sc_hd__nand3_2 _37147_ (.A(_15490_),
    .B(_15488_),
    .C(_15491_),
    .Y(_15492_));
 sky130_fd_sc_hd__buf_1 _37148_ (.A(_15492_),
    .X(_15493_));
 sky130_fd_sc_hd__a21oi_2 _37149_ (.A1(_15147_),
    .A2(_15141_),
    .B1(_14976_),
    .Y(_15494_));
 sky130_fd_sc_hd__a21o_2 _37150_ (.A1(_15489_),
    .A2(_15493_),
    .B1(_15494_),
    .X(_15495_));
 sky130_fd_sc_hd__nand3_2 _37151_ (.A(_15489_),
    .B(_15494_),
    .C(_15492_),
    .Y(_15496_));
 sky130_fd_sc_hd__a21boi_2 _37152_ (.A1(_15154_),
    .A2(_15163_),
    .B1_N(_15159_),
    .Y(_15497_));
 sky130_fd_sc_hd__nor3_2 _37153_ (.A(_15497_),
    .B(_15324_),
    .C(_15326_),
    .Y(_15498_));
 sky130_fd_sc_hd__a21o_2 _37154_ (.A1(_15328_),
    .A2(_15330_),
    .B1(_15498_),
    .X(_15499_));
 sky130_fd_sc_hd__a21oi_2 _37155_ (.A1(_15495_),
    .A2(_15496_),
    .B1(_15499_),
    .Y(_15500_));
 sky130_fd_sc_hd__a21oi_2 _37156_ (.A1(_15489_),
    .A2(_15493_),
    .B1(_15494_),
    .Y(_15501_));
 sky130_fd_sc_hd__a21oi_2 _37157_ (.A1(_15328_),
    .A2(_15330_),
    .B1(_15498_),
    .Y(_15502_));
 sky130_fd_sc_hd__nor3b_2 _37158_ (.A(_15501_),
    .B(_15502_),
    .C_N(_15496_),
    .Y(_15503_));
 sky130_fd_sc_hd__nor2_2 _37159_ (.A(_15500_),
    .B(_15503_),
    .Y(_15504_));
 sky130_fd_sc_hd__o21bai_2 _37160_ (.A1(_15334_),
    .A2(_15341_),
    .B1_N(_15336_),
    .Y(_15505_));
 sky130_fd_sc_hd__xor2_2 _37161_ (.A(_15504_),
    .B(_15505_),
    .X(_02670_));
 sky130_fd_sc_hd__a21oi_2 _37162_ (.A1(_15367_),
    .A2(_15368_),
    .B1(_15364_),
    .Y(_15506_));
 sky130_fd_sc_hd__o21ai_2 _37163_ (.A1(_15383_),
    .A2(_15506_),
    .B1(_15369_),
    .Y(_15507_));
 sky130_fd_sc_hd__and2_2 _37164_ (.A(_18704_),
    .B(_09755_),
    .X(_15508_));
 sky130_fd_sc_hd__buf_1 _37165_ (.A(_15508_),
    .X(_15509_));
 sky130_fd_sc_hd__a22oi_2 _37166_ (.A1(_18696_),
    .A2(_12292_),
    .B1(_12845_),
    .B2(_10673_),
    .Y(_15510_));
 sky130_fd_sc_hd__nand2_2 _37167_ (.A(_12477_),
    .B(_11441_),
    .Y(_15511_));
 sky130_fd_sc_hd__nor3_2 _37168_ (.A(_08314_),
    .B(_16970_),
    .C(_15511_),
    .Y(_15512_));
 sky130_fd_sc_hd__nor2_2 _37169_ (.A(_15510_),
    .B(_15512_),
    .Y(_15513_));
 sky130_fd_sc_hd__xnor2_2 _37170_ (.A(_15509_),
    .B(_15513_),
    .Y(_15514_));
 sky130_vsdinv _37171_ (.A(_15352_),
    .Y(_15515_));
 sky130_fd_sc_hd__a21oi_2 _37172_ (.A1(_15515_),
    .A2(_15351_),
    .B1(_15354_),
    .Y(_15516_));
 sky130_fd_sc_hd__nand2_2 _37173_ (.A(_15514_),
    .B(_15516_),
    .Y(_15517_));
 sky130_fd_sc_hd__buf_1 _37174_ (.A(_15512_),
    .X(_15518_));
 sky130_fd_sc_hd__o21bai_2 _37175_ (.A1(_15510_),
    .A2(_15518_),
    .B1_N(_15509_),
    .Y(_15519_));
 sky130_vsdinv _37176_ (.A(_15510_),
    .Y(_15520_));
 sky130_fd_sc_hd__nand3b_2 _37177_ (.A_N(_15512_),
    .B(_15520_),
    .C(_15509_),
    .Y(_15521_));
 sky130_fd_sc_hd__nand3b_2 _37178_ (.A_N(_15516_),
    .B(_15519_),
    .C(_15521_),
    .Y(_15522_));
 sky130_fd_sc_hd__buf_1 _37179_ (.A(_11736_),
    .X(_15523_));
 sky130_fd_sc_hd__and2_2 _37180_ (.A(_15017_),
    .B(_15523_),
    .X(_15524_));
 sky130_fd_sc_hd__a22oi_2 _37181_ (.A1(_18712_),
    .A2(_12839_),
    .B1(_15199_),
    .B2(_12330_),
    .Y(_15525_));
 sky130_fd_sc_hd__and4_2 _37182_ (.A(_14884_),
    .B(_15020_),
    .C(_10576_),
    .D(_10575_),
    .X(_15526_));
 sky130_fd_sc_hd__nor2_2 _37183_ (.A(_15525_),
    .B(_15526_),
    .Y(_15527_));
 sky130_fd_sc_hd__xor2_2 _37184_ (.A(_15524_),
    .B(_15527_),
    .X(_15528_));
 sky130_fd_sc_hd__a21o_2 _37185_ (.A1(_15517_),
    .A2(_15522_),
    .B1(_15528_),
    .X(_15529_));
 sky130_fd_sc_hd__nand3_2 _37186_ (.A(_15517_),
    .B(_15522_),
    .C(_15528_),
    .Y(_15530_));
 sky130_fd_sc_hd__o21ai_2 _37187_ (.A1(_15347_),
    .A2(_15357_),
    .B1(_15359_),
    .Y(_15531_));
 sky130_fd_sc_hd__a21oi_2 _37188_ (.A1(_15529_),
    .A2(_15530_),
    .B1(_15531_),
    .Y(_15532_));
 sky130_fd_sc_hd__nand3_2 _37189_ (.A(_15529_),
    .B(_15531_),
    .C(_15530_),
    .Y(_15533_));
 sky130_vsdinv _37190_ (.A(_15533_),
    .Y(_15534_));
 sky130_fd_sc_hd__o21a_2 _37191_ (.A1(_15373_),
    .A2(_15374_),
    .B1(_15377_),
    .X(_15535_));
 sky130_fd_sc_hd__nand2_2 _37192_ (.A(_14857_),
    .B(_10042_),
    .Y(_15536_));
 sky130_fd_sc_hd__nand2_2 _37193_ (.A(_18735_),
    .B(_10533_),
    .Y(_15537_));
 sky130_fd_sc_hd__xnor2_2 _37194_ (.A(_15536_),
    .B(_15537_),
    .Y(_15538_));
 sky130_fd_sc_hd__o21ai_2 _37195_ (.A1(_18743_),
    .A2(_19152_),
    .B1(_15538_),
    .Y(_15539_));
 sky130_fd_sc_hd__xor2_2 _37196_ (.A(_15536_),
    .B(_15537_),
    .X(_15540_));
 sky130_fd_sc_hd__nand3_2 _37197_ (.A(_15540_),
    .B(_08459_),
    .C(_13831_),
    .Y(_15541_));
 sky130_fd_sc_hd__a21o_2 _37198_ (.A1(_15345_),
    .A2(_15342_),
    .B1(_15344_),
    .X(_15542_));
 sky130_fd_sc_hd__a21o_2 _37199_ (.A1(_15539_),
    .A2(_15541_),
    .B1(_15542_),
    .X(_15543_));
 sky130_fd_sc_hd__nand3_2 _37200_ (.A(_15542_),
    .B(_15539_),
    .C(_15541_),
    .Y(_15544_));
 sky130_fd_sc_hd__nand2_2 _37201_ (.A(_15543_),
    .B(_15544_),
    .Y(_15545_));
 sky130_fd_sc_hd__xnor2_2 _37202_ (.A(_15535_),
    .B(_15545_),
    .Y(_15546_));
 sky130_fd_sc_hd__o21ai_2 _37203_ (.A1(_15532_),
    .A2(_15534_),
    .B1(_15546_),
    .Y(_15547_));
 sky130_fd_sc_hd__a21o_2 _37204_ (.A1(_15529_),
    .A2(_15530_),
    .B1(_15531_),
    .X(_15548_));
 sky130_fd_sc_hd__nand3b_2 _37205_ (.A_N(_15546_),
    .B(_15548_),
    .C(_15533_),
    .Y(_15549_));
 sky130_fd_sc_hd__nand3_2 _37206_ (.A(_15507_),
    .B(_15547_),
    .C(_15549_),
    .Y(_15550_));
 sky130_fd_sc_hd__a21o_2 _37207_ (.A1(_15547_),
    .A2(_15549_),
    .B1(_15507_),
    .X(_15551_));
 sky130_fd_sc_hd__o21a_2 _37208_ (.A1(_08219_),
    .A2(_10430_),
    .B1(_11204_),
    .X(_15552_));
 sky130_fd_sc_hd__nand3_2 _37209_ (.A(_14648_),
    .B(_12847_),
    .C(_10430_),
    .Y(_15553_));
 sky130_fd_sc_hd__a21oi_2 _37210_ (.A1(_15552_),
    .A2(_15553_),
    .B1(_15242_),
    .Y(_15554_));
 sky130_fd_sc_hd__and3_2 _37211_ (.A(_15552_),
    .B(_15241_),
    .C(_15553_),
    .X(_15555_));
 sky130_fd_sc_hd__nor2_2 _37212_ (.A(_15554_),
    .B(_15555_),
    .Y(_15556_));
 sky130_vsdinv _37213_ (.A(_15556_),
    .Y(_15557_));
 sky130_fd_sc_hd__buf_1 _37214_ (.A(_15057_),
    .X(_15558_));
 sky130_fd_sc_hd__nand3b_2 _37215_ (.A_N(_15395_),
    .B(_18755_),
    .C(_15558_),
    .Y(_15559_));
 sky130_fd_sc_hd__a21boi_2 _37216_ (.A1(_15397_),
    .A2(_15398_),
    .B1_N(_15559_),
    .Y(_15560_));
 sky130_fd_sc_hd__nand2_2 _37217_ (.A(_12527_),
    .B(_09793_),
    .Y(_15561_));
 sky130_fd_sc_hd__nand2_2 _37218_ (.A(_13305_),
    .B(_12871_),
    .Y(_15562_));
 sky130_fd_sc_hd__xor2_2 _37219_ (.A(_15561_),
    .B(_15562_),
    .X(_15563_));
 sky130_fd_sc_hd__nand3_2 _37220_ (.A(_15563_),
    .B(_08086_),
    .C(_19134_),
    .Y(_15564_));
 sky130_fd_sc_hd__xnor2_2 _37221_ (.A(_15561_),
    .B(_15562_),
    .Y(_15565_));
 sky130_fd_sc_hd__o21ai_2 _37222_ (.A1(_08232_),
    .A2(_12389_),
    .B1(_15565_),
    .Y(_15566_));
 sky130_fd_sc_hd__nand2_2 _37223_ (.A(_15564_),
    .B(_15566_),
    .Y(_15567_));
 sky130_fd_sc_hd__xnor2_2 _37224_ (.A(_15560_),
    .B(_15567_),
    .Y(_15568_));
 sky130_fd_sc_hd__nor2_2 _37225_ (.A(_15557_),
    .B(_15568_),
    .Y(_15569_));
 sky130_fd_sc_hd__nand2_2 _37226_ (.A(_15568_),
    .B(_15557_),
    .Y(_15570_));
 sky130_vsdinv _37227_ (.A(_15570_),
    .Y(_15571_));
 sky130_fd_sc_hd__a21bo_2 _37228_ (.A1(_15380_),
    .A2(_15372_),
    .B1_N(_15381_),
    .X(_15572_));
 sky130_fd_sc_hd__o21bai_2 _37229_ (.A1(_15569_),
    .A2(_15571_),
    .B1_N(_15572_),
    .Y(_15573_));
 sky130_fd_sc_hd__o21a_2 _37230_ (.A1(_15409_),
    .A2(_15411_),
    .B1(_15405_),
    .X(_15574_));
 sky130_vsdinv _37231_ (.A(_15574_),
    .Y(_15575_));
 sky130_fd_sc_hd__nand3b_2 _37232_ (.A_N(_15569_),
    .B(_15572_),
    .C(_15570_),
    .Y(_15576_));
 sky130_fd_sc_hd__nand3_2 _37233_ (.A(_15573_),
    .B(_15575_),
    .C(_15576_),
    .Y(_15577_));
 sky130_vsdinv _37234_ (.A(_15577_),
    .Y(_15578_));
 sky130_fd_sc_hd__a21oi_2 _37235_ (.A1(_15573_),
    .A2(_15576_),
    .B1(_15575_),
    .Y(_15579_));
 sky130_fd_sc_hd__o2bb2ai_2 _37236_ (.A1_N(_15550_),
    .A2_N(_15551_),
    .B1(_15578_),
    .B2(_15579_),
    .Y(_15580_));
 sky130_fd_sc_hd__nor2_2 _37237_ (.A(_15579_),
    .B(_15578_),
    .Y(_15581_));
 sky130_fd_sc_hd__nand3_2 _37238_ (.A(_15581_),
    .B(_15551_),
    .C(_15550_),
    .Y(_15582_));
 sky130_fd_sc_hd__o21ai_2 _37239_ (.A1(_15420_),
    .A2(_15422_),
    .B1(_15391_),
    .Y(_15583_));
 sky130_fd_sc_hd__a21oi_2 _37240_ (.A1(_15580_),
    .A2(_15582_),
    .B1(_15583_),
    .Y(_15584_));
 sky130_fd_sc_hd__nand3_2 _37241_ (.A(_15580_),
    .B(_15583_),
    .C(_15582_),
    .Y(_15585_));
 sky130_vsdinv _37242_ (.A(_15585_),
    .Y(_15586_));
 sky130_fd_sc_hd__nor2_2 _37243_ (.A(_15266_),
    .B(_15265_),
    .Y(_15587_));
 sky130_fd_sc_hd__nor2_2 _37244_ (.A(_15406_),
    .B(_15407_),
    .Y(_15588_));
 sky130_fd_sc_hd__o21ba_2 _37245_ (.A1(_15430_),
    .A2(_15408_),
    .B1_N(_15588_),
    .X(_15589_));
 sky130_fd_sc_hd__xnor2_2 _37246_ (.A(_15587_),
    .B(_15589_),
    .Y(_15590_));
 sky130_fd_sc_hd__nand2_2 _37247_ (.A(_15590_),
    .B(_15435_),
    .Y(_15591_));
 sky130_fd_sc_hd__xor2_2 _37248_ (.A(_15587_),
    .B(_15589_),
    .X(_15592_));
 sky130_fd_sc_hd__nand2_2 _37249_ (.A(_15592_),
    .B(_15271_),
    .Y(_15593_));
 sky130_fd_sc_hd__nand2_2 _37250_ (.A(_15437_),
    .B(_15433_),
    .Y(_15594_));
 sky130_fd_sc_hd__a21o_2 _37251_ (.A1(_15591_),
    .A2(_15593_),
    .B1(_15594_),
    .X(_15595_));
 sky130_fd_sc_hd__nand3_2 _37252_ (.A(_15594_),
    .B(_15591_),
    .C(_15593_),
    .Y(_15596_));
 sky130_fd_sc_hd__nand3_2 _37253_ (.A(_15595_),
    .B(_15114_),
    .C(_15596_),
    .Y(_15597_));
 sky130_vsdinv _37254_ (.A(_15597_),
    .Y(_15598_));
 sky130_fd_sc_hd__a21oi_2 _37255_ (.A1(_15595_),
    .A2(_15596_),
    .B1(_15114_),
    .Y(_15599_));
 sky130_fd_sc_hd__nand2_2 _37256_ (.A(_15418_),
    .B(_15413_),
    .Y(_15600_));
 sky130_fd_sc_hd__o21bai_2 _37257_ (.A1(_15598_),
    .A2(_15599_),
    .B1_N(_15600_),
    .Y(_15601_));
 sky130_fd_sc_hd__nand3b_2 _37258_ (.A_N(_15599_),
    .B(_15600_),
    .C(_15597_),
    .Y(_15602_));
 sky130_fd_sc_hd__o21a_2 _37259_ (.A1(_14653_),
    .A2(_15439_),
    .B1(_15443_),
    .X(_15603_));
 sky130_vsdinv _37260_ (.A(_15603_),
    .Y(_15604_));
 sky130_fd_sc_hd__a21o_2 _37261_ (.A1(_15601_),
    .A2(_15602_),
    .B1(_15604_),
    .X(_15605_));
 sky130_fd_sc_hd__nand3_2 _37262_ (.A(_15601_),
    .B(_15604_),
    .C(_15602_),
    .Y(_15606_));
 sky130_fd_sc_hd__nand2_2 _37263_ (.A(_15605_),
    .B(_15606_),
    .Y(_15607_));
 sky130_fd_sc_hd__o21ai_2 _37264_ (.A1(_15584_),
    .A2(_15586_),
    .B1(_15607_),
    .Y(_15608_));
 sky130_fd_sc_hd__a21o_2 _37265_ (.A1(_15580_),
    .A2(_15582_),
    .B1(_15583_),
    .X(_15609_));
 sky130_fd_sc_hd__nand3b_2 _37266_ (.A_N(_15607_),
    .B(_15609_),
    .C(_15585_),
    .Y(_15610_));
 sky130_fd_sc_hd__o21ai_2 _37267_ (.A1(_15453_),
    .A2(_15455_),
    .B1(_15429_),
    .Y(_15611_));
 sky130_fd_sc_hd__a21o_2 _37268_ (.A1(_15608_),
    .A2(_15610_),
    .B1(_15611_),
    .X(_15612_));
 sky130_fd_sc_hd__nand3_2 _37269_ (.A(_15608_),
    .B(_15611_),
    .C(_15610_),
    .Y(_15613_));
 sky130_fd_sc_hd__buf_1 _37270_ (.A(_15613_),
    .X(_15614_));
 sky130_fd_sc_hd__a21o_2 _37271_ (.A1(_15451_),
    .A2(_15446_),
    .B1(_15303_),
    .X(_15615_));
 sky130_fd_sc_hd__nand3_2 _37272_ (.A(_15451_),
    .B(_15303_),
    .C(_15446_),
    .Y(_15616_));
 sky130_fd_sc_hd__nand2_2 _37273_ (.A(_15615_),
    .B(_15616_),
    .Y(_15617_));
 sky130_fd_sc_hd__buf_1 _37274_ (.A(_15305_),
    .X(_15618_));
 sky130_fd_sc_hd__nand2_2 _37275_ (.A(_15617_),
    .B(_15618_),
    .Y(_15619_));
 sky130_fd_sc_hd__nand3_2 _37276_ (.A(_15615_),
    .B(_15616_),
    .C(_15307_),
    .Y(_15620_));
 sky130_fd_sc_hd__nand2_2 _37277_ (.A(_15619_),
    .B(_15620_),
    .Y(_15621_));
 sky130_fd_sc_hd__buf_1 _37278_ (.A(_15621_),
    .X(_15622_));
 sky130_fd_sc_hd__a21boi_2 _37279_ (.A1(_15612_),
    .A2(_15614_),
    .B1_N(_15622_),
    .Y(_15623_));
 sky130_fd_sc_hd__a21oi_2 _37280_ (.A1(_15608_),
    .A2(_15610_),
    .B1(_15611_),
    .Y(_15624_));
 sky130_fd_sc_hd__nor3b_2 _37281_ (.A(_15622_),
    .B(_15624_),
    .C_N(_15614_),
    .Y(_15625_));
 sky130_fd_sc_hd__o21ai_2 _37282_ (.A1(_15469_),
    .A2(_15471_),
    .B1(_15463_),
    .Y(_15626_));
 sky130_fd_sc_hd__o21bai_2 _37283_ (.A1(_15623_),
    .A2(_15625_),
    .B1_N(_15626_),
    .Y(_15627_));
 sky130_vsdinv _37284_ (.A(_15613_),
    .Y(_15628_));
 sky130_fd_sc_hd__o21ai_2 _37285_ (.A1(_15624_),
    .A2(_15628_),
    .B1(_15622_),
    .Y(_15629_));
 sky130_fd_sc_hd__nand3b_2 _37286_ (.A_N(_15621_),
    .B(_15612_),
    .C(_15614_),
    .Y(_15630_));
 sky130_fd_sc_hd__nand3_2 _37287_ (.A(_15629_),
    .B(_15626_),
    .C(_15630_),
    .Y(_15631_));
 sky130_fd_sc_hd__buf_1 _37288_ (.A(_15306_),
    .X(_15632_));
 sky130_fd_sc_hd__buf_1 _37289_ (.A(_15632_),
    .X(_15633_));
 sky130_fd_sc_hd__a21boi_2 _37290_ (.A1(_15633_),
    .A2(_15465_),
    .B1_N(_15464_),
    .Y(_15634_));
 sky130_fd_sc_hd__xor2_2 _37291_ (.A(_13467_),
    .B(_15634_),
    .X(_15635_));
 sky130_fd_sc_hd__a21oi_2 _37292_ (.A1(_15627_),
    .A2(_15631_),
    .B1(_15635_),
    .Y(_15636_));
 sky130_vsdinv _37293_ (.A(_15635_),
    .Y(_15637_));
 sky130_fd_sc_hd__a21oi_2 _37294_ (.A1(_15629_),
    .A2(_15630_),
    .B1(_15626_),
    .Y(_15638_));
 sky130_vsdinv _37295_ (.A(_15631_),
    .Y(_15639_));
 sky130_fd_sc_hd__nor3_2 _37296_ (.A(_15637_),
    .B(_15638_),
    .C(_15639_),
    .Y(_15640_));
 sky130_fd_sc_hd__o21ai_2 _37297_ (.A1(_15482_),
    .A2(_15483_),
    .B1(_15478_),
    .Y(_15641_));
 sky130_fd_sc_hd__o21bai_2 _37298_ (.A1(_15636_),
    .A2(_15640_),
    .B1_N(_15641_),
    .Y(_15642_));
 sky130_fd_sc_hd__o21bai_2 _37299_ (.A1(_15638_),
    .A2(_15639_),
    .B1_N(_15635_),
    .Y(_15643_));
 sky130_fd_sc_hd__nand3_2 _37300_ (.A(_15627_),
    .B(_15635_),
    .C(_15631_),
    .Y(_15644_));
 sky130_fd_sc_hd__nand3_2 _37301_ (.A(_15643_),
    .B(_15641_),
    .C(_15644_),
    .Y(_15645_));
 sky130_fd_sc_hd__a21oi_2 _37302_ (.A1(_15310_),
    .A2(_15302_),
    .B1(_15181_),
    .Y(_15646_));
 sky130_fd_sc_hd__a21oi_2 _37303_ (.A1(_15642_),
    .A2(_15645_),
    .B1(_15646_),
    .Y(_15647_));
 sky130_fd_sc_hd__nand3_2 _37304_ (.A(_15642_),
    .B(_15646_),
    .C(_15645_),
    .Y(_15648_));
 sky130_vsdinv _37305_ (.A(_15648_),
    .Y(_15649_));
 sky130_fd_sc_hd__a21boi_2 _37306_ (.A1(_15489_),
    .A2(_15494_),
    .B1_N(_15493_),
    .Y(_15650_));
 sky130_fd_sc_hd__o21ai_2 _37307_ (.A1(_15647_),
    .A2(_15649_),
    .B1(_15650_),
    .Y(_15651_));
 sky130_fd_sc_hd__nand2_2 _37308_ (.A(_15496_),
    .B(_15493_),
    .Y(_15652_));
 sky130_fd_sc_hd__a21o_2 _37309_ (.A1(_15642_),
    .A2(_15645_),
    .B1(_15646_),
    .X(_15653_));
 sky130_fd_sc_hd__nand3_2 _37310_ (.A(_15652_),
    .B(_15653_),
    .C(_15648_),
    .Y(_15654_));
 sky130_fd_sc_hd__nand2_2 _37311_ (.A(_15651_),
    .B(_15654_),
    .Y(_15655_));
 sky130_fd_sc_hd__nand3_2 _37312_ (.A(_15338_),
    .B(_15337_),
    .C(_15504_),
    .Y(_15656_));
 sky130_vsdinv _37313_ (.A(_15656_),
    .Y(_15657_));
 sky130_fd_sc_hd__nand3_2 _37314_ (.A(_15499_),
    .B(_15495_),
    .C(_15496_),
    .Y(_15658_));
 sky130_fd_sc_hd__o21ai_2 _37315_ (.A1(_15335_),
    .A2(_15500_),
    .B1(_15658_),
    .Y(_15659_));
 sky130_fd_sc_hd__a31oi_2 _37316_ (.A1(_15337_),
    .A2(_15504_),
    .A3(_15340_),
    .B1(_15659_),
    .Y(_15660_));
 sky130_fd_sc_hd__a21boi_2 _37317_ (.A1(_15004_),
    .A2(_15657_),
    .B1_N(_15660_),
    .Y(_15661_));
 sky130_fd_sc_hd__xor2_2 _37318_ (.A(_15655_),
    .B(_15661_),
    .X(_02671_));
 sky130_fd_sc_hd__nor3b_2 _37319_ (.A(_15510_),
    .B(_15518_),
    .C_N(_15508_),
    .Y(_15662_));
 sky130_fd_sc_hd__and2_2 _37320_ (.A(_10484_),
    .B(_08830_),
    .X(_15663_));
 sky130_fd_sc_hd__buf_1 _37321_ (.A(_15663_),
    .X(_15664_));
 sky130_fd_sc_hd__a22oi_2 _37322_ (.A1(_12477_),
    .A2(_09104_),
    .B1(_19191_),
    .B2(_14411_),
    .Y(_15665_));
 sky130_fd_sc_hd__and4_2 _37323_ (.A(_19191_),
    .B(_11322_),
    .C(_14871_),
    .D(_10070_),
    .X(_15666_));
 sky130_fd_sc_hd__nor2_2 _37324_ (.A(_15665_),
    .B(_15666_),
    .Y(_15667_));
 sky130_fd_sc_hd__xor2_2 _37325_ (.A(_15664_),
    .B(_15667_),
    .X(_15668_));
 sky130_fd_sc_hd__o21ai_2 _37326_ (.A1(_15518_),
    .A2(_15662_),
    .B1(_15668_),
    .Y(_15669_));
 sky130_fd_sc_hd__xnor2_2 _37327_ (.A(_15664_),
    .B(_15667_),
    .Y(_15670_));
 sky130_fd_sc_hd__a21oi_2 _37328_ (.A1(_15520_),
    .A2(_15509_),
    .B1(_15518_),
    .Y(_15671_));
 sky130_fd_sc_hd__nand2_2 _37329_ (.A(_15670_),
    .B(_15671_),
    .Y(_15672_));
 sky130_fd_sc_hd__and2_2 _37330_ (.A(_15017_),
    .B(_12596_),
    .X(_15673_));
 sky130_fd_sc_hd__a22oi_2 _37331_ (.A1(_15019_),
    .A2(_10583_),
    .B1(_15021_),
    .B2(_15523_),
    .Y(_15674_));
 sky130_fd_sc_hd__and4_2 _37332_ (.A(_15023_),
    .B(_15020_),
    .C(_10844_),
    .D(_10576_),
    .X(_15675_));
 sky130_fd_sc_hd__nor2_2 _37333_ (.A(_15674_),
    .B(_15675_),
    .Y(_15676_));
 sky130_fd_sc_hd__xor2_2 _37334_ (.A(_15673_),
    .B(_15676_),
    .X(_15677_));
 sky130_fd_sc_hd__a21o_2 _37335_ (.A1(_15669_),
    .A2(_15672_),
    .B1(_15677_),
    .X(_15678_));
 sky130_fd_sc_hd__nand3_2 _37336_ (.A(_15669_),
    .B(_15672_),
    .C(_15677_),
    .Y(_15679_));
 sky130_fd_sc_hd__nand2_2 _37337_ (.A(_15530_),
    .B(_15522_),
    .Y(_15680_));
 sky130_fd_sc_hd__a21oi_2 _37338_ (.A1(_15678_),
    .A2(_15679_),
    .B1(_15680_),
    .Y(_15681_));
 sky130_fd_sc_hd__nand3_2 _37339_ (.A(_15678_),
    .B(_15679_),
    .C(_15680_),
    .Y(_15682_));
 sky130_vsdinv _37340_ (.A(_15682_),
    .Y(_15683_));
 sky130_fd_sc_hd__o21a_2 _37341_ (.A1(_15536_),
    .A2(_15537_),
    .B1(_15541_),
    .X(_15684_));
 sky130_vsdinv _37342_ (.A(_15684_),
    .Y(_15685_));
 sky130_fd_sc_hd__nand2_2 _37343_ (.A(_12500_),
    .B(_12035_),
    .Y(_15686_));
 sky130_fd_sc_hd__nand2_2 _37344_ (.A(_12217_),
    .B(_13830_),
    .Y(_15687_));
 sky130_fd_sc_hd__xnor2_2 _37345_ (.A(_15686_),
    .B(_15687_),
    .Y(_15688_));
 sky130_fd_sc_hd__buf_1 _37346_ (.A(_15558_),
    .X(_15689_));
 sky130_fd_sc_hd__nand3b_2 _37347_ (.A_N(_15688_),
    .B(_08460_),
    .C(_15689_),
    .Y(_15690_));
 sky130_fd_sc_hd__o21ai_2 _37348_ (.A1(_18743_),
    .A2(_19146_),
    .B1(_15688_),
    .Y(_15691_));
 sky130_fd_sc_hd__a21o_2 _37349_ (.A1(_15527_),
    .A2(_15524_),
    .B1(_15526_),
    .X(_15692_));
 sky130_fd_sc_hd__a21o_2 _37350_ (.A1(_15690_),
    .A2(_15691_),
    .B1(_15692_),
    .X(_15693_));
 sky130_fd_sc_hd__nand3_2 _37351_ (.A(_15692_),
    .B(_15690_),
    .C(_15691_),
    .Y(_15694_));
 sky130_fd_sc_hd__nand2_2 _37352_ (.A(_15693_),
    .B(_15694_),
    .Y(_15695_));
 sky130_fd_sc_hd__xor2_2 _37353_ (.A(_15685_),
    .B(_15695_),
    .X(_15696_));
 sky130_fd_sc_hd__o21ai_2 _37354_ (.A1(_15681_),
    .A2(_15683_),
    .B1(_15696_),
    .Y(_15697_));
 sky130_fd_sc_hd__a21o_2 _37355_ (.A1(_15678_),
    .A2(_15679_),
    .B1(_15680_),
    .X(_15698_));
 sky130_fd_sc_hd__nand3b_2 _37356_ (.A_N(_15696_),
    .B(_15698_),
    .C(_15682_),
    .Y(_15699_));
 sky130_fd_sc_hd__o21ai_2 _37357_ (.A1(_15532_),
    .A2(_15546_),
    .B1(_15533_),
    .Y(_15700_));
 sky130_fd_sc_hd__a21oi_2 _37358_ (.A1(_15697_),
    .A2(_15699_),
    .B1(_15700_),
    .Y(_15701_));
 sky130_fd_sc_hd__nand3_2 _37359_ (.A(_15697_),
    .B(_15700_),
    .C(_15699_),
    .Y(_15702_));
 sky130_vsdinv _37360_ (.A(_15702_),
    .Y(_15703_));
 sky130_fd_sc_hd__nand3b_2 _37361_ (.A_N(_15535_),
    .B(_15543_),
    .C(_15544_),
    .Y(_15704_));
 sky130_fd_sc_hd__nand3b_2 _37362_ (.A_N(_15561_),
    .B(_18756_),
    .C(_10914_),
    .Y(_15705_));
 sky130_fd_sc_hd__nand2_2 _37363_ (.A(_15564_),
    .B(_15705_),
    .Y(_15706_));
 sky130_fd_sc_hd__nand2_2 _37364_ (.A(_10417_),
    .B(_11198_),
    .Y(_15707_));
 sky130_fd_sc_hd__nand2_2 _37365_ (.A(_12794_),
    .B(_10540_),
    .Y(_15708_));
 sky130_fd_sc_hd__xnor2_2 _37366_ (.A(_15707_),
    .B(_15708_),
    .Y(_15709_));
 sky130_fd_sc_hd__and2_2 _37367_ (.A(_11204_),
    .B(_08085_),
    .X(_15710_));
 sky130_vsdinv _37368_ (.A(_15710_),
    .Y(_15711_));
 sky130_fd_sc_hd__nand2_2 _37369_ (.A(_15709_),
    .B(_15711_),
    .Y(_15712_));
 sky130_fd_sc_hd__xor2_2 _37370_ (.A(_15707_),
    .B(_15708_),
    .X(_15713_));
 sky130_fd_sc_hd__nand2_2 _37371_ (.A(_15713_),
    .B(_15710_),
    .Y(_15714_));
 sky130_fd_sc_hd__nand3_2 _37372_ (.A(_15706_),
    .B(_15712_),
    .C(_15714_),
    .Y(_15715_));
 sky130_fd_sc_hd__nand2_2 _37373_ (.A(_15714_),
    .B(_15712_),
    .Y(_15716_));
 sky130_fd_sc_hd__nand3_2 _37374_ (.A(_15716_),
    .B(_15705_),
    .C(_15564_),
    .Y(_15717_));
 sky130_fd_sc_hd__buf_1 _37375_ (.A(_15556_),
    .X(_15718_));
 sky130_fd_sc_hd__a21oi_2 _37376_ (.A1(_15715_),
    .A2(_15717_),
    .B1(_15718_),
    .Y(_15719_));
 sky130_fd_sc_hd__buf_1 _37377_ (.A(_15556_),
    .X(_15720_));
 sky130_fd_sc_hd__and3_2 _37378_ (.A(_15717_),
    .B(_15715_),
    .C(_15720_),
    .X(_15721_));
 sky130_fd_sc_hd__a211o_2 _37379_ (.A1(_15704_),
    .A2(_15544_),
    .B1(_15719_),
    .C1(_15721_),
    .X(_15722_));
 sky130_fd_sc_hd__o211ai_2 _37380_ (.A1(_15719_),
    .A2(_15721_),
    .B1(_15544_),
    .C1(_15704_),
    .Y(_15723_));
 sky130_fd_sc_hd__nand3b_2 _37381_ (.A_N(_15560_),
    .B(_15566_),
    .C(_15564_),
    .Y(_15724_));
 sky130_fd_sc_hd__o21a_2 _37382_ (.A1(_15557_),
    .A2(_15568_),
    .B1(_15724_),
    .X(_15725_));
 sky130_fd_sc_hd__a21bo_2 _37383_ (.A1(_15722_),
    .A2(_15723_),
    .B1_N(_15725_),
    .X(_15726_));
 sky130_fd_sc_hd__nand3b_2 _37384_ (.A_N(_15725_),
    .B(_15722_),
    .C(_15723_),
    .Y(_15727_));
 sky130_fd_sc_hd__nand2_2 _37385_ (.A(_15726_),
    .B(_15727_),
    .Y(_15728_));
 sky130_fd_sc_hd__o21ai_2 _37386_ (.A1(_15701_),
    .A2(_15703_),
    .B1(_15728_),
    .Y(_15729_));
 sky130_fd_sc_hd__a21o_2 _37387_ (.A1(_15697_),
    .A2(_15699_),
    .B1(_15700_),
    .X(_15730_));
 sky130_fd_sc_hd__nand3b_2 _37388_ (.A_N(_15728_),
    .B(_15730_),
    .C(_15702_),
    .Y(_15731_));
 sky130_fd_sc_hd__and3_2 _37389_ (.A(_15507_),
    .B(_15547_),
    .C(_15549_),
    .X(_15732_));
 sky130_fd_sc_hd__a21o_2 _37390_ (.A1(_15581_),
    .A2(_15551_),
    .B1(_15732_),
    .X(_15733_));
 sky130_fd_sc_hd__a21o_2 _37391_ (.A1(_15729_),
    .A2(_15731_),
    .B1(_15733_),
    .X(_15734_));
 sky130_fd_sc_hd__nand3_2 _37392_ (.A(_15733_),
    .B(_15729_),
    .C(_15731_),
    .Y(_15735_));
 sky130_vsdinv _37393_ (.A(_15553_),
    .Y(_15736_));
 sky130_fd_sc_hd__a21oi_2 _37394_ (.A1(_15552_),
    .A2(_15242_),
    .B1(_15736_),
    .Y(_15737_));
 sky130_fd_sc_hd__o21a_2 _37395_ (.A1(_15266_),
    .A2(_15265_),
    .B1(_15737_),
    .X(_15738_));
 sky130_fd_sc_hd__nor3_2 _37396_ (.A(_15266_),
    .B(_15737_),
    .C(_15265_),
    .Y(_15739_));
 sky130_vsdinv _37397_ (.A(_15739_),
    .Y(_15740_));
 sky130_fd_sc_hd__nand3b_2 _37398_ (.A_N(_15738_),
    .B(_15740_),
    .C(_15275_),
    .Y(_15741_));
 sky130_fd_sc_hd__o21bai_2 _37399_ (.A1(_15739_),
    .A2(_15738_),
    .B1_N(_15275_),
    .Y(_15742_));
 sky130_fd_sc_hd__nor3_2 _37400_ (.A(_15099_),
    .B(_15100_),
    .C(_15589_),
    .Y(_15743_));
 sky130_fd_sc_hd__a221oi_2 _37401_ (.A1(_15741_),
    .A2(_15742_),
    .B1(_15590_),
    .B2(_15435_),
    .C1(_15743_),
    .Y(_15744_));
 sky130_vsdinv _37402_ (.A(_15744_),
    .Y(_15745_));
 sky130_fd_sc_hd__nor2_2 _37403_ (.A(_15271_),
    .B(_15592_),
    .Y(_15746_));
 sky130_fd_sc_hd__o211ai_2 _37404_ (.A1(_15743_),
    .A2(_15746_),
    .B1(_15741_),
    .C1(_15742_),
    .Y(_15747_));
 sky130_fd_sc_hd__a21oi_2 _37405_ (.A1(_15745_),
    .A2(_15747_),
    .B1(_14843_),
    .Y(_15748_));
 sky130_fd_sc_hd__nand3b_2 _37406_ (.A_N(_15744_),
    .B(_14656_),
    .C(_15747_),
    .Y(_15749_));
 sky130_vsdinv _37407_ (.A(_15749_),
    .Y(_15750_));
 sky130_fd_sc_hd__nand2_2 _37408_ (.A(_15577_),
    .B(_15576_),
    .Y(_15751_));
 sky130_fd_sc_hd__o21bai_2 _37409_ (.A1(_15748_),
    .A2(_15750_),
    .B1_N(_15751_),
    .Y(_15752_));
 sky130_fd_sc_hd__nand3b_2 _37410_ (.A_N(_15748_),
    .B(_15751_),
    .C(_15749_),
    .Y(_15753_));
 sky130_fd_sc_hd__a21boi_2 _37411_ (.A1(_15595_),
    .A2(_14849_),
    .B1_N(_15596_),
    .Y(_15754_));
 sky130_vsdinv _37412_ (.A(_15754_),
    .Y(_15755_));
 sky130_fd_sc_hd__a21o_2 _37413_ (.A1(_15752_),
    .A2(_15753_),
    .B1(_15755_),
    .X(_15756_));
 sky130_fd_sc_hd__nand3b_2 _37414_ (.A_N(_15754_),
    .B(_15752_),
    .C(_15753_),
    .Y(_15757_));
 sky130_fd_sc_hd__nand2_2 _37415_ (.A(_15756_),
    .B(_15757_),
    .Y(_15758_));
 sky130_fd_sc_hd__buf_1 _37416_ (.A(_15758_),
    .X(_15759_));
 sky130_fd_sc_hd__a21boi_2 _37417_ (.A1(_15734_),
    .A2(_15735_),
    .B1_N(_15759_),
    .Y(_15760_));
 sky130_fd_sc_hd__a21oi_2 _37418_ (.A1(_15729_),
    .A2(_15731_),
    .B1(_15733_),
    .Y(_15761_));
 sky130_vsdinv _37419_ (.A(_15735_),
    .Y(_15762_));
 sky130_fd_sc_hd__nor3_2 _37420_ (.A(_15761_),
    .B(_15759_),
    .C(_15762_),
    .Y(_15763_));
 sky130_fd_sc_hd__o21ai_2 _37421_ (.A1(_15607_),
    .A2(_15584_),
    .B1(_15585_),
    .Y(_15764_));
 sky130_fd_sc_hd__o21bai_2 _37422_ (.A1(_15760_),
    .A2(_15763_),
    .B1_N(_15764_),
    .Y(_15765_));
 sky130_fd_sc_hd__o21ai_2 _37423_ (.A1(_15761_),
    .A2(_15762_),
    .B1(_15759_),
    .Y(_15766_));
 sky130_fd_sc_hd__nand3b_2 _37424_ (.A_N(_15758_),
    .B(_15734_),
    .C(_15735_),
    .Y(_15767_));
 sky130_fd_sc_hd__nand3_2 _37425_ (.A(_15766_),
    .B(_15764_),
    .C(_15767_),
    .Y(_15768_));
 sky130_fd_sc_hd__buf_1 _37426_ (.A(_15768_),
    .X(_15769_));
 sky130_fd_sc_hd__a21o_2 _37427_ (.A1(_15606_),
    .A2(_15602_),
    .B1(_15142_),
    .X(_15770_));
 sky130_fd_sc_hd__nand3_2 _37428_ (.A(_15606_),
    .B(_15303_),
    .C(_15602_),
    .Y(_15771_));
 sky130_fd_sc_hd__a21oi_2 _37429_ (.A1(_15770_),
    .A2(_15771_),
    .B1(_15307_),
    .Y(_15772_));
 sky130_fd_sc_hd__nand3_2 _37430_ (.A(_15770_),
    .B(_15632_),
    .C(_15771_),
    .Y(_15773_));
 sky130_fd_sc_hd__or2b_2 _37431_ (.A(_15772_),
    .B_N(_15773_),
    .X(_15774_));
 sky130_fd_sc_hd__a21boi_2 _37432_ (.A1(_15765_),
    .A2(_15769_),
    .B1_N(_15774_),
    .Y(_15775_));
 sky130_fd_sc_hd__a21oi_2 _37433_ (.A1(_15766_),
    .A2(_15767_),
    .B1(_15764_),
    .Y(_15776_));
 sky130_fd_sc_hd__nor3b_2 _37434_ (.A(_15774_),
    .B(_15776_),
    .C_N(_15769_),
    .Y(_15777_));
 sky130_fd_sc_hd__o21ai_2 _37435_ (.A1(_15622_),
    .A2(_15624_),
    .B1(_15614_),
    .Y(_15778_));
 sky130_fd_sc_hd__o21bai_2 _37436_ (.A1(_15775_),
    .A2(_15777_),
    .B1_N(_15778_),
    .Y(_15779_));
 sky130_vsdinv _37437_ (.A(_15773_),
    .Y(_15780_));
 sky130_fd_sc_hd__o2bb2ai_2 _37438_ (.A1_N(_15769_),
    .A2_N(_15765_),
    .B1(_15780_),
    .B2(_15772_),
    .Y(_15781_));
 sky130_fd_sc_hd__nand3b_2 _37439_ (.A_N(_15774_),
    .B(_15765_),
    .C(_15769_),
    .Y(_15782_));
 sky130_fd_sc_hd__nand3_2 _37440_ (.A(_15781_),
    .B(_15778_),
    .C(_15782_),
    .Y(_15783_));
 sky130_fd_sc_hd__a21boi_2 _37441_ (.A1(_15632_),
    .A2(_15616_),
    .B1_N(_15615_),
    .Y(_15784_));
 sky130_fd_sc_hd__xor2_2 _37442_ (.A(_13467_),
    .B(_15784_),
    .X(_15785_));
 sky130_fd_sc_hd__a21o_2 _37443_ (.A1(_15779_),
    .A2(_15783_),
    .B1(_15785_),
    .X(_15786_));
 sky130_fd_sc_hd__o21ai_2 _37444_ (.A1(_15637_),
    .A2(_15638_),
    .B1(_15631_),
    .Y(_15787_));
 sky130_fd_sc_hd__nand3_2 _37445_ (.A(_15779_),
    .B(_15783_),
    .C(_15785_),
    .Y(_15788_));
 sky130_fd_sc_hd__nand3_2 _37446_ (.A(_15786_),
    .B(_15787_),
    .C(_15788_),
    .Y(_15789_));
 sky130_fd_sc_hd__a21oi_2 _37447_ (.A1(_15779_),
    .A2(_15783_),
    .B1(_15785_),
    .Y(_15790_));
 sky130_vsdinv _37448_ (.A(_15788_),
    .Y(_15791_));
 sky130_fd_sc_hd__o21bai_2 _37449_ (.A1(_15790_),
    .A2(_15791_),
    .B1_N(_15787_),
    .Y(_15792_));
 sky130_fd_sc_hd__buf_1 _37450_ (.A(_14976_),
    .X(_15793_));
 sky130_fd_sc_hd__buf_1 _37451_ (.A(_15793_),
    .X(_15794_));
 sky130_fd_sc_hd__o2bb2ai_2 _37452_ (.A1_N(_15789_),
    .A2_N(_15792_),
    .B1(_15794_),
    .B2(_15634_),
    .Y(_15795_));
 sky130_fd_sc_hd__a21oi_2 _37453_ (.A1(_15468_),
    .A2(_15464_),
    .B1(_15793_),
    .Y(_15796_));
 sky130_fd_sc_hd__nand3_2 _37454_ (.A(_15792_),
    .B(_15796_),
    .C(_15789_),
    .Y(_15797_));
 sky130_fd_sc_hd__a21boi_2 _37455_ (.A1(_15642_),
    .A2(_15646_),
    .B1_N(_15645_),
    .Y(_15798_));
 sky130_fd_sc_hd__a21boi_2 _37456_ (.A1(_15795_),
    .A2(_15797_),
    .B1_N(_15798_),
    .Y(_15799_));
 sky130_fd_sc_hd__a21oi_2 _37457_ (.A1(_15792_),
    .A2(_15789_),
    .B1(_15796_),
    .Y(_15800_));
 sky130_fd_sc_hd__nor3b_2 _37458_ (.A(_15798_),
    .B(_15800_),
    .C_N(_15797_),
    .Y(_15801_));
 sky130_fd_sc_hd__nor2_2 _37459_ (.A(_15799_),
    .B(_15801_),
    .Y(_15802_));
 sky130_fd_sc_hd__o21a_2 _37460_ (.A1(_15655_),
    .A2(_15661_),
    .B1(_15654_),
    .X(_15803_));
 sky130_fd_sc_hd__xnor2_2 _37461_ (.A(_15802_),
    .B(_15803_),
    .Y(_02672_));
 sky130_vsdinv _37462_ (.A(_15665_),
    .Y(_15804_));
 sky130_fd_sc_hd__a21oi_2 _37463_ (.A1(_15804_),
    .A2(_15664_),
    .B1(_15666_),
    .Y(_15805_));
 sky130_vsdinv _37464_ (.A(_15805_),
    .Y(_15806_));
 sky130_fd_sc_hd__and2_2 _37465_ (.A(_18705_),
    .B(_10583_),
    .X(_15807_));
 sky130_fd_sc_hd__a22oi_2 _37466_ (.A1(_12477_),
    .A2(_10575_),
    .B1(_19186_),
    .B2(_10673_),
    .Y(_15808_));
 sky130_fd_sc_hd__nand2_2 _37467_ (.A(_10482_),
    .B(_10077_),
    .Y(_15809_));
 sky130_fd_sc_hd__nor3_2 _37468_ (.A(_08827_),
    .B(_16970_),
    .C(_15809_),
    .Y(_15810_));
 sky130_fd_sc_hd__nor2_2 _37469_ (.A(_15808_),
    .B(_15810_),
    .Y(_15811_));
 sky130_fd_sc_hd__xor2_2 _37470_ (.A(_15807_),
    .B(_15811_),
    .X(_15812_));
 sky130_fd_sc_hd__nor2_2 _37471_ (.A(_15806_),
    .B(_15812_),
    .Y(_15813_));
 sky130_fd_sc_hd__nand2_2 _37472_ (.A(_15812_),
    .B(_15806_),
    .Y(_15814_));
 sky130_vsdinv _37473_ (.A(_15814_),
    .Y(_15815_));
 sky130_fd_sc_hd__and2_2 _37474_ (.A(_15017_),
    .B(_13580_),
    .X(_15816_));
 sky130_fd_sc_hd__a22oi_2 _37475_ (.A1(_15019_),
    .A2(_15523_),
    .B1(_15021_),
    .B2(_10043_),
    .Y(_15817_));
 sky130_fd_sc_hd__and4_2 _37476_ (.A(_15023_),
    .B(_18718_),
    .C(_10849_),
    .D(_10844_),
    .X(_15818_));
 sky130_fd_sc_hd__nor2_2 _37477_ (.A(_15817_),
    .B(_15818_),
    .Y(_15819_));
 sky130_fd_sc_hd__xor2_2 _37478_ (.A(_15816_),
    .B(_15819_),
    .X(_15820_));
 sky130_fd_sc_hd__o21bai_2 _37479_ (.A1(_15813_),
    .A2(_15815_),
    .B1_N(_15820_),
    .Y(_15821_));
 sky130_fd_sc_hd__nand3b_2 _37480_ (.A_N(_15813_),
    .B(_15814_),
    .C(_15820_),
    .Y(_15822_));
 sky130_fd_sc_hd__nand2_2 _37481_ (.A(_15679_),
    .B(_15669_),
    .Y(_15823_));
 sky130_fd_sc_hd__a21oi_2 _37482_ (.A1(_15821_),
    .A2(_15822_),
    .B1(_15823_),
    .Y(_15824_));
 sky130_fd_sc_hd__nand3_2 _37483_ (.A(_15823_),
    .B(_15821_),
    .C(_15822_),
    .Y(_15825_));
 sky130_vsdinv _37484_ (.A(_15825_),
    .Y(_15826_));
 sky130_fd_sc_hd__buf_1 _37485_ (.A(_13831_),
    .X(_15827_));
 sky130_fd_sc_hd__nand3b_2 _37486_ (.A_N(_15686_),
    .B(_18737_),
    .C(_15827_),
    .Y(_15828_));
 sky130_fd_sc_hd__o31a_2 _37487_ (.A1(_18743_),
    .A2(_19147_),
    .A3(_15688_),
    .B1(_15828_),
    .X(_15829_));
 sky130_vsdinv _37488_ (.A(_15829_),
    .Y(_15830_));
 sky130_fd_sc_hd__nand2_2 _37489_ (.A(_18729_),
    .B(_13830_),
    .Y(_15831_));
 sky130_fd_sc_hd__nand2_2 _37490_ (.A(_11042_),
    .B(_15057_),
    .Y(_15832_));
 sky130_fd_sc_hd__xor2_2 _37491_ (.A(_15831_),
    .B(_15832_),
    .X(_15833_));
 sky130_fd_sc_hd__a21o_2 _37492_ (.A1(_15376_),
    .A2(_10915_),
    .B1(_15833_),
    .X(_15834_));
 sky130_fd_sc_hd__nand3_2 _37493_ (.A(_15833_),
    .B(_08460_),
    .C(_10915_),
    .Y(_15835_));
 sky130_fd_sc_hd__a21o_2 _37494_ (.A1(_15676_),
    .A2(_15673_),
    .B1(_15675_),
    .X(_15836_));
 sky130_fd_sc_hd__a21o_2 _37495_ (.A1(_15834_),
    .A2(_15835_),
    .B1(_15836_),
    .X(_15837_));
 sky130_fd_sc_hd__nand3_2 _37496_ (.A(_15836_),
    .B(_15834_),
    .C(_15835_),
    .Y(_15838_));
 sky130_fd_sc_hd__nand2_2 _37497_ (.A(_15837_),
    .B(_15838_),
    .Y(_15839_));
 sky130_fd_sc_hd__xor2_2 _37498_ (.A(_15830_),
    .B(_15839_),
    .X(_15840_));
 sky130_fd_sc_hd__o21ai_2 _37499_ (.A1(_15824_),
    .A2(_15826_),
    .B1(_15840_),
    .Y(_15841_));
 sky130_fd_sc_hd__a21o_2 _37500_ (.A1(_15821_),
    .A2(_15822_),
    .B1(_15823_),
    .X(_15842_));
 sky130_fd_sc_hd__nand3b_2 _37501_ (.A_N(_15840_),
    .B(_15842_),
    .C(_15825_),
    .Y(_15843_));
 sky130_fd_sc_hd__o21ai_2 _37502_ (.A1(_15696_),
    .A2(_15681_),
    .B1(_15682_),
    .Y(_15844_));
 sky130_fd_sc_hd__a21o_2 _37503_ (.A1(_15841_),
    .A2(_15843_),
    .B1(_15844_),
    .X(_15845_));
 sky130_fd_sc_hd__nand3_2 _37504_ (.A(_15841_),
    .B(_15843_),
    .C(_15844_),
    .Y(_15846_));
 sky130_fd_sc_hd__a21boi_2 _37505_ (.A1(_15718_),
    .A2(_15717_),
    .B1_N(_15715_),
    .Y(_15847_));
 sky130_fd_sc_hd__nand2_2 _37506_ (.A(_14245_),
    .B(_12905_),
    .Y(_15848_));
 sky130_fd_sc_hd__nand2_2 _37507_ (.A(_12368_),
    .B(_11968_),
    .Y(_15849_));
 sky130_fd_sc_hd__xnor2_2 _37508_ (.A(_15848_),
    .B(_15849_),
    .Y(_15850_));
 sky130_fd_sc_hd__nand3b_2 _37509_ (.A_N(_15850_),
    .B(_14831_),
    .C(_07847_),
    .Y(_15851_));
 sky130_fd_sc_hd__nand2_2 _37510_ (.A(_15850_),
    .B(_15711_),
    .Y(_15852_));
 sky130_fd_sc_hd__o21ai_2 _37511_ (.A1(_15707_),
    .A2(_15708_),
    .B1(_15714_),
    .Y(_15853_));
 sky130_fd_sc_hd__a21o_2 _37512_ (.A1(_15851_),
    .A2(_15852_),
    .B1(_15853_),
    .X(_15854_));
 sky130_fd_sc_hd__nand3_2 _37513_ (.A(_15853_),
    .B(_15851_),
    .C(_15852_),
    .Y(_15855_));
 sky130_fd_sc_hd__a21o_2 _37514_ (.A1(_15854_),
    .A2(_15855_),
    .B1(_15720_),
    .X(_15856_));
 sky130_fd_sc_hd__nand3_2 _37515_ (.A(_15854_),
    .B(_15720_),
    .C(_15855_),
    .Y(_15857_));
 sky130_fd_sc_hd__a21bo_2 _37516_ (.A1(_15693_),
    .A2(_15685_),
    .B1_N(_15694_),
    .X(_15858_));
 sky130_fd_sc_hd__a21o_2 _37517_ (.A1(_15856_),
    .A2(_15857_),
    .B1(_15858_),
    .X(_15859_));
 sky130_fd_sc_hd__nand3_2 _37518_ (.A(_15858_),
    .B(_15856_),
    .C(_15857_),
    .Y(_15860_));
 sky130_fd_sc_hd__nand2_2 _37519_ (.A(_15859_),
    .B(_15860_),
    .Y(_15861_));
 sky130_fd_sc_hd__xnor2_2 _37520_ (.A(_15847_),
    .B(_15861_),
    .Y(_15862_));
 sky130_fd_sc_hd__buf_1 _37521_ (.A(_15862_),
    .X(_15863_));
 sky130_fd_sc_hd__a21boi_2 _37522_ (.A1(_15845_),
    .A2(_15846_),
    .B1_N(_15863_),
    .Y(_15864_));
 sky130_fd_sc_hd__a21oi_2 _37523_ (.A1(_15841_),
    .A2(_15843_),
    .B1(_15844_),
    .Y(_15865_));
 sky130_vsdinv _37524_ (.A(_15846_),
    .Y(_15866_));
 sky130_fd_sc_hd__nor3_2 _37525_ (.A(_15863_),
    .B(_15865_),
    .C(_15866_),
    .Y(_15867_));
 sky130_fd_sc_hd__o21ai_2 _37526_ (.A1(_15728_),
    .A2(_15701_),
    .B1(_15702_),
    .Y(_15868_));
 sky130_fd_sc_hd__o21bai_2 _37527_ (.A1(_15864_),
    .A2(_15867_),
    .B1_N(_15868_),
    .Y(_15869_));
 sky130_fd_sc_hd__o21ai_2 _37528_ (.A1(_15865_),
    .A2(_15866_),
    .B1(_15863_),
    .Y(_15870_));
 sky130_fd_sc_hd__nand3b_2 _37529_ (.A_N(_15862_),
    .B(_15845_),
    .C(_15846_),
    .Y(_15871_));
 sky130_fd_sc_hd__nand3_2 _37530_ (.A(_15870_),
    .B(_15871_),
    .C(_15868_),
    .Y(_15872_));
 sky130_fd_sc_hd__o2111ai_2 _37531_ (.A1(_16963_),
    .A2(_18782_),
    .B1(_14634_),
    .C1(_14827_),
    .D1(_15737_),
    .Y(_15873_));
 sky130_fd_sc_hd__a21bo_2 _37532_ (.A1(_15739_),
    .A2(_15272_),
    .B1_N(_15873_),
    .X(_15874_));
 sky130_fd_sc_hd__xnor2_2 _37533_ (.A(_15874_),
    .B(_14651_),
    .Y(_15875_));
 sky130_vsdinv _37534_ (.A(_15875_),
    .Y(_15876_));
 sky130_fd_sc_hd__a21o_2 _37535_ (.A1(_15727_),
    .A2(_15722_),
    .B1(_15876_),
    .X(_15877_));
 sky130_fd_sc_hd__buf_1 _37536_ (.A(_15876_),
    .X(_15878_));
 sky130_fd_sc_hd__nand3_2 _37537_ (.A(_15727_),
    .B(_15722_),
    .C(_15878_),
    .Y(_15879_));
 sky130_fd_sc_hd__o211a_2 _37538_ (.A1(_15736_),
    .A2(_15555_),
    .B1(_15435_),
    .C1(_15587_),
    .X(_15880_));
 sky130_fd_sc_hd__a31oi_2 _37539_ (.A1(_15745_),
    .A2(_15747_),
    .A3(_15114_),
    .B1(_15880_),
    .Y(_15881_));
 sky130_fd_sc_hd__a21bo_2 _37540_ (.A1(_15877_),
    .A2(_15879_),
    .B1_N(_15881_),
    .X(_15882_));
 sky130_fd_sc_hd__nand3b_2 _37541_ (.A_N(_15881_),
    .B(_15877_),
    .C(_15879_),
    .Y(_15883_));
 sky130_fd_sc_hd__nand2_2 _37542_ (.A(_15882_),
    .B(_15883_),
    .Y(_15884_));
 sky130_vsdinv _37543_ (.A(_15884_),
    .Y(_15885_));
 sky130_fd_sc_hd__a21oi_2 _37544_ (.A1(_15869_),
    .A2(_15872_),
    .B1(_15885_),
    .Y(_15886_));
 sky130_fd_sc_hd__nand3_2 _37545_ (.A(_15869_),
    .B(_15885_),
    .C(_15872_),
    .Y(_15887_));
 sky130_vsdinv _37546_ (.A(_15887_),
    .Y(_15888_));
 sky130_fd_sc_hd__o21ai_2 _37547_ (.A1(_15761_),
    .A2(_15759_),
    .B1(_15735_),
    .Y(_15889_));
 sky130_fd_sc_hd__o21bai_2 _37548_ (.A1(_15886_),
    .A2(_15888_),
    .B1_N(_15889_),
    .Y(_15890_));
 sky130_fd_sc_hd__a21oi_2 _37549_ (.A1(_15870_),
    .A2(_15871_),
    .B1(_15868_),
    .Y(_15891_));
 sky130_fd_sc_hd__and3_2 _37550_ (.A(_15870_),
    .B(_15871_),
    .C(_15868_),
    .X(_15892_));
 sky130_fd_sc_hd__o21bai_2 _37551_ (.A1(_15891_),
    .A2(_15892_),
    .B1_N(_15885_),
    .Y(_15893_));
 sky130_fd_sc_hd__nand3_2 _37552_ (.A(_15893_),
    .B(_15887_),
    .C(_15889_),
    .Y(_15894_));
 sky130_fd_sc_hd__a21o_2 _37553_ (.A1(_15757_),
    .A2(_15753_),
    .B1(_15140_),
    .X(_15895_));
 sky130_fd_sc_hd__nand3_2 _37554_ (.A(_15757_),
    .B(_15142_),
    .C(_15753_),
    .Y(_15896_));
 sky130_fd_sc_hd__a21o_2 _37555_ (.A1(_15895_),
    .A2(_15896_),
    .B1(_15309_),
    .X(_15897_));
 sky130_fd_sc_hd__nand3_2 _37556_ (.A(_15895_),
    .B(_15309_),
    .C(_15896_),
    .Y(_15898_));
 sky130_fd_sc_hd__nand2_2 _37557_ (.A(_15897_),
    .B(_15898_),
    .Y(_15899_));
 sky130_fd_sc_hd__buf_1 _37558_ (.A(_15899_),
    .X(_15900_));
 sky130_fd_sc_hd__a21boi_2 _37559_ (.A1(_15890_),
    .A2(_15894_),
    .B1_N(_15900_),
    .Y(_15901_));
 sky130_fd_sc_hd__a21oi_2 _37560_ (.A1(_15893_),
    .A2(_15887_),
    .B1(_15889_),
    .Y(_15902_));
 sky130_vsdinv _37561_ (.A(_15894_),
    .Y(_15903_));
 sky130_fd_sc_hd__nor3_2 _37562_ (.A(_15900_),
    .B(_15902_),
    .C(_15903_),
    .Y(_15904_));
 sky130_fd_sc_hd__o21ai_2 _37563_ (.A1(_15774_),
    .A2(_15776_),
    .B1(_15768_),
    .Y(_15905_));
 sky130_fd_sc_hd__o21bai_2 _37564_ (.A1(_15901_),
    .A2(_15904_),
    .B1_N(_15905_),
    .Y(_15906_));
 sky130_fd_sc_hd__o21ai_2 _37565_ (.A1(_15902_),
    .A2(_15903_),
    .B1(_15900_),
    .Y(_15907_));
 sky130_fd_sc_hd__nand3b_2 _37566_ (.A_N(_15899_),
    .B(_15890_),
    .C(_15894_),
    .Y(_15908_));
 sky130_fd_sc_hd__nand3_2 _37567_ (.A(_15907_),
    .B(_15908_),
    .C(_15905_),
    .Y(_15909_));
 sky130_fd_sc_hd__a21boi_2 _37568_ (.A1(_15632_),
    .A2(_15771_),
    .B1_N(_15770_),
    .Y(_15910_));
 sky130_fd_sc_hd__xor2_2 _37569_ (.A(_13467_),
    .B(_15910_),
    .X(_15911_));
 sky130_fd_sc_hd__a21o_2 _37570_ (.A1(_15906_),
    .A2(_15909_),
    .B1(_15911_),
    .X(_15912_));
 sky130_fd_sc_hd__nand3_2 _37571_ (.A(_15906_),
    .B(_15911_),
    .C(_15909_),
    .Y(_15913_));
 sky130_vsdinv _37572_ (.A(_15785_),
    .Y(_15914_));
 sky130_fd_sc_hd__a21oi_2 _37573_ (.A1(_15781_),
    .A2(_15782_),
    .B1(_15778_),
    .Y(_15915_));
 sky130_fd_sc_hd__o21ai_2 _37574_ (.A1(_15914_),
    .A2(_15915_),
    .B1(_15783_),
    .Y(_15916_));
 sky130_fd_sc_hd__nand3_2 _37575_ (.A(_15912_),
    .B(_15913_),
    .C(_15916_),
    .Y(_15917_));
 sky130_fd_sc_hd__buf_1 _37576_ (.A(_15917_),
    .X(_15918_));
 sky130_fd_sc_hd__a21oi_2 _37577_ (.A1(_15906_),
    .A2(_15909_),
    .B1(_15911_),
    .Y(_15919_));
 sky130_vsdinv _37578_ (.A(_15913_),
    .Y(_15920_));
 sky130_fd_sc_hd__o21bai_2 _37579_ (.A1(_15919_),
    .A2(_15920_),
    .B1_N(_15916_),
    .Y(_15921_));
 sky130_fd_sc_hd__buf_1 _37580_ (.A(_15182_),
    .X(_15922_));
 sky130_fd_sc_hd__o2bb2ai_2 _37581_ (.A1_N(_15918_),
    .A2_N(_15921_),
    .B1(_15922_),
    .B2(_15784_),
    .Y(_15923_));
 sky130_fd_sc_hd__a21oi_2 _37582_ (.A1(_15620_),
    .A2(_15615_),
    .B1(_15181_),
    .Y(_15924_));
 sky130_fd_sc_hd__nand3_2 _37583_ (.A(_15921_),
    .B(_15924_),
    .C(_15917_),
    .Y(_15925_));
 sky130_fd_sc_hd__a21boi_2 _37584_ (.A1(_15792_),
    .A2(_15796_),
    .B1_N(_15789_),
    .Y(_15926_));
 sky130_fd_sc_hd__a21boi_2 _37585_ (.A1(_15923_),
    .A2(_15925_),
    .B1_N(_15926_),
    .Y(_15927_));
 sky130_fd_sc_hd__a21oi_2 _37586_ (.A1(_15921_),
    .A2(_15918_),
    .B1(_15924_),
    .Y(_15928_));
 sky130_fd_sc_hd__nor3b_2 _37587_ (.A(_15926_),
    .B(_15928_),
    .C_N(_15925_),
    .Y(_15929_));
 sky130_fd_sc_hd__nor2_2 _37588_ (.A(_15927_),
    .B(_15929_),
    .Y(_15930_));
 sky130_fd_sc_hd__a21bo_2 _37589_ (.A1(_15003_),
    .A2(_15657_),
    .B1_N(_15660_),
    .X(_15931_));
 sky130_fd_sc_hd__nor3_2 _37590_ (.A(_15801_),
    .B(_15799_),
    .C(_15655_),
    .Y(_15932_));
 sky130_fd_sc_hd__nand3b_2 _37591_ (.A_N(_15798_),
    .B(_15797_),
    .C(_15795_),
    .Y(_15933_));
 sky130_fd_sc_hd__a21oi_2 _37592_ (.A1(_15933_),
    .A2(_15654_),
    .B1(_15799_),
    .Y(_15934_));
 sky130_fd_sc_hd__a21o_2 _37593_ (.A1(_15931_),
    .A2(_15932_),
    .B1(_15934_),
    .X(_15935_));
 sky130_fd_sc_hd__xor2_2 _37594_ (.A(_15930_),
    .B(_15935_),
    .X(_02673_));
 sky130_fd_sc_hd__and2_2 _37595_ (.A(_18705_),
    .B(_15523_),
    .X(_15936_));
 sky130_fd_sc_hd__nand2_2 _37596_ (.A(_14871_),
    .B(_12842_),
    .Y(_15937_));
 sky130_fd_sc_hd__nand2_2 _37597_ (.A(_19181_),
    .B(_14411_),
    .Y(_15938_));
 sky130_fd_sc_hd__xor2_2 _37598_ (.A(_15937_),
    .B(_15938_),
    .X(_15939_));
 sky130_fd_sc_hd__xnor2_2 _37599_ (.A(_15936_),
    .B(_15939_),
    .Y(_15940_));
 sky130_vsdinv _37600_ (.A(_15808_),
    .Y(_15941_));
 sky130_fd_sc_hd__a21oi_2 _37601_ (.A1(_15941_),
    .A2(_15807_),
    .B1(_15810_),
    .Y(_15942_));
 sky130_fd_sc_hd__nand2_2 _37602_ (.A(_15940_),
    .B(_15942_),
    .Y(_15943_));
 sky130_fd_sc_hd__xor2_2 _37603_ (.A(_15936_),
    .B(_15939_),
    .X(_15944_));
 sky130_vsdinv _37604_ (.A(_15942_),
    .Y(_15945_));
 sky130_fd_sc_hd__nand2_2 _37605_ (.A(_15944_),
    .B(_15945_),
    .Y(_15946_));
 sky130_fd_sc_hd__and2_2 _37606_ (.A(_14701_),
    .B(_13831_),
    .X(_15947_));
 sky130_fd_sc_hd__a22oi_2 _37607_ (.A1(_15019_),
    .A2(_12596_),
    .B1(_15021_),
    .B2(_13369_),
    .Y(_15948_));
 sky130_fd_sc_hd__and4_2 _37608_ (.A(_18712_),
    .B(_15199_),
    .C(_10052_),
    .D(_09809_),
    .X(_15949_));
 sky130_fd_sc_hd__nor2_2 _37609_ (.A(_15948_),
    .B(_15949_),
    .Y(_15950_));
 sky130_fd_sc_hd__xor2_2 _37610_ (.A(_15947_),
    .B(_15950_),
    .X(_15951_));
 sky130_fd_sc_hd__a21oi_2 _37611_ (.A1(_15943_),
    .A2(_15946_),
    .B1(_15951_),
    .Y(_15952_));
 sky130_fd_sc_hd__nand3_2 _37612_ (.A(_15943_),
    .B(_15946_),
    .C(_15951_),
    .Y(_15953_));
 sky130_vsdinv _37613_ (.A(_15953_),
    .Y(_15954_));
 sky130_vsdinv _37614_ (.A(_15820_),
    .Y(_15955_));
 sky130_fd_sc_hd__o21ai_2 _37615_ (.A1(_15955_),
    .A2(_15813_),
    .B1(_15814_),
    .Y(_15956_));
 sky130_fd_sc_hd__o21bai_2 _37616_ (.A1(_15952_),
    .A2(_15954_),
    .B1_N(_15956_),
    .Y(_15957_));
 sky130_fd_sc_hd__a21o_2 _37617_ (.A1(_15943_),
    .A2(_15946_),
    .B1(_15951_),
    .X(_15958_));
 sky130_fd_sc_hd__nand3_2 _37618_ (.A(_15958_),
    .B(_15953_),
    .C(_15956_),
    .Y(_15959_));
 sky130_fd_sc_hd__o21a_2 _37619_ (.A1(_15831_),
    .A2(_15832_),
    .B1(_15835_),
    .X(_15960_));
 sky130_vsdinv _37620_ (.A(_15960_),
    .Y(_15961_));
 sky130_fd_sc_hd__nand2_2 _37621_ (.A(_18729_),
    .B(_12069_),
    .Y(_15962_));
 sky130_fd_sc_hd__nand2_2 _37622_ (.A(_11042_),
    .B(_10897_),
    .Y(_15963_));
 sky130_fd_sc_hd__xor2_2 _37623_ (.A(_15962_),
    .B(_15963_),
    .X(_15964_));
 sky130_fd_sc_hd__a21o_2 _37624_ (.A1(_15376_),
    .A2(_19135_),
    .B1(_15964_),
    .X(_15965_));
 sky130_fd_sc_hd__nand3_2 _37625_ (.A(_15964_),
    .B(_15376_),
    .C(_19135_),
    .Y(_15966_));
 sky130_fd_sc_hd__a21o_2 _37626_ (.A1(_15819_),
    .A2(_15816_),
    .B1(_15818_),
    .X(_15967_));
 sky130_fd_sc_hd__a21oi_2 _37627_ (.A1(_15965_),
    .A2(_15966_),
    .B1(_15967_),
    .Y(_15968_));
 sky130_fd_sc_hd__nand3_2 _37628_ (.A(_15967_),
    .B(_15965_),
    .C(_15966_),
    .Y(_15969_));
 sky130_vsdinv _37629_ (.A(_15969_),
    .Y(_15970_));
 sky130_fd_sc_hd__nor2_2 _37630_ (.A(_15968_),
    .B(_15970_),
    .Y(_15971_));
 sky130_fd_sc_hd__xor2_2 _37631_ (.A(_15961_),
    .B(_15971_),
    .X(_15972_));
 sky130_fd_sc_hd__a21oi_2 _37632_ (.A1(_15957_),
    .A2(_15959_),
    .B1(_15972_),
    .Y(_15973_));
 sky130_fd_sc_hd__nand3_2 _37633_ (.A(_15972_),
    .B(_15957_),
    .C(_15959_),
    .Y(_15974_));
 sky130_vsdinv _37634_ (.A(_15974_),
    .Y(_15975_));
 sky130_fd_sc_hd__o21ai_2 _37635_ (.A1(_15840_),
    .A2(_15824_),
    .B1(_15825_),
    .Y(_15976_));
 sky130_fd_sc_hd__o21bai_2 _37636_ (.A1(_15973_),
    .A2(_15975_),
    .B1_N(_15976_),
    .Y(_15977_));
 sky130_fd_sc_hd__a21o_2 _37637_ (.A1(_15957_),
    .A2(_15959_),
    .B1(_15972_),
    .X(_15978_));
 sky130_fd_sc_hd__nand3_2 _37638_ (.A(_15978_),
    .B(_15974_),
    .C(_15976_),
    .Y(_15979_));
 sky130_fd_sc_hd__buf_1 _37639_ (.A(_14648_),
    .X(_15980_));
 sky130_fd_sc_hd__buf_1 _37640_ (.A(_15980_),
    .X(_15981_));
 sky130_fd_sc_hd__nand3b_2 _37641_ (.A_N(_15848_),
    .B(_15981_),
    .C(_18756_),
    .Y(_15982_));
 sky130_fd_sc_hd__o21a_2 _37642_ (.A1(_18749_),
    .A2(_10734_),
    .B1(_14830_),
    .X(_15983_));
 sky130_fd_sc_hd__nand3_2 _37643_ (.A(_14830_),
    .B(_18750_),
    .C(_12791_),
    .Y(_15984_));
 sky130_fd_sc_hd__nand2_2 _37644_ (.A(_15983_),
    .B(_15984_),
    .Y(_15985_));
 sky130_fd_sc_hd__xor2_2 _37645_ (.A(_15710_),
    .B(_15985_),
    .X(_15986_));
 sky130_fd_sc_hd__a21bo_2 _37646_ (.A1(_15982_),
    .A2(_15851_),
    .B1_N(_15986_),
    .X(_15987_));
 sky130_fd_sc_hd__nand3b_2 _37647_ (.A_N(_15986_),
    .B(_15982_),
    .C(_15851_),
    .Y(_15988_));
 sky130_fd_sc_hd__nand2_2 _37648_ (.A(_15987_),
    .B(_15988_),
    .Y(_15989_));
 sky130_fd_sc_hd__nand2_2 _37649_ (.A(_15989_),
    .B(_15718_),
    .Y(_15990_));
 sky130_fd_sc_hd__nand3_2 _37650_ (.A(_15987_),
    .B(_15557_),
    .C(_15988_),
    .Y(_15991_));
 sky130_fd_sc_hd__a21boi_2 _37651_ (.A1(_15837_),
    .A2(_15830_),
    .B1_N(_15838_),
    .Y(_15992_));
 sky130_fd_sc_hd__a21bo_2 _37652_ (.A1(_15990_),
    .A2(_15991_),
    .B1_N(_15992_),
    .X(_15993_));
 sky130_fd_sc_hd__nand3b_2 _37653_ (.A_N(_15992_),
    .B(_15990_),
    .C(_15991_),
    .Y(_15994_));
 sky130_fd_sc_hd__buf_1 _37654_ (.A(_15718_),
    .X(_15995_));
 sky130_fd_sc_hd__a21boi_2 _37655_ (.A1(_15854_),
    .A2(_15995_),
    .B1_N(_15855_),
    .Y(_15996_));
 sky130_fd_sc_hd__a21bo_2 _37656_ (.A1(_15993_),
    .A2(_15994_),
    .B1_N(_15996_),
    .X(_15997_));
 sky130_fd_sc_hd__nand3b_2 _37657_ (.A_N(_15996_),
    .B(_15993_),
    .C(_15994_),
    .Y(_15998_));
 sky130_fd_sc_hd__nand2_2 _37658_ (.A(_15997_),
    .B(_15998_),
    .Y(_15999_));
 sky130_fd_sc_hd__buf_1 _37659_ (.A(_15999_),
    .X(_16000_));
 sky130_fd_sc_hd__a21boi_2 _37660_ (.A1(_15977_),
    .A2(_15979_),
    .B1_N(_16000_),
    .Y(_16001_));
 sky130_fd_sc_hd__a21oi_2 _37661_ (.A1(_15978_),
    .A2(_15974_),
    .B1(_15976_),
    .Y(_16002_));
 sky130_vsdinv _37662_ (.A(_15979_),
    .Y(_16003_));
 sky130_fd_sc_hd__nor3_2 _37663_ (.A(_16000_),
    .B(_16002_),
    .C(_16003_),
    .Y(_16004_));
 sky130_fd_sc_hd__o21ai_2 _37664_ (.A1(_15863_),
    .A2(_15865_),
    .B1(_15846_),
    .Y(_16005_));
 sky130_fd_sc_hd__o21bai_2 _37665_ (.A1(_16001_),
    .A2(_16004_),
    .B1_N(_16005_),
    .Y(_16006_));
 sky130_fd_sc_hd__o21ai_2 _37666_ (.A1(_16002_),
    .A2(_16003_),
    .B1(_16000_),
    .Y(_16007_));
 sky130_fd_sc_hd__nand3b_2 _37667_ (.A_N(_15999_),
    .B(_15977_),
    .C(_15979_),
    .Y(_16008_));
 sky130_fd_sc_hd__nand3_2 _37668_ (.A(_16007_),
    .B(_16005_),
    .C(_16008_),
    .Y(_16009_));
 sky130_fd_sc_hd__a21oi_2 _37669_ (.A1(_14849_),
    .A2(_15873_),
    .B1(_15880_),
    .Y(_16010_));
 sky130_vsdinv _37670_ (.A(_16010_),
    .Y(_16011_));
 sky130_fd_sc_hd__nand3b_2 _37671_ (.A_N(_15847_),
    .B(_15859_),
    .C(_15860_),
    .Y(_16012_));
 sky130_fd_sc_hd__a21o_2 _37672_ (.A1(_16012_),
    .A2(_15860_),
    .B1(_15876_),
    .X(_16013_));
 sky130_fd_sc_hd__nand3_2 _37673_ (.A(_16012_),
    .B(_15860_),
    .C(_15878_),
    .Y(_16014_));
 sky130_fd_sc_hd__nand2_2 _37674_ (.A(_16013_),
    .B(_16014_),
    .Y(_16015_));
 sky130_fd_sc_hd__xor2_2 _37675_ (.A(_16011_),
    .B(_16015_),
    .X(_16016_));
 sky130_fd_sc_hd__buf_1 _37676_ (.A(_16016_),
    .X(_16017_));
 sky130_fd_sc_hd__a21boi_2 _37677_ (.A1(_16006_),
    .A2(_16009_),
    .B1_N(_16017_),
    .Y(_16018_));
 sky130_fd_sc_hd__a21oi_2 _37678_ (.A1(_16007_),
    .A2(_16008_),
    .B1(_16005_),
    .Y(_16019_));
 sky130_vsdinv _37679_ (.A(_16009_),
    .Y(_16020_));
 sky130_fd_sc_hd__nor3_2 _37680_ (.A(_16017_),
    .B(_16019_),
    .C(_16020_),
    .Y(_16021_));
 sky130_fd_sc_hd__o21ai_2 _37681_ (.A1(_15884_),
    .A2(_15891_),
    .B1(_15872_),
    .Y(_16022_));
 sky130_fd_sc_hd__o21bai_2 _37682_ (.A1(_16018_),
    .A2(_16021_),
    .B1_N(_16022_),
    .Y(_16023_));
 sky130_fd_sc_hd__o21ai_2 _37683_ (.A1(_16019_),
    .A2(_16020_),
    .B1(_16017_),
    .Y(_16024_));
 sky130_fd_sc_hd__nand3b_2 _37684_ (.A_N(_16016_),
    .B(_16006_),
    .C(_16009_),
    .Y(_16025_));
 sky130_fd_sc_hd__nand3_2 _37685_ (.A(_16024_),
    .B(_16022_),
    .C(_16025_),
    .Y(_16026_));
 sky130_fd_sc_hd__buf_1 _37686_ (.A(_15139_),
    .X(_16027_));
 sky130_fd_sc_hd__a21oi_2 _37687_ (.A1(_15883_),
    .A2(_15877_),
    .B1(_16027_),
    .Y(_16028_));
 sky130_fd_sc_hd__o211a_2 _37688_ (.A1(_15135_),
    .A2(_15137_),
    .B1(_15877_),
    .C1(_15883_),
    .X(_16029_));
 sky130_fd_sc_hd__nor3_2 _37689_ (.A(_15618_),
    .B(_16028_),
    .C(_16029_),
    .Y(_16030_));
 sky130_fd_sc_hd__o21a_2 _37690_ (.A1(_16028_),
    .A2(_16029_),
    .B1(_15305_),
    .X(_16031_));
 sky130_fd_sc_hd__nor2_2 _37691_ (.A(_16030_),
    .B(_16031_),
    .Y(_16032_));
 sky130_fd_sc_hd__a21oi_2 _37692_ (.A1(_16023_),
    .A2(_16026_),
    .B1(_16032_),
    .Y(_16033_));
 sky130_fd_sc_hd__nand3_2 _37693_ (.A(_16023_),
    .B(_16026_),
    .C(_16032_),
    .Y(_16034_));
 sky130_vsdinv _37694_ (.A(_16034_),
    .Y(_16035_));
 sky130_fd_sc_hd__o21ai_2 _37695_ (.A1(_15900_),
    .A2(_15902_),
    .B1(_15894_),
    .Y(_16036_));
 sky130_fd_sc_hd__o21bai_2 _37696_ (.A1(_16033_),
    .A2(_16035_),
    .B1_N(_16036_),
    .Y(_16037_));
 sky130_fd_sc_hd__o2bb2ai_2 _37697_ (.A1_N(_16026_),
    .A2_N(_16023_),
    .B1(_16030_),
    .B2(_16031_),
    .Y(_16038_));
 sky130_fd_sc_hd__nand3_2 _37698_ (.A(_16038_),
    .B(_16036_),
    .C(_16034_),
    .Y(_16039_));
 sky130_fd_sc_hd__buf_1 _37699_ (.A(_15160_),
    .X(_16040_));
 sky130_fd_sc_hd__nand2_2 _37700_ (.A(_15898_),
    .B(_15895_),
    .Y(_16041_));
 sky130_fd_sc_hd__xor2_2 _37701_ (.A(_16040_),
    .B(_16041_),
    .X(_16042_));
 sky130_fd_sc_hd__a21oi_2 _37702_ (.A1(_16037_),
    .A2(_16039_),
    .B1(_16042_),
    .Y(_16043_));
 sky130_fd_sc_hd__nand3_2 _37703_ (.A(_16037_),
    .B(_16039_),
    .C(_16042_),
    .Y(_16044_));
 sky130_vsdinv _37704_ (.A(_16044_),
    .Y(_16045_));
 sky130_vsdinv _37705_ (.A(_15911_),
    .Y(_16046_));
 sky130_fd_sc_hd__a21oi_2 _37706_ (.A1(_15907_),
    .A2(_15908_),
    .B1(_15905_),
    .Y(_16047_));
 sky130_fd_sc_hd__o21ai_2 _37707_ (.A1(_16046_),
    .A2(_16047_),
    .B1(_15909_),
    .Y(_16048_));
 sky130_fd_sc_hd__o21bai_2 _37708_ (.A1(_16043_),
    .A2(_16045_),
    .B1_N(_16048_),
    .Y(_16049_));
 sky130_fd_sc_hd__a21o_2 _37709_ (.A1(_16037_),
    .A2(_16039_),
    .B1(_16042_),
    .X(_16050_));
 sky130_fd_sc_hd__nand3_2 _37710_ (.A(_16050_),
    .B(_16048_),
    .C(_16044_),
    .Y(_16051_));
 sky130_fd_sc_hd__a21oi_2 _37711_ (.A1(_15773_),
    .A2(_15770_),
    .B1(_14976_),
    .Y(_16052_));
 sky130_fd_sc_hd__a21oi_2 _37712_ (.A1(_16049_),
    .A2(_16051_),
    .B1(_16052_),
    .Y(_16053_));
 sky130_fd_sc_hd__nand3_2 _37713_ (.A(_16049_),
    .B(_16052_),
    .C(_16051_),
    .Y(_16054_));
 sky130_vsdinv _37714_ (.A(_16054_),
    .Y(_16055_));
 sky130_fd_sc_hd__a21boi_2 _37715_ (.A1(_15921_),
    .A2(_15924_),
    .B1_N(_15918_),
    .Y(_16056_));
 sky130_fd_sc_hd__o21ai_2 _37716_ (.A1(_16053_),
    .A2(_16055_),
    .B1(_16056_),
    .Y(_16057_));
 sky130_fd_sc_hd__nand2_2 _37717_ (.A(_15925_),
    .B(_15918_),
    .Y(_16058_));
 sky130_fd_sc_hd__o2bb2ai_2 _37718_ (.A1_N(_16051_),
    .A2_N(_16049_),
    .B1(_15182_),
    .B2(_15910_),
    .Y(_16059_));
 sky130_fd_sc_hd__nand3_2 _37719_ (.A(_16058_),
    .B(_16054_),
    .C(_16059_),
    .Y(_16060_));
 sky130_fd_sc_hd__nand2_2 _37720_ (.A(_16057_),
    .B(_16060_),
    .Y(_16061_));
 sky130_fd_sc_hd__a21oi_2 _37721_ (.A1(_15935_),
    .A2(_15930_),
    .B1(_15929_),
    .Y(_16062_));
 sky130_fd_sc_hd__xor2_2 _37722_ (.A(_16061_),
    .B(_16062_),
    .X(_02674_));
 sky130_fd_sc_hd__buf_1 _37723_ (.A(_14701_),
    .X(_16063_));
 sky130_fd_sc_hd__buf_1 _37724_ (.A(_15558_),
    .X(_16064_));
 sky130_fd_sc_hd__and2_2 _37725_ (.A(_16063_),
    .B(_16064_),
    .X(_16065_));
 sky130_fd_sc_hd__buf_1 _37726_ (.A(_18713_),
    .X(_16066_));
 sky130_fd_sc_hd__buf_1 _37727_ (.A(_13580_),
    .X(_16067_));
 sky130_fd_sc_hd__buf_1 _37728_ (.A(_18719_),
    .X(_16068_));
 sky130_fd_sc_hd__a22oi_2 _37729_ (.A1(_16066_),
    .A2(_16067_),
    .B1(_16068_),
    .B2(_15827_),
    .Y(_16069_));
 sky130_fd_sc_hd__buf_1 _37730_ (.A(_13113_),
    .X(_16070_));
 sky130_fd_sc_hd__and4_2 _37731_ (.A(_18713_),
    .B(_18719_),
    .C(_16070_),
    .D(_16067_),
    .X(_16071_));
 sky130_fd_sc_hd__nor2_2 _37732_ (.A(_16069_),
    .B(_16071_),
    .Y(_16072_));
 sky130_fd_sc_hd__xor2_2 _37733_ (.A(_16065_),
    .B(_16072_),
    .X(_16073_));
 sky130_fd_sc_hd__nor3_2 _37734_ (.A(_12329_),
    .B(_16971_),
    .C(_15937_),
    .Y(_16074_));
 sky130_fd_sc_hd__a21o_2 _37735_ (.A1(_15939_),
    .A2(_15936_),
    .B1(_16074_),
    .X(_16075_));
 sky130_fd_sc_hd__and2_2 _37736_ (.A(_18706_),
    .B(_14666_),
    .X(_16076_));
 sky130_fd_sc_hd__nand2_2 _37737_ (.A(_18696_),
    .B(_12859_),
    .Y(_16077_));
 sky130_fd_sc_hd__nand2_2 _37738_ (.A(_19175_),
    .B(_11289_),
    .Y(_16078_));
 sky130_fd_sc_hd__xor2_2 _37739_ (.A(_16077_),
    .B(_16078_),
    .X(_16079_));
 sky130_fd_sc_hd__xor2_2 _37740_ (.A(_16076_),
    .B(_16079_),
    .X(_16080_));
 sky130_fd_sc_hd__xor2_2 _37741_ (.A(_16075_),
    .B(_16080_),
    .X(_16081_));
 sky130_fd_sc_hd__xor2_2 _37742_ (.A(_16073_),
    .B(_16081_),
    .X(_16082_));
 sky130_fd_sc_hd__nand3b_2 _37743_ (.A_N(_16082_),
    .B(_15946_),
    .C(_15953_),
    .Y(_16083_));
 sky130_fd_sc_hd__nor2_2 _37744_ (.A(_15942_),
    .B(_15940_),
    .Y(_16084_));
 sky130_fd_sc_hd__o21ai_2 _37745_ (.A1(_16084_),
    .A2(_15954_),
    .B1(_16082_),
    .Y(_16085_));
 sky130_fd_sc_hd__o21a_2 _37746_ (.A1(_15962_),
    .A2(_15963_),
    .B1(_15966_),
    .X(_16086_));
 sky130_fd_sc_hd__a21o_2 _37747_ (.A1(_15950_),
    .A2(_15947_),
    .B1(_15949_),
    .X(_16087_));
 sky130_fd_sc_hd__nand2_2 _37748_ (.A(_18729_),
    .B(_11199_),
    .Y(_16088_));
 sky130_fd_sc_hd__nand2_2 _37749_ (.A(_18736_),
    .B(_10900_),
    .Y(_16089_));
 sky130_fd_sc_hd__xor2_2 _37750_ (.A(_16088_),
    .B(_16089_),
    .X(_16090_));
 sky130_fd_sc_hd__a21o_2 _37751_ (.A1(_15981_),
    .A2(_08460_),
    .B1(_16090_),
    .X(_16091_));
 sky130_fd_sc_hd__and2_2 _37752_ (.A(_14830_),
    .B(_13508_),
    .X(_16092_));
 sky130_fd_sc_hd__nand2_2 _37753_ (.A(_16090_),
    .B(_16092_),
    .Y(_16093_));
 sky130_fd_sc_hd__nand2_2 _37754_ (.A(_16091_),
    .B(_16093_),
    .Y(_16094_));
 sky130_fd_sc_hd__xor2_2 _37755_ (.A(_16087_),
    .B(_16094_),
    .X(_16095_));
 sky130_fd_sc_hd__xor2_2 _37756_ (.A(_16086_),
    .B(_16095_),
    .X(_16096_));
 sky130_fd_sc_hd__a21o_2 _37757_ (.A1(_16083_),
    .A2(_16085_),
    .B1(_16096_),
    .X(_16097_));
 sky130_fd_sc_hd__nand3_2 _37758_ (.A(_16083_),
    .B(_16085_),
    .C(_16096_),
    .Y(_16098_));
 sky130_fd_sc_hd__nand2_2 _37759_ (.A(_15974_),
    .B(_15959_),
    .Y(_16099_));
 sky130_fd_sc_hd__a21o_2 _37760_ (.A1(_16097_),
    .A2(_16098_),
    .B1(_16099_),
    .X(_16100_));
 sky130_fd_sc_hd__nand3_2 _37761_ (.A(_16097_),
    .B(_16098_),
    .C(_16099_),
    .Y(_16101_));
 sky130_fd_sc_hd__and4_2 _37762_ (.A(_15980_),
    .B(_18750_),
    .C(_18755_),
    .D(_08086_),
    .X(_16102_));
 sky130_fd_sc_hd__a21oi_2 _37763_ (.A1(_15989_),
    .A2(_15995_),
    .B1(_16102_),
    .Y(_16103_));
 sky130_fd_sc_hd__o31ai_2 _37764_ (.A1(_18750_),
    .A2(_18756_),
    .A3(_07847_),
    .B1(_14831_),
    .Y(_16104_));
 sky130_fd_sc_hd__nor2_2 _37765_ (.A(_16102_),
    .B(_16104_),
    .Y(_16105_));
 sky130_fd_sc_hd__xor2_2 _37766_ (.A(_16105_),
    .B(_15720_),
    .X(_16106_));
 sky130_fd_sc_hd__buf_1 _37767_ (.A(_16106_),
    .X(_16107_));
 sky130_fd_sc_hd__o21ai_2 _37768_ (.A1(_15960_),
    .A2(_15968_),
    .B1(_15969_),
    .Y(_16108_));
 sky130_fd_sc_hd__xnor2_2 _37769_ (.A(_16107_),
    .B(_16108_),
    .Y(_16109_));
 sky130_fd_sc_hd__xor2_2 _37770_ (.A(_16103_),
    .B(_16109_),
    .X(_16110_));
 sky130_fd_sc_hd__a21oi_2 _37771_ (.A1(_16100_),
    .A2(_16101_),
    .B1(_16110_),
    .Y(_16111_));
 sky130_fd_sc_hd__nand3_2 _37772_ (.A(_16100_),
    .B(_16101_),
    .C(_16110_),
    .Y(_16112_));
 sky130_vsdinv _37773_ (.A(_16112_),
    .Y(_16113_));
 sky130_fd_sc_hd__o21ai_2 _37774_ (.A1(_16000_),
    .A2(_16002_),
    .B1(_15979_),
    .Y(_16114_));
 sky130_fd_sc_hd__o21bai_2 _37775_ (.A1(_16111_),
    .A2(_16113_),
    .B1_N(_16114_),
    .Y(_16115_));
 sky130_fd_sc_hd__a21o_2 _37776_ (.A1(_16100_),
    .A2(_16101_),
    .B1(_16110_),
    .X(_16116_));
 sky130_fd_sc_hd__nand3_2 _37777_ (.A(_16116_),
    .B(_16112_),
    .C(_16114_),
    .Y(_16117_));
 sky130_fd_sc_hd__buf_1 _37778_ (.A(_16011_),
    .X(_16118_));
 sky130_fd_sc_hd__buf_1 _37779_ (.A(_16118_),
    .X(_16119_));
 sky130_fd_sc_hd__buf_1 _37780_ (.A(_15878_),
    .X(_16120_));
 sky130_fd_sc_hd__a21o_2 _37781_ (.A1(_15998_),
    .A2(_15994_),
    .B1(_16120_),
    .X(_16121_));
 sky130_fd_sc_hd__buf_1 _37782_ (.A(_15878_),
    .X(_16122_));
 sky130_fd_sc_hd__nand3_2 _37783_ (.A(_15998_),
    .B(_16122_),
    .C(_15994_),
    .Y(_16123_));
 sky130_fd_sc_hd__nand2_2 _37784_ (.A(_16121_),
    .B(_16123_),
    .Y(_16124_));
 sky130_fd_sc_hd__xor2_2 _37785_ (.A(_16119_),
    .B(_16124_),
    .X(_16125_));
 sky130_fd_sc_hd__a21boi_2 _37786_ (.A1(_16115_),
    .A2(_16117_),
    .B1_N(_16125_),
    .Y(_16126_));
 sky130_fd_sc_hd__nand3b_2 _37787_ (.A_N(_16125_),
    .B(_16115_),
    .C(_16117_),
    .Y(_16127_));
 sky130_vsdinv _37788_ (.A(_16127_),
    .Y(_16128_));
 sky130_fd_sc_hd__o21ai_2 _37789_ (.A1(_16017_),
    .A2(_16019_),
    .B1(_16009_),
    .Y(_16129_));
 sky130_fd_sc_hd__o21bai_2 _37790_ (.A1(_16126_),
    .A2(_16128_),
    .B1_N(_16129_),
    .Y(_16130_));
 sky130_fd_sc_hd__a21oi_2 _37791_ (.A1(_16116_),
    .A2(_16112_),
    .B1(_16114_),
    .Y(_16131_));
 sky130_vsdinv _37792_ (.A(_16117_),
    .Y(_16132_));
 sky130_fd_sc_hd__o21ai_2 _37793_ (.A1(_16131_),
    .A2(_16132_),
    .B1(_16125_),
    .Y(_16133_));
 sky130_fd_sc_hd__nand3_2 _37794_ (.A(_16133_),
    .B(_16127_),
    .C(_16129_),
    .Y(_16134_));
 sky130_fd_sc_hd__buf_1 _37795_ (.A(_16010_),
    .X(_16135_));
 sky130_fd_sc_hd__o21ai_2 _37796_ (.A1(_16135_),
    .A2(_16015_),
    .B1(_16013_),
    .Y(_16136_));
 sky130_fd_sc_hd__xor2_2 _37797_ (.A(_15138_),
    .B(_16136_),
    .X(_16137_));
 sky130_fd_sc_hd__xor2_2 _37798_ (.A(_15633_),
    .B(_16137_),
    .X(_16138_));
 sky130_fd_sc_hd__a21oi_2 _37799_ (.A1(_16130_),
    .A2(_16134_),
    .B1(_16138_),
    .Y(_16139_));
 sky130_fd_sc_hd__nand3_2 _37800_ (.A(_16130_),
    .B(_16138_),
    .C(_16134_),
    .Y(_16140_));
 sky130_vsdinv _37801_ (.A(_16140_),
    .Y(_16141_));
 sky130_fd_sc_hd__nand2_2 _37802_ (.A(_16034_),
    .B(_16026_),
    .Y(_16142_));
 sky130_fd_sc_hd__o21bai_2 _37803_ (.A1(_16139_),
    .A2(_16141_),
    .B1_N(_16142_),
    .Y(_16143_));
 sky130_fd_sc_hd__a21oi_2 _37804_ (.A1(_16133_),
    .A2(_16127_),
    .B1(_16129_),
    .Y(_16144_));
 sky130_vsdinv _37805_ (.A(_16134_),
    .Y(_16145_));
 sky130_fd_sc_hd__o21bai_2 _37806_ (.A1(_16144_),
    .A2(_16145_),
    .B1_N(_16138_),
    .Y(_16146_));
 sky130_fd_sc_hd__nand3_2 _37807_ (.A(_16146_),
    .B(_16140_),
    .C(_16142_),
    .Y(_16147_));
 sky130_fd_sc_hd__buf_1 _37808_ (.A(_15618_),
    .X(_16148_));
 sky130_fd_sc_hd__buf_1 _37809_ (.A(_16148_),
    .X(_16149_));
 sky130_fd_sc_hd__o21ba_2 _37810_ (.A1(_16149_),
    .A2(_16029_),
    .B1_N(_16028_),
    .X(_16150_));
 sky130_fd_sc_hd__xor2_2 _37811_ (.A(_14812_),
    .B(_16150_),
    .X(_16151_));
 sky130_fd_sc_hd__a21oi_2 _37812_ (.A1(_16143_),
    .A2(_16147_),
    .B1(_16151_),
    .Y(_16152_));
 sky130_fd_sc_hd__nand3_2 _37813_ (.A(_16143_),
    .B(_16147_),
    .C(_16151_),
    .Y(_16153_));
 sky130_vsdinv _37814_ (.A(_16153_),
    .Y(_16154_));
 sky130_fd_sc_hd__nand2_2 _37815_ (.A(_16044_),
    .B(_16039_),
    .Y(_16155_));
 sky130_fd_sc_hd__o21bai_2 _37816_ (.A1(_16152_),
    .A2(_16154_),
    .B1_N(_16155_),
    .Y(_16156_));
 sky130_fd_sc_hd__a21oi_2 _37817_ (.A1(_16146_),
    .A2(_16140_),
    .B1(_16142_),
    .Y(_16157_));
 sky130_vsdinv _37818_ (.A(_16147_),
    .Y(_16158_));
 sky130_fd_sc_hd__o21bai_2 _37819_ (.A1(_16157_),
    .A2(_16158_),
    .B1_N(_16151_),
    .Y(_16159_));
 sky130_fd_sc_hd__nand3_2 _37820_ (.A(_16159_),
    .B(_16153_),
    .C(_16155_),
    .Y(_16160_));
 sky130_fd_sc_hd__a21oi_2 _37821_ (.A1(_15898_),
    .A2(_15895_),
    .B1(_15794_),
    .Y(_16161_));
 sky130_fd_sc_hd__a21oi_2 _37822_ (.A1(_16156_),
    .A2(_16160_),
    .B1(_16161_),
    .Y(_16162_));
 sky130_fd_sc_hd__nand3_2 _37823_ (.A(_16156_),
    .B(_16161_),
    .C(_16160_),
    .Y(_16163_));
 sky130_vsdinv _37824_ (.A(_16163_),
    .Y(_16164_));
 sky130_fd_sc_hd__nand2_2 _37825_ (.A(_16054_),
    .B(_16051_),
    .Y(_16165_));
 sky130_fd_sc_hd__o21bai_2 _37826_ (.A1(_16162_),
    .A2(_16164_),
    .B1_N(_16165_),
    .Y(_16166_));
 sky130_fd_sc_hd__a21o_2 _37827_ (.A1(_16156_),
    .A2(_16160_),
    .B1(_16161_),
    .X(_16167_));
 sky130_fd_sc_hd__nand3_2 _37828_ (.A(_16167_),
    .B(_16163_),
    .C(_16165_),
    .Y(_16168_));
 sky130_fd_sc_hd__nand2_2 _37829_ (.A(_16166_),
    .B(_16168_),
    .Y(_16169_));
 sky130_fd_sc_hd__nor3_2 _37830_ (.A(_15929_),
    .B(_15927_),
    .C(_16061_),
    .Y(_16170_));
 sky130_fd_sc_hd__nand2_2 _37831_ (.A(_16170_),
    .B(_15932_),
    .Y(_16171_));
 sky130_fd_sc_hd__nor2_2 _37832_ (.A(_16171_),
    .B(_15656_),
    .Y(_16172_));
 sky130_fd_sc_hd__a21boi_2 _37833_ (.A1(_15929_),
    .A2(_16057_),
    .B1_N(_16060_),
    .Y(_16173_));
 sky130_fd_sc_hd__a21boi_2 _37834_ (.A1(_16170_),
    .A2(_15934_),
    .B1_N(_16173_),
    .Y(_16174_));
 sky130_fd_sc_hd__o21ai_2 _37835_ (.A1(_16171_),
    .A2(_15660_),
    .B1(_16174_),
    .Y(_16175_));
 sky130_fd_sc_hd__a21oi_2 _37836_ (.A1(_15003_),
    .A2(_16172_),
    .B1(_16175_),
    .Y(_16176_));
 sky130_fd_sc_hd__xor2_2 _37837_ (.A(_16169_),
    .B(_16176_),
    .X(_02675_));
 sky130_fd_sc_hd__and2_2 _37838_ (.A(_16080_),
    .B(_16075_),
    .X(_16177_));
 sky130_fd_sc_hd__a21o_2 _37839_ (.A1(_16081_),
    .A2(_16073_),
    .B1(_16177_),
    .X(_16178_));
 sky130_fd_sc_hd__buf_1 _37840_ (.A(_10914_),
    .X(_16179_));
 sky130_fd_sc_hd__and2_2 _37841_ (.A(_16063_),
    .B(_16179_),
    .X(_16180_));
 sky130_fd_sc_hd__a22oi_2 _37842_ (.A1(_16066_),
    .A2(_15827_),
    .B1(_16068_),
    .B2(_15689_),
    .Y(_16181_));
 sky130_fd_sc_hd__and4_2 _37843_ (.A(_18713_),
    .B(_16068_),
    .C(_15558_),
    .D(_16070_),
    .X(_16182_));
 sky130_fd_sc_hd__nor2_2 _37844_ (.A(_16181_),
    .B(_16182_),
    .Y(_16183_));
 sky130_fd_sc_hd__xor2_2 _37845_ (.A(_16180_),
    .B(_16183_),
    .X(_16184_));
 sky130_fd_sc_hd__nor3_2 _37846_ (.A(_12330_),
    .B(_16971_),
    .C(_16077_),
    .Y(_16185_));
 sky130_fd_sc_hd__a21o_2 _37847_ (.A1(_16079_),
    .A2(_16076_),
    .B1(_16185_),
    .X(_16186_));
 sky130_fd_sc_hd__and2_2 _37848_ (.A(_18705_),
    .B(_16067_),
    .X(_16187_));
 sky130_fd_sc_hd__nand2_2 _37849_ (.A(_18696_),
    .B(_12596_),
    .Y(_16188_));
 sky130_fd_sc_hd__nand2_2 _37850_ (.A(_19169_),
    .B(_11289_),
    .Y(_16189_));
 sky130_fd_sc_hd__xor2_2 _37851_ (.A(_16188_),
    .B(_16189_),
    .X(_16190_));
 sky130_fd_sc_hd__xor2_2 _37852_ (.A(_16187_),
    .B(_16190_),
    .X(_16191_));
 sky130_fd_sc_hd__xor2_2 _37853_ (.A(_16186_),
    .B(_16191_),
    .X(_16192_));
 sky130_fd_sc_hd__xor2_2 _37854_ (.A(_16184_),
    .B(_16192_),
    .X(_16193_));
 sky130_fd_sc_hd__nor2_2 _37855_ (.A(_16178_),
    .B(_16193_),
    .Y(_16194_));
 sky130_fd_sc_hd__nand2_2 _37856_ (.A(_16193_),
    .B(_16178_),
    .Y(_16195_));
 sky130_vsdinv _37857_ (.A(_16195_),
    .Y(_16196_));
 sky130_fd_sc_hd__o21a_2 _37858_ (.A1(_16088_),
    .A2(_16089_),
    .B1(_16093_),
    .X(_16197_));
 sky130_fd_sc_hd__a21o_2 _37859_ (.A1(_16072_),
    .A2(_16065_),
    .B1(_16071_),
    .X(_16198_));
 sky130_vsdinv _37860_ (.A(_16092_),
    .Y(_16199_));
 sky130_fd_sc_hd__nand2_2 _37861_ (.A(_18730_),
    .B(_19134_),
    .Y(_16200_));
 sky130_fd_sc_hd__nand2_2 _37862_ (.A(_15980_),
    .B(_14716_),
    .Y(_16201_));
 sky130_fd_sc_hd__xor2_2 _37863_ (.A(_16200_),
    .B(_16201_),
    .X(_16202_));
 sky130_fd_sc_hd__xor2_2 _37864_ (.A(_16199_),
    .B(_16202_),
    .X(_16203_));
 sky130_fd_sc_hd__xnor2_2 _37865_ (.A(_16198_),
    .B(_16203_),
    .Y(_16204_));
 sky130_fd_sc_hd__xnor2_2 _37866_ (.A(_16197_),
    .B(_16204_),
    .Y(_16205_));
 sky130_fd_sc_hd__o21bai_2 _37867_ (.A1(_16194_),
    .A2(_16196_),
    .B1_N(_16205_),
    .Y(_16206_));
 sky130_fd_sc_hd__nand3b_2 _37868_ (.A_N(_16194_),
    .B(_16195_),
    .C(_16205_),
    .Y(_16207_));
 sky130_fd_sc_hd__nand2_2 _37869_ (.A(_16098_),
    .B(_16085_),
    .Y(_16208_));
 sky130_fd_sc_hd__a21o_2 _37870_ (.A1(_16206_),
    .A2(_16207_),
    .B1(_16208_),
    .X(_16209_));
 sky130_fd_sc_hd__nand3_2 _37871_ (.A(_16208_),
    .B(_16206_),
    .C(_16207_),
    .Y(_16210_));
 sky130_fd_sc_hd__nand2_2 _37872_ (.A(_16209_),
    .B(_16210_),
    .Y(_16211_));
 sky130_fd_sc_hd__or2_2 _37873_ (.A(_16086_),
    .B(_16095_),
    .X(_16212_));
 sky130_fd_sc_hd__nand3_2 _37874_ (.A(_16087_),
    .B(_16091_),
    .C(_16093_),
    .Y(_16213_));
 sky130_vsdinv _37875_ (.A(_16106_),
    .Y(_16214_));
 sky130_fd_sc_hd__a21o_2 _37876_ (.A1(_16212_),
    .A2(_16213_),
    .B1(_16214_),
    .X(_16215_));
 sky130_fd_sc_hd__buf_1 _37877_ (.A(_16214_),
    .X(_16216_));
 sky130_fd_sc_hd__o211ai_2 _37878_ (.A1(_16086_),
    .A2(_16095_),
    .B1(_16213_),
    .C1(_16216_),
    .Y(_16217_));
 sky130_fd_sc_hd__a21oi_2 _37879_ (.A1(_15995_),
    .A2(_16105_),
    .B1(_16102_),
    .Y(_16218_));
 sky130_vsdinv _37880_ (.A(_16218_),
    .Y(_16219_));
 sky130_fd_sc_hd__a21o_2 _37881_ (.A1(_16215_),
    .A2(_16217_),
    .B1(_16219_),
    .X(_16220_));
 sky130_fd_sc_hd__nand3_2 _37882_ (.A(_16215_),
    .B(_16219_),
    .C(_16217_),
    .Y(_16221_));
 sky130_fd_sc_hd__and2_2 _37883_ (.A(_16220_),
    .B(_16221_),
    .X(_16222_));
 sky130_vsdinv _37884_ (.A(_16222_),
    .Y(_16223_));
 sky130_fd_sc_hd__nand2_2 _37885_ (.A(_16211_),
    .B(_16223_),
    .Y(_16224_));
 sky130_fd_sc_hd__nand3_2 _37886_ (.A(_16209_),
    .B(_16222_),
    .C(_16210_),
    .Y(_16225_));
 sky130_vsdinv _37887_ (.A(_16110_),
    .Y(_16226_));
 sky130_fd_sc_hd__a21oi_2 _37888_ (.A1(_16097_),
    .A2(_16098_),
    .B1(_16099_),
    .Y(_16227_));
 sky130_fd_sc_hd__o21ai_2 _37889_ (.A1(_16226_),
    .A2(_16227_),
    .B1(_16101_),
    .Y(_16228_));
 sky130_fd_sc_hd__nand3_2 _37890_ (.A(_16224_),
    .B(_16225_),
    .C(_16228_),
    .Y(_16229_));
 sky130_fd_sc_hd__a21o_2 _37891_ (.A1(_16224_),
    .A2(_16225_),
    .B1(_16228_),
    .X(_16230_));
 sky130_fd_sc_hd__and2_2 _37892_ (.A(_16108_),
    .B(_16106_),
    .X(_16231_));
 sky130_fd_sc_hd__o21bai_2 _37893_ (.A1(_16103_),
    .A2(_16109_),
    .B1_N(_16231_),
    .Y(_16232_));
 sky130_fd_sc_hd__or2b_2 _37894_ (.A(_16232_),
    .B_N(_16120_),
    .X(_16233_));
 sky130_fd_sc_hd__nand2_2 _37895_ (.A(_16232_),
    .B(_15875_),
    .Y(_16234_));
 sky130_fd_sc_hd__and3_2 _37896_ (.A(_16233_),
    .B(_16118_),
    .C(_16234_),
    .X(_16235_));
 sky130_fd_sc_hd__buf_1 _37897_ (.A(_16118_),
    .X(_16236_));
 sky130_fd_sc_hd__a21oi_2 _37898_ (.A1(_16233_),
    .A2(_16234_),
    .B1(_16236_),
    .Y(_16237_));
 sky130_fd_sc_hd__o2bb2ai_2 _37899_ (.A1_N(_16229_),
    .A2_N(_16230_),
    .B1(_16235_),
    .B2(_16237_),
    .Y(_16238_));
 sky130_fd_sc_hd__o21ai_2 _37900_ (.A1(_16125_),
    .A2(_16131_),
    .B1(_16117_),
    .Y(_16239_));
 sky130_fd_sc_hd__nor2_2 _37901_ (.A(_16237_),
    .B(_16235_),
    .Y(_16240_));
 sky130_fd_sc_hd__nand3_2 _37902_ (.A(_16230_),
    .B(_16229_),
    .C(_16240_),
    .Y(_16241_));
 sky130_fd_sc_hd__nand3_2 _37903_ (.A(_16238_),
    .B(_16239_),
    .C(_16241_),
    .Y(_16242_));
 sky130_fd_sc_hd__a21oi_2 _37904_ (.A1(_16230_),
    .A2(_16229_),
    .B1(_16240_),
    .Y(_16243_));
 sky130_vsdinv _37905_ (.A(_16241_),
    .Y(_16244_));
 sky130_fd_sc_hd__o21bai_2 _37906_ (.A1(_16243_),
    .A2(_16244_),
    .B1_N(_16239_),
    .Y(_16245_));
 sky130_fd_sc_hd__nand3_2 _37907_ (.A(_16121_),
    .B(_16236_),
    .C(_16123_),
    .Y(_16246_));
 sky130_fd_sc_hd__buf_1 _37908_ (.A(_16027_),
    .X(_16247_));
 sky130_fd_sc_hd__a21oi_2 _37909_ (.A1(_16246_),
    .A2(_16121_),
    .B1(_16247_),
    .Y(_16248_));
 sky130_fd_sc_hd__o211a_2 _37910_ (.A1(_15135_),
    .A2(_15137_),
    .B1(_16121_),
    .C1(_16246_),
    .X(_16249_));
 sky130_fd_sc_hd__nor3_2 _37911_ (.A(_16148_),
    .B(_16248_),
    .C(_16249_),
    .Y(_16250_));
 sky130_fd_sc_hd__o21a_2 _37912_ (.A1(_16248_),
    .A2(_16249_),
    .B1(_15618_),
    .X(_16251_));
 sky130_fd_sc_hd__o2bb2ai_2 _37913_ (.A1_N(_16242_),
    .A2_N(_16245_),
    .B1(_16250_),
    .B2(_16251_),
    .Y(_16252_));
 sky130_fd_sc_hd__nor2_2 _37914_ (.A(_16250_),
    .B(_16251_),
    .Y(_16253_));
 sky130_fd_sc_hd__nand3_2 _37915_ (.A(_16245_),
    .B(_16242_),
    .C(_16253_),
    .Y(_16254_));
 sky130_vsdinv _37916_ (.A(_16138_),
    .Y(_16255_));
 sky130_fd_sc_hd__o21ai_2 _37917_ (.A1(_16255_),
    .A2(_16144_),
    .B1(_16134_),
    .Y(_16256_));
 sky130_fd_sc_hd__a21oi_2 _37918_ (.A1(_16252_),
    .A2(_16254_),
    .B1(_16256_),
    .Y(_16257_));
 sky130_fd_sc_hd__nand3_2 _37919_ (.A(_16252_),
    .B(_16256_),
    .C(_16254_),
    .Y(_16258_));
 sky130_vsdinv _37920_ (.A(_16258_),
    .Y(_16259_));
 sky130_fd_sc_hd__buf_1 _37921_ (.A(_15633_),
    .X(_16260_));
 sky130_fd_sc_hd__and2_2 _37922_ (.A(_16136_),
    .B(_15138_),
    .X(_16261_));
 sky130_fd_sc_hd__a21oi_2 _37923_ (.A1(_16137_),
    .A2(_16260_),
    .B1(_16261_),
    .Y(_16262_));
 sky130_fd_sc_hd__xor2_2 _37924_ (.A(_14975_),
    .B(_16262_),
    .X(_16263_));
 sky130_fd_sc_hd__o21bai_2 _37925_ (.A1(_16257_),
    .A2(_16259_),
    .B1_N(_16263_),
    .Y(_16264_));
 sky130_vsdinv _37926_ (.A(_16151_),
    .Y(_16265_));
 sky130_fd_sc_hd__o21ai_2 _37927_ (.A1(_16265_),
    .A2(_16157_),
    .B1(_16147_),
    .Y(_16266_));
 sky130_fd_sc_hd__a21oi_2 _37928_ (.A1(_16245_),
    .A2(_16242_),
    .B1(_16253_),
    .Y(_16267_));
 sky130_vsdinv _37929_ (.A(_16254_),
    .Y(_16268_));
 sky130_fd_sc_hd__o21bai_2 _37930_ (.A1(_16267_),
    .A2(_16268_),
    .B1_N(_16256_),
    .Y(_16269_));
 sky130_fd_sc_hd__nand3_2 _37931_ (.A(_16269_),
    .B(_16258_),
    .C(_16263_),
    .Y(_16270_));
 sky130_fd_sc_hd__nand3_2 _37932_ (.A(_16264_),
    .B(_16266_),
    .C(_16270_),
    .Y(_16271_));
 sky130_fd_sc_hd__a21oi_2 _37933_ (.A1(_16269_),
    .A2(_16258_),
    .B1(_16263_),
    .Y(_16272_));
 sky130_vsdinv _37934_ (.A(_16270_),
    .Y(_16273_));
 sky130_fd_sc_hd__o21bai_2 _37935_ (.A1(_16272_),
    .A2(_16273_),
    .B1_N(_16266_),
    .Y(_16274_));
 sky130_fd_sc_hd__o2bb2ai_2 _37936_ (.A1_N(_16271_),
    .A2_N(_16274_),
    .B1(_15922_),
    .B2(_16150_),
    .Y(_16275_));
 sky130_fd_sc_hd__nor2_2 _37937_ (.A(_15794_),
    .B(_16150_),
    .Y(_16276_));
 sky130_fd_sc_hd__nand3_2 _37938_ (.A(_16274_),
    .B(_16276_),
    .C(_16271_),
    .Y(_16277_));
 sky130_vsdinv _37939_ (.A(_16161_),
    .Y(_16278_));
 sky130_fd_sc_hd__a21oi_2 _37940_ (.A1(_16159_),
    .A2(_16153_),
    .B1(_16155_),
    .Y(_16279_));
 sky130_fd_sc_hd__o21ai_2 _37941_ (.A1(_16278_),
    .A2(_16279_),
    .B1(_16160_),
    .Y(_16280_));
 sky130_fd_sc_hd__a21o_2 _37942_ (.A1(_16275_),
    .A2(_16277_),
    .B1(_16280_),
    .X(_16281_));
 sky130_fd_sc_hd__nand3_2 _37943_ (.A(_16275_),
    .B(_16280_),
    .C(_16277_),
    .Y(_16282_));
 sky130_fd_sc_hd__nand2_2 _37944_ (.A(_16281_),
    .B(_16282_),
    .Y(_16283_));
 sky130_fd_sc_hd__o21ai_2 _37945_ (.A1(_16169_),
    .A2(_16176_),
    .B1(_16168_),
    .Y(_16284_));
 sky130_fd_sc_hd__xnor2_2 _37946_ (.A(_16283_),
    .B(_16284_),
    .Y(_02676_));
 sky130_fd_sc_hd__and2_2 _37947_ (.A(_16191_),
    .B(_16186_),
    .X(_16285_));
 sky130_fd_sc_hd__a21o_2 _37948_ (.A1(_16192_),
    .A2(_16184_),
    .B1(_16285_),
    .X(_16286_));
 sky130_fd_sc_hd__and2_2 _37949_ (.A(_16063_),
    .B(_19136_),
    .X(_16287_));
 sky130_fd_sc_hd__a22oi_2 _37950_ (.A1(_18714_),
    .A2(_16064_),
    .B1(_18720_),
    .B2(_16179_),
    .Y(_16288_));
 sky130_fd_sc_hd__and4_2 _37951_ (.A(_16066_),
    .B(_16068_),
    .C(_10915_),
    .D(_15689_),
    .X(_16289_));
 sky130_fd_sc_hd__nor2_2 _37952_ (.A(_16288_),
    .B(_16289_),
    .Y(_16290_));
 sky130_fd_sc_hd__xor2_2 _37953_ (.A(_16287_),
    .B(_16290_),
    .X(_16291_));
 sky130_fd_sc_hd__nor3_2 _37954_ (.A(_12859_),
    .B(_16971_),
    .C(_16188_),
    .Y(_16292_));
 sky130_fd_sc_hd__a21o_2 _37955_ (.A1(_16190_),
    .A2(_16187_),
    .B1(_16292_),
    .X(_16293_));
 sky130_fd_sc_hd__and2_2 _37956_ (.A(_18706_),
    .B(_16070_),
    .X(_16294_));
 sky130_fd_sc_hd__nand2_2 _37957_ (.A(_18697_),
    .B(_13369_),
    .Y(_16295_));
 sky130_fd_sc_hd__nand2_2 _37958_ (.A(_19164_),
    .B(_11290_),
    .Y(_16296_));
 sky130_fd_sc_hd__xor2_2 _37959_ (.A(_16295_),
    .B(_16296_),
    .X(_16297_));
 sky130_fd_sc_hd__xor2_2 _37960_ (.A(_16294_),
    .B(_16297_),
    .X(_16298_));
 sky130_fd_sc_hd__xor2_2 _37961_ (.A(_16293_),
    .B(_16298_),
    .X(_16299_));
 sky130_fd_sc_hd__xor2_2 _37962_ (.A(_16291_),
    .B(_16299_),
    .X(_16300_));
 sky130_fd_sc_hd__nor2_2 _37963_ (.A(_16286_),
    .B(_16300_),
    .Y(_16301_));
 sky130_fd_sc_hd__nand2_2 _37964_ (.A(_16300_),
    .B(_16286_),
    .Y(_16302_));
 sky130_vsdinv _37965_ (.A(_16302_),
    .Y(_16303_));
 sky130_fd_sc_hd__nor2_2 _37966_ (.A(_16200_),
    .B(_16201_),
    .Y(_16304_));
 sky130_fd_sc_hd__a21oi_2 _37967_ (.A1(_16202_),
    .A2(_16092_),
    .B1(_16304_),
    .Y(_16305_));
 sky130_fd_sc_hd__a21o_2 _37968_ (.A1(_16183_),
    .A2(_16180_),
    .B1(_16182_),
    .X(_16306_));
 sky130_fd_sc_hd__nand2_2 _37969_ (.A(_15980_),
    .B(_18730_),
    .Y(_16307_));
 sky130_fd_sc_hd__xnor2_2 _37970_ (.A(_16201_),
    .B(_16307_),
    .Y(_16308_));
 sky130_fd_sc_hd__xor2_2 _37971_ (.A(_16199_),
    .B(_16308_),
    .X(_16309_));
 sky130_fd_sc_hd__xnor2_2 _37972_ (.A(_16306_),
    .B(_16309_),
    .Y(_16310_));
 sky130_fd_sc_hd__xor2_2 _37973_ (.A(_16305_),
    .B(_16310_),
    .X(_16311_));
 sky130_fd_sc_hd__o21bai_2 _37974_ (.A1(_16301_),
    .A2(_16303_),
    .B1_N(_16311_),
    .Y(_16312_));
 sky130_fd_sc_hd__nand3b_2 _37975_ (.A_N(_16301_),
    .B(_16302_),
    .C(_16311_),
    .Y(_16313_));
 sky130_fd_sc_hd__nand2_2 _37976_ (.A(_16207_),
    .B(_16195_),
    .Y(_16314_));
 sky130_fd_sc_hd__a21o_2 _37977_ (.A1(_16312_),
    .A2(_16313_),
    .B1(_16314_),
    .X(_16315_));
 sky130_fd_sc_hd__nand3_2 _37978_ (.A(_16314_),
    .B(_16312_),
    .C(_16313_),
    .Y(_16316_));
 sky130_fd_sc_hd__or2b_2 _37979_ (.A(_16197_),
    .B_N(_16204_),
    .X(_16317_));
 sky130_fd_sc_hd__or2b_2 _37980_ (.A(_16203_),
    .B_N(_16198_),
    .X(_16318_));
 sky130_fd_sc_hd__a21o_2 _37981_ (.A1(_16317_),
    .A2(_16318_),
    .B1(_16216_),
    .X(_16319_));
 sky130_fd_sc_hd__nand3_2 _37982_ (.A(_16317_),
    .B(_16216_),
    .C(_16318_),
    .Y(_16320_));
 sky130_fd_sc_hd__nand2_2 _37983_ (.A(_16319_),
    .B(_16320_),
    .Y(_16321_));
 sky130_fd_sc_hd__xor2_2 _37984_ (.A(_16218_),
    .B(_16321_),
    .X(_16322_));
 sky130_fd_sc_hd__a21o_2 _37985_ (.A1(_16315_),
    .A2(_16316_),
    .B1(_16322_),
    .X(_16323_));
 sky130_fd_sc_hd__nand3_2 _37986_ (.A(_16315_),
    .B(_16316_),
    .C(_16322_),
    .Y(_16324_));
 sky130_fd_sc_hd__a21oi_2 _37987_ (.A1(_16206_),
    .A2(_16207_),
    .B1(_16208_),
    .Y(_16325_));
 sky130_fd_sc_hd__o21ai_2 _37988_ (.A1(_16325_),
    .A2(_16223_),
    .B1(_16210_),
    .Y(_16326_));
 sky130_fd_sc_hd__nand3_2 _37989_ (.A(_16323_),
    .B(_16324_),
    .C(_16326_),
    .Y(_16327_));
 sky130_fd_sc_hd__a21oi_2 _37990_ (.A1(_16315_),
    .A2(_16316_),
    .B1(_16322_),
    .Y(_16328_));
 sky130_vsdinv _37991_ (.A(_16324_),
    .Y(_16329_));
 sky130_fd_sc_hd__o21bai_2 _37992_ (.A1(_16328_),
    .A2(_16329_),
    .B1_N(_16326_),
    .Y(_16330_));
 sky130_fd_sc_hd__a21o_2 _37993_ (.A1(_16221_),
    .A2(_16215_),
    .B1(_16120_),
    .X(_16331_));
 sky130_fd_sc_hd__nand3_2 _37994_ (.A(_16221_),
    .B(_16120_),
    .C(_16215_),
    .Y(_16332_));
 sky130_fd_sc_hd__and3_2 _37995_ (.A(_16331_),
    .B(_16118_),
    .C(_16332_),
    .X(_16333_));
 sky130_fd_sc_hd__a21oi_2 _37996_ (.A1(_16331_),
    .A2(_16332_),
    .B1(_16236_),
    .Y(_16334_));
 sky130_fd_sc_hd__o2bb2ai_2 _37997_ (.A1_N(_16327_),
    .A2_N(_16330_),
    .B1(_16333_),
    .B2(_16334_),
    .Y(_16335_));
 sky130_fd_sc_hd__nor2_2 _37998_ (.A(_16334_),
    .B(_16333_),
    .Y(_16336_));
 sky130_fd_sc_hd__nand3_2 _37999_ (.A(_16330_),
    .B(_16327_),
    .C(_16336_),
    .Y(_16337_));
 sky130_vsdinv _38000_ (.A(_16240_),
    .Y(_16338_));
 sky130_fd_sc_hd__a21oi_2 _38001_ (.A1(_16224_),
    .A2(_16225_),
    .B1(_16228_),
    .Y(_16339_));
 sky130_fd_sc_hd__o21ai_2 _38002_ (.A1(_16338_),
    .A2(_16339_),
    .B1(_16229_),
    .Y(_16340_));
 sky130_fd_sc_hd__nand3_2 _38003_ (.A(_16335_),
    .B(_16337_),
    .C(_16340_),
    .Y(_16341_));
 sky130_fd_sc_hd__a21oi_2 _38004_ (.A1(_16330_),
    .A2(_16327_),
    .B1(_16336_),
    .Y(_16342_));
 sky130_vsdinv _38005_ (.A(_16337_),
    .Y(_16343_));
 sky130_fd_sc_hd__o21bai_2 _38006_ (.A1(_16342_),
    .A2(_16343_),
    .B1_N(_16340_),
    .Y(_16344_));
 sky130_fd_sc_hd__a21boi_2 _38007_ (.A1(_16233_),
    .A2(_16236_),
    .B1_N(_16234_),
    .Y(_16345_));
 sky130_fd_sc_hd__nor2_2 _38008_ (.A(_16027_),
    .B(_16345_),
    .Y(_16346_));
 sky130_fd_sc_hd__nand2_2 _38009_ (.A(_16345_),
    .B(_16027_),
    .Y(_16347_));
 sky130_fd_sc_hd__nor3b_2 _38010_ (.A(_16148_),
    .B(_16346_),
    .C_N(_16347_),
    .Y(_16348_));
 sky130_vsdinv _38011_ (.A(_16346_),
    .Y(_16349_));
 sky130_fd_sc_hd__a21oi_2 _38012_ (.A1(_16349_),
    .A2(_16347_),
    .B1(_15633_),
    .Y(_16350_));
 sky130_fd_sc_hd__o2bb2ai_2 _38013_ (.A1_N(_16341_),
    .A2_N(_16344_),
    .B1(_16348_),
    .B2(_16350_),
    .Y(_16351_));
 sky130_fd_sc_hd__nor2_2 _38014_ (.A(_16348_),
    .B(_16350_),
    .Y(_16352_));
 sky130_fd_sc_hd__nand3_2 _38015_ (.A(_16344_),
    .B(_16352_),
    .C(_16341_),
    .Y(_16353_));
 sky130_vsdinv _38016_ (.A(_16253_),
    .Y(_16354_));
 sky130_fd_sc_hd__a21oi_2 _38017_ (.A1(_16238_),
    .A2(_16241_),
    .B1(_16239_),
    .Y(_16355_));
 sky130_fd_sc_hd__o21ai_2 _38018_ (.A1(_16354_),
    .A2(_16355_),
    .B1(_16242_),
    .Y(_16356_));
 sky130_fd_sc_hd__a21oi_2 _38019_ (.A1(_16351_),
    .A2(_16353_),
    .B1(_16356_),
    .Y(_16357_));
 sky130_fd_sc_hd__nand3_2 _38020_ (.A(_16351_),
    .B(_16356_),
    .C(_16353_),
    .Y(_16358_));
 sky130_vsdinv _38021_ (.A(_16358_),
    .Y(_16359_));
 sky130_fd_sc_hd__o21ba_2 _38022_ (.A1(_16149_),
    .A2(_16249_),
    .B1_N(_16248_),
    .X(_16360_));
 sky130_fd_sc_hd__xor2_2 _38023_ (.A(_14975_),
    .B(_16360_),
    .X(_16361_));
 sky130_fd_sc_hd__o21bai_2 _38024_ (.A1(_16357_),
    .A2(_16359_),
    .B1_N(_16361_),
    .Y(_16362_));
 sky130_fd_sc_hd__a21o_2 _38025_ (.A1(_16351_),
    .A2(_16353_),
    .B1(_16356_),
    .X(_16363_));
 sky130_fd_sc_hd__nand3_2 _38026_ (.A(_16363_),
    .B(_16358_),
    .C(_16361_),
    .Y(_16364_));
 sky130_vsdinv _38027_ (.A(_16263_),
    .Y(_16365_));
 sky130_fd_sc_hd__o21ai_2 _38028_ (.A1(_16365_),
    .A2(_16257_),
    .B1(_16258_),
    .Y(_16366_));
 sky130_fd_sc_hd__a21oi_2 _38029_ (.A1(_16362_),
    .A2(_16364_),
    .B1(_16366_),
    .Y(_16367_));
 sky130_fd_sc_hd__nand3_2 _38030_ (.A(_16362_),
    .B(_16366_),
    .C(_16364_),
    .Y(_16368_));
 sky130_vsdinv _38031_ (.A(_16368_),
    .Y(_16369_));
 sky130_fd_sc_hd__nor2_2 _38032_ (.A(_15182_),
    .B(_16262_),
    .Y(_16370_));
 sky130_fd_sc_hd__o21bai_2 _38033_ (.A1(_16367_),
    .A2(_16369_),
    .B1_N(_16370_),
    .Y(_16371_));
 sky130_fd_sc_hd__a21o_2 _38034_ (.A1(_16362_),
    .A2(_16364_),
    .B1(_16366_),
    .X(_16372_));
 sky130_fd_sc_hd__nand3_2 _38035_ (.A(_16372_),
    .B(_16370_),
    .C(_16368_),
    .Y(_16373_));
 sky130_vsdinv _38036_ (.A(_16276_),
    .Y(_16374_));
 sky130_fd_sc_hd__a21oi_2 _38037_ (.A1(_16264_),
    .A2(_16270_),
    .B1(_16266_),
    .Y(_16375_));
 sky130_fd_sc_hd__o21ai_2 _38038_ (.A1(_16374_),
    .A2(_16375_),
    .B1(_16271_),
    .Y(_16376_));
 sky130_fd_sc_hd__a21o_2 _38039_ (.A1(_16371_),
    .A2(_16373_),
    .B1(_16376_),
    .X(_16377_));
 sky130_fd_sc_hd__nand3_2 _38040_ (.A(_16371_),
    .B(_16376_),
    .C(_16373_),
    .Y(_16378_));
 sky130_fd_sc_hd__nand2_2 _38041_ (.A(_16377_),
    .B(_16378_),
    .Y(_16379_));
 sky130_fd_sc_hd__a21oi_2 _38042_ (.A1(_16275_),
    .A2(_16277_),
    .B1(_16280_),
    .Y(_16380_));
 sky130_fd_sc_hd__a21oi_2 _38043_ (.A1(_16168_),
    .A2(_16282_),
    .B1(_16380_),
    .Y(_16381_));
 sky130_fd_sc_hd__nor3_2 _38044_ (.A(_16169_),
    .B(_16283_),
    .C(_16176_),
    .Y(_16382_));
 sky130_fd_sc_hd__nor2_2 _38045_ (.A(_16381_),
    .B(_16382_),
    .Y(_16383_));
 sky130_fd_sc_hd__xor2_2 _38046_ (.A(_16379_),
    .B(_16383_),
    .X(_02677_));
 sky130_fd_sc_hd__nand2_2 _38047_ (.A(_16313_),
    .B(_16302_),
    .Y(_16384_));
 sky130_fd_sc_hd__and2_2 _38048_ (.A(_16298_),
    .B(_16293_),
    .X(_16385_));
 sky130_fd_sc_hd__a21o_2 _38049_ (.A1(_16299_),
    .A2(_16291_),
    .B1(_16385_),
    .X(_16386_));
 sky130_fd_sc_hd__buf_1 _38050_ (.A(_14831_),
    .X(_16387_));
 sky130_fd_sc_hd__nand2_2 _38051_ (.A(_16387_),
    .B(_16063_),
    .Y(_16388_));
 sky130_fd_sc_hd__nand2_2 _38052_ (.A(_18714_),
    .B(_16179_),
    .Y(_16389_));
 sky130_fd_sc_hd__nand2_2 _38053_ (.A(_18720_),
    .B(_19136_),
    .Y(_16390_));
 sky130_fd_sc_hd__xnor2_2 _38054_ (.A(_16389_),
    .B(_16390_),
    .Y(_16391_));
 sky130_fd_sc_hd__xor2_2 _38055_ (.A(_16388_),
    .B(_16391_),
    .X(_16392_));
 sky130_fd_sc_hd__nor3_2 _38056_ (.A(_14666_),
    .B(_16972_),
    .C(_16295_),
    .Y(_16393_));
 sky130_fd_sc_hd__a21o_2 _38057_ (.A1(_16297_),
    .A2(_16294_),
    .B1(_16393_),
    .X(_16394_));
 sky130_fd_sc_hd__and2_2 _38058_ (.A(_18706_),
    .B(_16064_),
    .X(_16395_));
 sky130_fd_sc_hd__nand2_2 _38059_ (.A(_18697_),
    .B(_16070_),
    .Y(_16396_));
 sky130_fd_sc_hd__nand2_2 _38060_ (.A(_19159_),
    .B(_11290_),
    .Y(_16397_));
 sky130_fd_sc_hd__xor2_2 _38061_ (.A(_16396_),
    .B(_16397_),
    .X(_16398_));
 sky130_fd_sc_hd__xor2_2 _38062_ (.A(_16395_),
    .B(_16398_),
    .X(_16399_));
 sky130_fd_sc_hd__xor2_2 _38063_ (.A(_16394_),
    .B(_16399_),
    .X(_16400_));
 sky130_fd_sc_hd__xor2_2 _38064_ (.A(_16392_),
    .B(_16400_),
    .X(_16401_));
 sky130_fd_sc_hd__nor2_2 _38065_ (.A(_16386_),
    .B(_16401_),
    .Y(_16402_));
 sky130_fd_sc_hd__nand2_2 _38066_ (.A(_16401_),
    .B(_16386_),
    .Y(_16403_));
 sky130_vsdinv _38067_ (.A(_16403_),
    .Y(_16404_));
 sky130_fd_sc_hd__nand3_2 _38068_ (.A(_16387_),
    .B(_18730_),
    .C(_18737_),
    .Y(_16405_));
 sky130_fd_sc_hd__o21a_2 _38069_ (.A1(_16199_),
    .A2(_16308_),
    .B1(_16405_),
    .X(_16406_));
 sky130_fd_sc_hd__buf_1 _38070_ (.A(_16406_),
    .X(_16407_));
 sky130_fd_sc_hd__a21o_2 _38071_ (.A1(_16290_),
    .A2(_16287_),
    .B1(_16289_),
    .X(_16408_));
 sky130_fd_sc_hd__xnor2_2 _38072_ (.A(_16408_),
    .B(_16309_),
    .Y(_16409_));
 sky130_fd_sc_hd__xor2_2 _38073_ (.A(_16407_),
    .B(_16409_),
    .X(_16410_));
 sky130_fd_sc_hd__o21bai_2 _38074_ (.A1(_16402_),
    .A2(_16404_),
    .B1_N(_16410_),
    .Y(_16411_));
 sky130_fd_sc_hd__nand3b_2 _38075_ (.A_N(_16402_),
    .B(_16403_),
    .C(_16410_),
    .Y(_16412_));
 sky130_fd_sc_hd__nand3_2 _38076_ (.A(_16384_),
    .B(_16411_),
    .C(_16412_),
    .Y(_16413_));
 sky130_fd_sc_hd__a21o_2 _38077_ (.A1(_16411_),
    .A2(_16412_),
    .B1(_16384_),
    .X(_16414_));
 sky130_fd_sc_hd__or2_2 _38078_ (.A(_16305_),
    .B(_16310_),
    .X(_16415_));
 sky130_fd_sc_hd__buf_1 _38079_ (.A(_16309_),
    .X(_16416_));
 sky130_fd_sc_hd__nand2_2 _38080_ (.A(_16416_),
    .B(_16306_),
    .Y(_16417_));
 sky130_fd_sc_hd__buf_1 _38081_ (.A(_16214_),
    .X(_16418_));
 sky130_fd_sc_hd__a21o_2 _38082_ (.A1(_16415_),
    .A2(_16417_),
    .B1(_16418_),
    .X(_16419_));
 sky130_fd_sc_hd__o211ai_2 _38083_ (.A1(_16305_),
    .A2(_16310_),
    .B1(_16216_),
    .C1(_16417_),
    .Y(_16420_));
 sky130_fd_sc_hd__and3_2 _38084_ (.A(_16419_),
    .B(_16219_),
    .C(_16420_),
    .X(_16421_));
 sky130_fd_sc_hd__buf_1 _38085_ (.A(_16219_),
    .X(_16422_));
 sky130_fd_sc_hd__a21oi_2 _38086_ (.A1(_16419_),
    .A2(_16420_),
    .B1(_16422_),
    .Y(_16423_));
 sky130_fd_sc_hd__o2bb2ai_2 _38087_ (.A1_N(_16413_),
    .A2_N(_16414_),
    .B1(_16421_),
    .B2(_16423_),
    .Y(_16424_));
 sky130_fd_sc_hd__a21o_2 _38088_ (.A1(_16419_),
    .A2(_16420_),
    .B1(_16422_),
    .X(_16425_));
 sky130_fd_sc_hd__and2b_2 _38089_ (.A_N(_16421_),
    .B(_16425_),
    .X(_16426_));
 sky130_fd_sc_hd__nand3_2 _38090_ (.A(_16414_),
    .B(_16413_),
    .C(_16426_),
    .Y(_16427_));
 sky130_fd_sc_hd__nand2_2 _38091_ (.A(_16324_),
    .B(_16316_),
    .Y(_16428_));
 sky130_fd_sc_hd__a21o_2 _38092_ (.A1(_16424_),
    .A2(_16427_),
    .B1(_16428_),
    .X(_16429_));
 sky130_fd_sc_hd__nand3_2 _38093_ (.A(_16428_),
    .B(_16424_),
    .C(_16427_),
    .Y(_16430_));
 sky130_fd_sc_hd__nand3_2 _38094_ (.A(_16319_),
    .B(_16422_),
    .C(_16320_),
    .Y(_16431_));
 sky130_fd_sc_hd__a21o_2 _38095_ (.A1(_16431_),
    .A2(_16319_),
    .B1(_16122_),
    .X(_16432_));
 sky130_fd_sc_hd__nand3_2 _38096_ (.A(_16431_),
    .B(_16122_),
    .C(_16319_),
    .Y(_16433_));
 sky130_fd_sc_hd__nand2_2 _38097_ (.A(_16432_),
    .B(_16433_),
    .Y(_16434_));
 sky130_fd_sc_hd__xor2_2 _38098_ (.A(_16135_),
    .B(_16434_),
    .X(_16435_));
 sky130_fd_sc_hd__a21oi_2 _38099_ (.A1(_16429_),
    .A2(_16430_),
    .B1(_16435_),
    .Y(_16436_));
 sky130_fd_sc_hd__nand3_2 _38100_ (.A(_16429_),
    .B(_16430_),
    .C(_16435_),
    .Y(_16437_));
 sky130_vsdinv _38101_ (.A(_16437_),
    .Y(_16438_));
 sky130_fd_sc_hd__nand2_2 _38102_ (.A(_16337_),
    .B(_16327_),
    .Y(_16439_));
 sky130_fd_sc_hd__o21bai_2 _38103_ (.A1(_16436_),
    .A2(_16438_),
    .B1_N(_16439_),
    .Y(_16440_));
 sky130_fd_sc_hd__a21o_2 _38104_ (.A1(_16429_),
    .A2(_16430_),
    .B1(_16435_),
    .X(_16441_));
 sky130_fd_sc_hd__nand3_2 _38105_ (.A(_16441_),
    .B(_16439_),
    .C(_16437_),
    .Y(_16442_));
 sky130_fd_sc_hd__a21boi_2 _38106_ (.A1(_16119_),
    .A2(_16332_),
    .B1_N(_16331_),
    .Y(_16443_));
 sky130_fd_sc_hd__nor2_2 _38107_ (.A(_16247_),
    .B(_16443_),
    .Y(_16444_));
 sky130_fd_sc_hd__nand2_2 _38108_ (.A(_16443_),
    .B(_16247_),
    .Y(_16445_));
 sky130_fd_sc_hd__nor3b_2 _38109_ (.A(_16148_),
    .B(_16444_),
    .C_N(_16445_),
    .Y(_16446_));
 sky130_vsdinv _38110_ (.A(_16444_),
    .Y(_16447_));
 sky130_fd_sc_hd__a21oi_2 _38111_ (.A1(_16447_),
    .A2(_16445_),
    .B1(_16260_),
    .Y(_16448_));
 sky130_fd_sc_hd__nor2_2 _38112_ (.A(_16446_),
    .B(_16448_),
    .Y(_16449_));
 sky130_fd_sc_hd__a21oi_2 _38113_ (.A1(_16440_),
    .A2(_16442_),
    .B1(_16449_),
    .Y(_16450_));
 sky130_fd_sc_hd__nand3_2 _38114_ (.A(_16440_),
    .B(_16449_),
    .C(_16442_),
    .Y(_16451_));
 sky130_fd_sc_hd__nand2_2 _38115_ (.A(_16353_),
    .B(_16341_),
    .Y(_16452_));
 sky130_fd_sc_hd__nand3b_2 _38116_ (.A_N(_16450_),
    .B(_16451_),
    .C(_16452_),
    .Y(_16453_));
 sky130_vsdinv _38117_ (.A(_16451_),
    .Y(_16454_));
 sky130_fd_sc_hd__o21bai_2 _38118_ (.A1(_16450_),
    .A2(_16454_),
    .B1_N(_16452_),
    .Y(_16455_));
 sky130_fd_sc_hd__a21oi_2 _38119_ (.A1(_16347_),
    .A2(_16260_),
    .B1(_16346_),
    .Y(_16456_));
 sky130_fd_sc_hd__nor2_2 _38120_ (.A(_14812_),
    .B(_16456_),
    .Y(_16457_));
 sky130_fd_sc_hd__buf_1 _38121_ (.A(_16260_),
    .X(_16458_));
 sky130_fd_sc_hd__a211oi_2 _38122_ (.A1(_16347_),
    .A2(_16458_),
    .B1(_16040_),
    .C1(_16346_),
    .Y(_16459_));
 sky130_fd_sc_hd__o2bb2ai_2 _38123_ (.A1_N(_16453_),
    .A2_N(_16455_),
    .B1(_16457_),
    .B2(_16459_),
    .Y(_16460_));
 sky130_fd_sc_hd__nor2_2 _38124_ (.A(_16459_),
    .B(_16457_),
    .Y(_16461_));
 sky130_fd_sc_hd__nand3_2 _38125_ (.A(_16455_),
    .B(_16453_),
    .C(_16461_),
    .Y(_16462_));
 sky130_vsdinv _38126_ (.A(_16361_),
    .Y(_16463_));
 sky130_fd_sc_hd__o21ai_2 _38127_ (.A1(_16463_),
    .A2(_16357_),
    .B1(_16358_),
    .Y(_16464_));
 sky130_fd_sc_hd__a21oi_2 _38128_ (.A1(_16460_),
    .A2(_16462_),
    .B1(_16464_),
    .Y(_16465_));
 sky130_fd_sc_hd__nand3_2 _38129_ (.A(_16460_),
    .B(_16462_),
    .C(_16464_),
    .Y(_16466_));
 sky130_vsdinv _38130_ (.A(_16466_),
    .Y(_16467_));
 sky130_fd_sc_hd__nor2_2 _38131_ (.A(_15794_),
    .B(_16360_),
    .Y(_16468_));
 sky130_fd_sc_hd__o21bai_2 _38132_ (.A1(_16465_),
    .A2(_16467_),
    .B1_N(_16468_),
    .Y(_16469_));
 sky130_fd_sc_hd__a21o_2 _38133_ (.A1(_16460_),
    .A2(_16462_),
    .B1(_16464_),
    .X(_16470_));
 sky130_fd_sc_hd__nand3_2 _38134_ (.A(_16470_),
    .B(_16468_),
    .C(_16466_),
    .Y(_16471_));
 sky130_vsdinv _38135_ (.A(_16370_),
    .Y(_16472_));
 sky130_fd_sc_hd__o21ai_2 _38136_ (.A1(_16472_),
    .A2(_16367_),
    .B1(_16368_),
    .Y(_16473_));
 sky130_fd_sc_hd__a21oi_2 _38137_ (.A1(_16469_),
    .A2(_16471_),
    .B1(_16473_),
    .Y(_16474_));
 sky130_fd_sc_hd__nand3_2 _38138_ (.A(_16469_),
    .B(_16471_),
    .C(_16473_),
    .Y(_16475_));
 sky130_vsdinv _38139_ (.A(_16475_),
    .Y(_16476_));
 sky130_fd_sc_hd__nor2_2 _38140_ (.A(_16474_),
    .B(_16476_),
    .Y(_16477_));
 sky130_fd_sc_hd__a21oi_2 _38141_ (.A1(_16371_),
    .A2(_16373_),
    .B1(_16376_),
    .Y(_16478_));
 sky130_vsdinv _38142_ (.A(_16378_),
    .Y(_16479_));
 sky130_fd_sc_hd__o21bai_2 _38143_ (.A1(_16478_),
    .A2(_16383_),
    .B1_N(_16479_),
    .Y(_16480_));
 sky130_fd_sc_hd__xor2_2 _38144_ (.A(_16477_),
    .B(_16480_),
    .X(_02678_));
 sky130_fd_sc_hd__buf_1 _38145_ (.A(_16388_),
    .X(_16481_));
 sky130_fd_sc_hd__nor2_2 _38146_ (.A(_16389_),
    .B(_16390_),
    .Y(_16482_));
 sky130_fd_sc_hd__o21bai_2 _38147_ (.A1(_16481_),
    .A2(_16391_),
    .B1_N(_16482_),
    .Y(_16483_));
 sky130_fd_sc_hd__xnor2_2 _38148_ (.A(_16483_),
    .B(_16416_),
    .Y(_16484_));
 sky130_fd_sc_hd__xnor2_2 _38149_ (.A(_16407_),
    .B(_16484_),
    .Y(_16485_));
 sky130_fd_sc_hd__and2_2 _38150_ (.A(_16399_),
    .B(_16394_),
    .X(_16486_));
 sky130_fd_sc_hd__a21o_2 _38151_ (.A1(_16400_),
    .A2(_16392_),
    .B1(_16486_),
    .X(_16487_));
 sky130_fd_sc_hd__nand2_2 _38152_ (.A(_18714_),
    .B(_19137_),
    .Y(_16488_));
 sky130_fd_sc_hd__nand2_2 _38153_ (.A(_15981_),
    .B(_18720_),
    .Y(_16489_));
 sky130_fd_sc_hd__xnor2_2 _38154_ (.A(_16488_),
    .B(_16489_),
    .Y(_16490_));
 sky130_fd_sc_hd__xor2_2 _38155_ (.A(_16481_),
    .B(_16490_),
    .X(_16491_));
 sky130_fd_sc_hd__nor3_2 _38156_ (.A(_16067_),
    .B(_16972_),
    .C(_16396_),
    .Y(_16492_));
 sky130_fd_sc_hd__a21o_2 _38157_ (.A1(_16398_),
    .A2(_16395_),
    .B1(_16492_),
    .X(_16493_));
 sky130_fd_sc_hd__and2_2 _38158_ (.A(_18707_),
    .B(_10916_),
    .X(_16494_));
 sky130_fd_sc_hd__nand2_2 _38159_ (.A(_18698_),
    .B(_15689_),
    .Y(_16495_));
 sky130_fd_sc_hd__nand2_2 _38160_ (.A(_19152_),
    .B(_11291_),
    .Y(_16496_));
 sky130_fd_sc_hd__xor2_2 _38161_ (.A(_16495_),
    .B(_16496_),
    .X(_16497_));
 sky130_fd_sc_hd__xor2_2 _38162_ (.A(_16494_),
    .B(_16497_),
    .X(_16498_));
 sky130_fd_sc_hd__xor2_2 _38163_ (.A(_16493_),
    .B(_16498_),
    .X(_16499_));
 sky130_fd_sc_hd__xor2_2 _38164_ (.A(_16491_),
    .B(_16499_),
    .X(_16500_));
 sky130_fd_sc_hd__xnor2_2 _38165_ (.A(_16487_),
    .B(_16500_),
    .Y(_16501_));
 sky130_fd_sc_hd__xor2_2 _38166_ (.A(_16485_),
    .B(_16501_),
    .X(_16502_));
 sky130_fd_sc_hd__a21bo_2 _38167_ (.A1(_16403_),
    .A2(_16412_),
    .B1_N(_16502_),
    .X(_16503_));
 sky130_fd_sc_hd__nand3b_2 _38168_ (.A_N(_16502_),
    .B(_16403_),
    .C(_16412_),
    .Y(_16504_));
 sky130_fd_sc_hd__buf_1 _38169_ (.A(_16218_),
    .X(_16505_));
 sky130_fd_sc_hd__and2_2 _38170_ (.A(_16416_),
    .B(_16408_),
    .X(_16506_));
 sky130_fd_sc_hd__o21bai_2 _38171_ (.A1(_16407_),
    .A2(_16409_),
    .B1_N(_16506_),
    .Y(_16507_));
 sky130_fd_sc_hd__xor2_2 _38172_ (.A(_16418_),
    .B(_16507_),
    .X(_16508_));
 sky130_fd_sc_hd__xor2_2 _38173_ (.A(_16505_),
    .B(_16508_),
    .X(_16509_));
 sky130_fd_sc_hd__a21o_2 _38174_ (.A1(_16503_),
    .A2(_16504_),
    .B1(_16509_),
    .X(_16510_));
 sky130_fd_sc_hd__nand3_2 _38175_ (.A(_16503_),
    .B(_16504_),
    .C(_16509_),
    .Y(_16511_));
 sky130_fd_sc_hd__nand2_2 _38176_ (.A(_16427_),
    .B(_16413_),
    .Y(_16512_));
 sky130_fd_sc_hd__a21o_2 _38177_ (.A1(_16510_),
    .A2(_16511_),
    .B1(_16512_),
    .X(_16513_));
 sky130_fd_sc_hd__nand3_2 _38178_ (.A(_16510_),
    .B(_16511_),
    .C(_16512_),
    .Y(_16514_));
 sky130_fd_sc_hd__buf_1 _38179_ (.A(_16135_),
    .X(_16515_));
 sky130_fd_sc_hd__buf_1 _38180_ (.A(_16122_),
    .X(_16516_));
 sky130_fd_sc_hd__buf_1 _38181_ (.A(_16422_),
    .X(_16517_));
 sky130_fd_sc_hd__a21bo_2 _38182_ (.A1(_16517_),
    .A2(_16420_),
    .B1_N(_16419_),
    .X(_16518_));
 sky130_fd_sc_hd__xor2_2 _38183_ (.A(_16516_),
    .B(_16518_),
    .X(_16519_));
 sky130_fd_sc_hd__xor2_2 _38184_ (.A(_16515_),
    .B(_16519_),
    .X(_16520_));
 sky130_fd_sc_hd__a21o_2 _38185_ (.A1(_16513_),
    .A2(_16514_),
    .B1(_16520_),
    .X(_16521_));
 sky130_fd_sc_hd__nand3_2 _38186_ (.A(_16513_),
    .B(_16514_),
    .C(_16520_),
    .Y(_16522_));
 sky130_fd_sc_hd__nand2_2 _38187_ (.A(_16437_),
    .B(_16430_),
    .Y(_16523_));
 sky130_fd_sc_hd__a21o_2 _38188_ (.A1(_16521_),
    .A2(_16522_),
    .B1(_16523_),
    .X(_16524_));
 sky130_fd_sc_hd__nand3_2 _38189_ (.A(_16521_),
    .B(_16522_),
    .C(_16523_),
    .Y(_16525_));
 sky130_fd_sc_hd__buf_1 _38190_ (.A(_16247_),
    .X(_16526_));
 sky130_fd_sc_hd__a21boi_2 _38191_ (.A1(_16119_),
    .A2(_16433_),
    .B1_N(_16432_),
    .Y(_16527_));
 sky130_fd_sc_hd__xor2_2 _38192_ (.A(_16526_),
    .B(_16527_),
    .X(_16528_));
 sky130_fd_sc_hd__xor2_2 _38193_ (.A(_16458_),
    .B(_16528_),
    .X(_16529_));
 sky130_fd_sc_hd__a21oi_2 _38194_ (.A1(_16524_),
    .A2(_16525_),
    .B1(_16529_),
    .Y(_16530_));
 sky130_fd_sc_hd__nand3_2 _38195_ (.A(_16524_),
    .B(_16525_),
    .C(_16529_),
    .Y(_16531_));
 sky130_vsdinv _38196_ (.A(_16531_),
    .Y(_16532_));
 sky130_fd_sc_hd__nand2_2 _38197_ (.A(_16451_),
    .B(_16442_),
    .Y(_16533_));
 sky130_fd_sc_hd__o21bai_2 _38198_ (.A1(_16530_),
    .A2(_16532_),
    .B1_N(_16533_),
    .Y(_16534_));
 sky130_fd_sc_hd__a21o_2 _38199_ (.A1(_16524_),
    .A2(_16525_),
    .B1(_16529_),
    .X(_16535_));
 sky130_fd_sc_hd__nand3_2 _38200_ (.A(_16535_),
    .B(_16531_),
    .C(_16533_),
    .Y(_16536_));
 sky130_fd_sc_hd__a21oi_2 _38201_ (.A1(_16445_),
    .A2(_16458_),
    .B1(_16444_),
    .Y(_16537_));
 sky130_fd_sc_hd__xor2_2 _38202_ (.A(_15793_),
    .B(_16537_),
    .X(_16538_));
 sky130_fd_sc_hd__a21oi_2 _38203_ (.A1(_16534_),
    .A2(_16536_),
    .B1(_16538_),
    .Y(_16539_));
 sky130_fd_sc_hd__nand3_2 _38204_ (.A(_16534_),
    .B(_16536_),
    .C(_16538_),
    .Y(_16540_));
 sky130_fd_sc_hd__nand2_2 _38205_ (.A(_16462_),
    .B(_16453_),
    .Y(_16541_));
 sky130_fd_sc_hd__nand3b_2 _38206_ (.A_N(_16539_),
    .B(_16540_),
    .C(_16541_),
    .Y(_16542_));
 sky130_vsdinv _38207_ (.A(_16540_),
    .Y(_16543_));
 sky130_fd_sc_hd__o21bai_2 _38208_ (.A1(_16539_),
    .A2(_16543_),
    .B1_N(_16541_),
    .Y(_16544_));
 sky130_fd_sc_hd__buf_1 _38209_ (.A(_15922_),
    .X(_16545_));
 sky130_fd_sc_hd__o2bb2ai_2 _38210_ (.A1_N(_16542_),
    .A2_N(_16544_),
    .B1(_16545_),
    .B2(_16456_),
    .Y(_16546_));
 sky130_fd_sc_hd__nand3_2 _38211_ (.A(_16544_),
    .B(_16542_),
    .C(_16457_),
    .Y(_16547_));
 sky130_fd_sc_hd__a21o_2 _38212_ (.A1(_16470_),
    .A2(_16468_),
    .B1(_16467_),
    .X(_16548_));
 sky130_fd_sc_hd__a21o_2 _38213_ (.A1(_16546_),
    .A2(_16547_),
    .B1(_16548_),
    .X(_16549_));
 sky130_fd_sc_hd__nand3_2 _38214_ (.A(_16546_),
    .B(_16547_),
    .C(_16548_),
    .Y(_16550_));
 sky130_fd_sc_hd__nand2_2 _38215_ (.A(_16549_),
    .B(_16550_),
    .Y(_16551_));
 sky130_fd_sc_hd__nor2_2 _38216_ (.A(_16169_),
    .B(_16283_),
    .Y(_16552_));
 sky130_fd_sc_hd__a21o_2 _38217_ (.A1(_16469_),
    .A2(_16471_),
    .B1(_16473_),
    .X(_16553_));
 sky130_fd_sc_hd__nand2_2 _38218_ (.A(_16553_),
    .B(_16475_),
    .Y(_16554_));
 sky130_fd_sc_hd__nor2_2 _38219_ (.A(_16379_),
    .B(_16554_),
    .Y(_16555_));
 sky130_fd_sc_hd__nand2_2 _38220_ (.A(_16552_),
    .B(_16555_),
    .Y(_16556_));
 sky130_fd_sc_hd__nor2_2 _38221_ (.A(_16478_),
    .B(_16479_),
    .Y(_16557_));
 sky130_fd_sc_hd__nand3_2 _38222_ (.A(_16477_),
    .B(_16381_),
    .C(_16557_),
    .Y(_16558_));
 sky130_fd_sc_hd__a21oi_2 _38223_ (.A1(_16553_),
    .A2(_16479_),
    .B1(_16476_),
    .Y(_16559_));
 sky130_fd_sc_hd__nand2_2 _38224_ (.A(_16558_),
    .B(_16559_),
    .Y(_16560_));
 sky130_fd_sc_hd__o21bai_2 _38225_ (.A1(_16556_),
    .A2(_16176_),
    .B1_N(_16560_),
    .Y(_16561_));
 sky130_fd_sc_hd__xnor2_2 _38226_ (.A(_16551_),
    .B(_16561_),
    .Y(_02679_));
 sky130_fd_sc_hd__nand2_2 _38227_ (.A(_16522_),
    .B(_16514_),
    .Y(_16562_));
 sky130_fd_sc_hd__buf_1 _38228_ (.A(_16406_),
    .X(_16563_));
 sky130_fd_sc_hd__buf_1 _38229_ (.A(_16309_),
    .X(_16564_));
 sky130_fd_sc_hd__and2_2 _38230_ (.A(_16564_),
    .B(_16483_),
    .X(_16565_));
 sky130_fd_sc_hd__o21bai_2 _38231_ (.A1(_16563_),
    .A2(_16484_),
    .B1_N(_16565_),
    .Y(_16566_));
 sky130_fd_sc_hd__xor2_2 _38232_ (.A(_16418_),
    .B(_16566_),
    .X(_16567_));
 sky130_fd_sc_hd__xor2_2 _38233_ (.A(_16517_),
    .B(_16567_),
    .X(_16568_));
 sky130_fd_sc_hd__nand2_2 _38234_ (.A(_16500_),
    .B(_16487_),
    .Y(_16569_));
 sky130_fd_sc_hd__o21ai_2 _38235_ (.A1(_16485_),
    .A2(_16501_),
    .B1(_16569_),
    .Y(_16570_));
 sky130_fd_sc_hd__nor2_2 _38236_ (.A(_16488_),
    .B(_16489_),
    .Y(_16571_));
 sky130_fd_sc_hd__o21ba_2 _38237_ (.A1(_16481_),
    .A2(_16490_),
    .B1_N(_16571_),
    .X(_16572_));
 sky130_fd_sc_hd__xor2_2 _38238_ (.A(_16572_),
    .B(_16564_),
    .X(_16573_));
 sky130_fd_sc_hd__xnor2_2 _38239_ (.A(_16407_),
    .B(_16573_),
    .Y(_16574_));
 sky130_fd_sc_hd__and2_2 _38240_ (.A(_16498_),
    .B(_16493_),
    .X(_16575_));
 sky130_fd_sc_hd__a21o_2 _38241_ (.A1(_16499_),
    .A2(_16491_),
    .B1(_16575_),
    .X(_16576_));
 sky130_fd_sc_hd__nand2_2 _38242_ (.A(_15981_),
    .B(_16066_),
    .Y(_16577_));
 sky130_fd_sc_hd__xnor2_2 _38243_ (.A(_16489_),
    .B(_16577_),
    .Y(_16578_));
 sky130_fd_sc_hd__xor2_2 _38244_ (.A(_16388_),
    .B(_16578_),
    .X(_16579_));
 sky130_fd_sc_hd__nor3_2 _38245_ (.A(_15827_),
    .B(_16972_),
    .C(_16495_),
    .Y(_16580_));
 sky130_fd_sc_hd__a21o_2 _38246_ (.A1(_16497_),
    .A2(_16494_),
    .B1(_16580_),
    .X(_16581_));
 sky130_fd_sc_hd__and2_2 _38247_ (.A(_18707_),
    .B(_19136_),
    .X(_16582_));
 sky130_fd_sc_hd__nand2_2 _38248_ (.A(_18697_),
    .B(_16179_),
    .Y(_16583_));
 sky130_fd_sc_hd__nand2_2 _38249_ (.A(_19147_),
    .B(_11290_),
    .Y(_16584_));
 sky130_fd_sc_hd__xor2_2 _38250_ (.A(_16583_),
    .B(_16584_),
    .X(_16585_));
 sky130_fd_sc_hd__xor2_2 _38251_ (.A(_16582_),
    .B(_16585_),
    .X(_16586_));
 sky130_fd_sc_hd__xor2_2 _38252_ (.A(_16581_),
    .B(_16586_),
    .X(_16587_));
 sky130_fd_sc_hd__xor2_2 _38253_ (.A(_16579_),
    .B(_16587_),
    .X(_16588_));
 sky130_fd_sc_hd__xnor2_2 _38254_ (.A(_16576_),
    .B(_16588_),
    .Y(_16589_));
 sky130_fd_sc_hd__xor2_2 _38255_ (.A(_16574_),
    .B(_16589_),
    .X(_16590_));
 sky130_fd_sc_hd__xnor2_2 _38256_ (.A(_16570_),
    .B(_16590_),
    .Y(_16591_));
 sky130_fd_sc_hd__nor2_2 _38257_ (.A(_16568_),
    .B(_16591_),
    .Y(_16592_));
 sky130_fd_sc_hd__nand2_2 _38258_ (.A(_16591_),
    .B(_16568_),
    .Y(_16593_));
 sky130_vsdinv _38259_ (.A(_16593_),
    .Y(_16594_));
 sky130_fd_sc_hd__nand2_2 _38260_ (.A(_16511_),
    .B(_16503_),
    .Y(_16595_));
 sky130_fd_sc_hd__o21bai_2 _38261_ (.A1(_16592_),
    .A2(_16594_),
    .B1_N(_16595_),
    .Y(_16596_));
 sky130_fd_sc_hd__nand3b_2 _38262_ (.A_N(_16592_),
    .B(_16595_),
    .C(_16593_),
    .Y(_16597_));
 sky130_fd_sc_hd__or2b_2 _38263_ (.A(_16508_),
    .B_N(_16517_),
    .X(_16598_));
 sky130_fd_sc_hd__nand2_2 _38264_ (.A(_16507_),
    .B(_16107_),
    .Y(_16599_));
 sky130_fd_sc_hd__a21o_2 _38265_ (.A1(_16598_),
    .A2(_16599_),
    .B1(_16516_),
    .X(_16600_));
 sky130_fd_sc_hd__o211ai_2 _38266_ (.A1(_16505_),
    .A2(_16508_),
    .B1(_16516_),
    .C1(_16599_),
    .Y(_16601_));
 sky130_fd_sc_hd__nand2_2 _38267_ (.A(_16600_),
    .B(_16601_),
    .Y(_16602_));
 sky130_fd_sc_hd__xor2_2 _38268_ (.A(_16515_),
    .B(_16602_),
    .X(_16603_));
 sky130_fd_sc_hd__a21o_2 _38269_ (.A1(_16596_),
    .A2(_16597_),
    .B1(_16603_),
    .X(_16604_));
 sky130_fd_sc_hd__nand3_2 _38270_ (.A(_16596_),
    .B(_16597_),
    .C(_16603_),
    .Y(_16605_));
 sky130_fd_sc_hd__nand3_2 _38271_ (.A(_16562_),
    .B(_16604_),
    .C(_16605_),
    .Y(_16606_));
 sky130_fd_sc_hd__a21o_2 _38272_ (.A1(_16604_),
    .A2(_16605_),
    .B1(_16562_),
    .X(_16607_));
 sky130_fd_sc_hd__buf_1 _38273_ (.A(_16149_),
    .X(_16608_));
 sky130_fd_sc_hd__and2_2 _38274_ (.A(_16518_),
    .B(_15875_),
    .X(_16609_));
 sky130_fd_sc_hd__o21ba_2 _38275_ (.A1(_16135_),
    .A2(_16519_),
    .B1_N(_16609_),
    .X(_16610_));
 sky130_fd_sc_hd__nor2_2 _38276_ (.A(_16526_),
    .B(_16610_),
    .Y(_16611_));
 sky130_fd_sc_hd__o21a_2 _38277_ (.A1(_15135_),
    .A2(_15137_),
    .B1(_16610_),
    .X(_16612_));
 sky130_fd_sc_hd__nor3_2 _38278_ (.A(_16608_),
    .B(_16611_),
    .C(_16612_),
    .Y(_16613_));
 sky130_fd_sc_hd__o21a_2 _38279_ (.A1(_16611_),
    .A2(_16612_),
    .B1(_16149_),
    .X(_16614_));
 sky130_fd_sc_hd__o2bb2ai_2 _38280_ (.A1_N(_16606_),
    .A2_N(_16607_),
    .B1(_16613_),
    .B2(_16614_),
    .Y(_16615_));
 sky130_fd_sc_hd__nor2_2 _38281_ (.A(_16613_),
    .B(_16614_),
    .Y(_16616_));
 sky130_fd_sc_hd__nand3_2 _38282_ (.A(_16607_),
    .B(_16606_),
    .C(_16616_),
    .Y(_16617_));
 sky130_fd_sc_hd__and3_2 _38283_ (.A(_16521_),
    .B(_16522_),
    .C(_16523_),
    .X(_16618_));
 sky130_fd_sc_hd__a21o_2 _38284_ (.A1(_16524_),
    .A2(_16529_),
    .B1(_16618_),
    .X(_16619_));
 sky130_fd_sc_hd__a21o_2 _38285_ (.A1(_16615_),
    .A2(_16617_),
    .B1(_16619_),
    .X(_16620_));
 sky130_fd_sc_hd__nand3_2 _38286_ (.A(_16619_),
    .B(_16617_),
    .C(_16615_),
    .Y(_16621_));
 sky130_fd_sc_hd__buf_1 _38287_ (.A(_16621_),
    .X(_16622_));
 sky130_fd_sc_hd__nor2_2 _38288_ (.A(_16526_),
    .B(_16527_),
    .Y(_16623_));
 sky130_fd_sc_hd__a21oi_2 _38289_ (.A1(_16528_),
    .A2(_16458_),
    .B1(_16623_),
    .Y(_16624_));
 sky130_fd_sc_hd__xor2_2 _38290_ (.A(_15793_),
    .B(_16624_),
    .X(_16625_));
 sky130_fd_sc_hd__a21oi_2 _38291_ (.A1(_16620_),
    .A2(_16622_),
    .B1(_16625_),
    .Y(_16626_));
 sky130_vsdinv _38292_ (.A(_16625_),
    .Y(_16627_));
 sky130_fd_sc_hd__a21oi_2 _38293_ (.A1(_16615_),
    .A2(_16617_),
    .B1(_16619_),
    .Y(_16628_));
 sky130_fd_sc_hd__nor3b_2 _38294_ (.A(_16627_),
    .B(_16628_),
    .C_N(_16621_),
    .Y(_16629_));
 sky130_vsdinv _38295_ (.A(_16538_),
    .Y(_16630_));
 sky130_fd_sc_hd__a21oi_2 _38296_ (.A1(_16535_),
    .A2(_16531_),
    .B1(_16533_),
    .Y(_16631_));
 sky130_fd_sc_hd__o21ai_2 _38297_ (.A1(_16630_),
    .A2(_16631_),
    .B1(_16536_),
    .Y(_16632_));
 sky130_fd_sc_hd__o21bai_2 _38298_ (.A1(_16626_),
    .A2(_16629_),
    .B1_N(_16632_),
    .Y(_16633_));
 sky130_fd_sc_hd__a21o_2 _38299_ (.A1(_16620_),
    .A2(_16622_),
    .B1(_16625_),
    .X(_16634_));
 sky130_fd_sc_hd__nand3_2 _38300_ (.A(_16620_),
    .B(_16622_),
    .C(_16625_),
    .Y(_16635_));
 sky130_fd_sc_hd__nand3_2 _38301_ (.A(_16634_),
    .B(_16632_),
    .C(_16635_),
    .Y(_16636_));
 sky130_fd_sc_hd__nor2_2 _38302_ (.A(_15922_),
    .B(_16537_),
    .Y(_16637_));
 sky130_fd_sc_hd__a21oi_2 _38303_ (.A1(_16633_),
    .A2(_16636_),
    .B1(_16637_),
    .Y(_16638_));
 sky130_fd_sc_hd__nand3_2 _38304_ (.A(_16633_),
    .B(_16637_),
    .C(_16636_),
    .Y(_16639_));
 sky130_vsdinv _38305_ (.A(_16639_),
    .Y(_16640_));
 sky130_fd_sc_hd__a21boi_2 _38306_ (.A1(_16544_),
    .A2(_16457_),
    .B1_N(_16542_),
    .Y(_16641_));
 sky130_fd_sc_hd__o21ai_2 _38307_ (.A1(_16638_),
    .A2(_16640_),
    .B1(_16641_),
    .Y(_16642_));
 sky130_fd_sc_hd__nand2_2 _38308_ (.A(_16547_),
    .B(_16542_),
    .Y(_16643_));
 sky130_fd_sc_hd__o2bb2ai_2 _38309_ (.A1_N(_16636_),
    .A2_N(_16633_),
    .B1(_16545_),
    .B2(_16537_),
    .Y(_16644_));
 sky130_fd_sc_hd__nand3_2 _38310_ (.A(_16643_),
    .B(_16644_),
    .C(_16639_),
    .Y(_16645_));
 sky130_fd_sc_hd__nand2_2 _38311_ (.A(_16642_),
    .B(_16645_),
    .Y(_16646_));
 sky130_fd_sc_hd__a21boi_2 _38312_ (.A1(_16561_),
    .A2(_16549_),
    .B1_N(_16550_),
    .Y(_16647_));
 sky130_fd_sc_hd__xor2_2 _38313_ (.A(_16646_),
    .B(_16647_),
    .X(_02680_));
 sky130_fd_sc_hd__a21boi_2 _38314_ (.A1(_16596_),
    .A2(_16603_),
    .B1_N(_16597_),
    .Y(_16648_));
 sky130_fd_sc_hd__nand2_2 _38315_ (.A(_16566_),
    .B(_16107_),
    .Y(_16649_));
 sky130_fd_sc_hd__o21a_2 _38316_ (.A1(_16505_),
    .A2(_16567_),
    .B1(_16649_),
    .X(_16650_));
 sky130_fd_sc_hd__xor2_2 _38317_ (.A(_15875_),
    .B(_16650_),
    .X(_16651_));
 sky130_fd_sc_hd__xor2_2 _38318_ (.A(_16515_),
    .B(_16651_),
    .X(_16652_));
 sky130_vsdinv _38319_ (.A(_16652_),
    .Y(_16653_));
 sky130_fd_sc_hd__or2b_2 _38320_ (.A(_16572_),
    .B_N(_16564_),
    .X(_16654_));
 sky130_fd_sc_hd__o21a_2 _38321_ (.A1(_16563_),
    .A2(_16573_),
    .B1(_16654_),
    .X(_16655_));
 sky130_fd_sc_hd__xor2_2 _38322_ (.A(_16107_),
    .B(_16655_),
    .X(_16656_));
 sky130_fd_sc_hd__xor2_2 _38323_ (.A(_16517_),
    .B(_16656_),
    .X(_16657_));
 sky130_fd_sc_hd__nand2_2 _38324_ (.A(_16588_),
    .B(_16576_),
    .Y(_16658_));
 sky130_fd_sc_hd__o21ai_2 _38325_ (.A1(_16574_),
    .A2(_16589_),
    .B1(_16658_),
    .Y(_16659_));
 sky130_fd_sc_hd__nor2_2 _38326_ (.A(_16481_),
    .B(_16578_),
    .Y(_16660_));
 sky130_fd_sc_hd__o21bai_2 _38327_ (.A1(_16489_),
    .A2(_16577_),
    .B1_N(_16660_),
    .Y(_16661_));
 sky130_fd_sc_hd__xnor2_2 _38328_ (.A(_16416_),
    .B(_16661_),
    .Y(_16662_));
 sky130_fd_sc_hd__xnor2_2 _38329_ (.A(_16563_),
    .B(_16662_),
    .Y(_16663_));
 sky130_fd_sc_hd__buf_1 _38330_ (.A(_16579_),
    .X(_16664_));
 sky130_fd_sc_hd__and2_2 _38331_ (.A(_16586_),
    .B(_16581_),
    .X(_16665_));
 sky130_fd_sc_hd__a21o_2 _38332_ (.A1(_16587_),
    .A2(_16664_),
    .B1(_16665_),
    .X(_16666_));
 sky130_fd_sc_hd__nor3_2 _38333_ (.A(_16064_),
    .B(_16973_),
    .C(_16583_),
    .Y(_16667_));
 sky130_fd_sc_hd__a21o_2 _38334_ (.A1(_16585_),
    .A2(_16582_),
    .B1(_16667_),
    .X(_16668_));
 sky130_fd_sc_hd__and2_2 _38335_ (.A(_16387_),
    .B(_18707_),
    .X(_16669_));
 sky130_fd_sc_hd__nand2_2 _38336_ (.A(_18698_),
    .B(_19135_),
    .Y(_16670_));
 sky130_fd_sc_hd__nand2_2 _38337_ (.A(_19141_),
    .B(_11291_),
    .Y(_16671_));
 sky130_fd_sc_hd__xor2_2 _38338_ (.A(_16670_),
    .B(_16671_),
    .X(_16672_));
 sky130_fd_sc_hd__xor2_2 _38339_ (.A(_16669_),
    .B(_16672_),
    .X(_16673_));
 sky130_fd_sc_hd__xor2_2 _38340_ (.A(_16668_),
    .B(_16673_),
    .X(_16674_));
 sky130_fd_sc_hd__xor2_2 _38341_ (.A(_16664_),
    .B(_16674_),
    .X(_16675_));
 sky130_fd_sc_hd__xnor2_2 _38342_ (.A(_16666_),
    .B(_16675_),
    .Y(_16676_));
 sky130_fd_sc_hd__xor2_2 _38343_ (.A(_16663_),
    .B(_16676_),
    .X(_16677_));
 sky130_fd_sc_hd__xnor2_2 _38344_ (.A(_16659_),
    .B(_16677_),
    .Y(_16678_));
 sky130_fd_sc_hd__xor2_2 _38345_ (.A(_16657_),
    .B(_16678_),
    .X(_16679_));
 sky130_fd_sc_hd__a21o_2 _38346_ (.A1(_16590_),
    .A2(_16570_),
    .B1(_16592_),
    .X(_16680_));
 sky130_fd_sc_hd__xnor2_2 _38347_ (.A(_16679_),
    .B(_16680_),
    .Y(_16681_));
 sky130_fd_sc_hd__nor2_2 _38348_ (.A(_16653_),
    .B(_16681_),
    .Y(_16682_));
 sky130_fd_sc_hd__and2_2 _38349_ (.A(_16681_),
    .B(_16653_),
    .X(_16683_));
 sky130_fd_sc_hd__nor3_2 _38350_ (.A(_16648_),
    .B(_16682_),
    .C(_16683_),
    .Y(_16684_));
 sky130_vsdinv _38351_ (.A(_16684_),
    .Y(_16685_));
 sky130_fd_sc_hd__o21ai_2 _38352_ (.A1(_16682_),
    .A2(_16683_),
    .B1(_16648_),
    .Y(_16686_));
 sky130_fd_sc_hd__a21boi_2 _38353_ (.A1(_16119_),
    .A2(_16601_),
    .B1_N(_16600_),
    .Y(_16687_));
 sky130_fd_sc_hd__xor2_2 _38354_ (.A(_15138_),
    .B(_16687_),
    .X(_16688_));
 sky130_fd_sc_hd__xor2_2 _38355_ (.A(_16608_),
    .B(_16688_),
    .X(_16689_));
 sky130_fd_sc_hd__a21oi_2 _38356_ (.A1(_16685_),
    .A2(_16686_),
    .B1(_16689_),
    .Y(_16690_));
 sky130_fd_sc_hd__nand3b_2 _38357_ (.A_N(_16684_),
    .B(_16686_),
    .C(_16689_),
    .Y(_16691_));
 sky130_vsdinv _38358_ (.A(_16691_),
    .Y(_16692_));
 sky130_fd_sc_hd__nand2_2 _38359_ (.A(_16617_),
    .B(_16606_),
    .Y(_16693_));
 sky130_fd_sc_hd__o21bai_2 _38360_ (.A1(_16690_),
    .A2(_16692_),
    .B1_N(_16693_),
    .Y(_16694_));
 sky130_fd_sc_hd__a21o_2 _38361_ (.A1(_16685_),
    .A2(_16686_),
    .B1(_16689_),
    .X(_16695_));
 sky130_fd_sc_hd__nand3_2 _38362_ (.A(_16695_),
    .B(_16691_),
    .C(_16693_),
    .Y(_16696_));
 sky130_fd_sc_hd__buf_1 _38363_ (.A(_16696_),
    .X(_16697_));
 sky130_fd_sc_hd__o21ba_2 _38364_ (.A1(_16608_),
    .A2(_16612_),
    .B1_N(_16611_),
    .X(_16698_));
 sky130_fd_sc_hd__xor2_2 _38365_ (.A(_16040_),
    .B(_16698_),
    .X(_16699_));
 sky130_fd_sc_hd__a21boi_2 _38366_ (.A1(_16694_),
    .A2(_16697_),
    .B1_N(_16699_),
    .Y(_16700_));
 sky130_fd_sc_hd__nand3b_2 _38367_ (.A_N(_16699_),
    .B(_16694_),
    .C(_16696_),
    .Y(_16701_));
 sky130_vsdinv _38368_ (.A(_16701_),
    .Y(_16702_));
 sky130_fd_sc_hd__o21ai_2 _38369_ (.A1(_16627_),
    .A2(_16628_),
    .B1(_16622_),
    .Y(_16703_));
 sky130_fd_sc_hd__o21bai_2 _38370_ (.A1(_16700_),
    .A2(_16702_),
    .B1_N(_16703_),
    .Y(_16704_));
 sky130_fd_sc_hd__a21bo_2 _38371_ (.A1(_16694_),
    .A2(_16697_),
    .B1_N(_16699_),
    .X(_16705_));
 sky130_fd_sc_hd__nand3_2 _38372_ (.A(_16705_),
    .B(_16701_),
    .C(_16703_),
    .Y(_16706_));
 sky130_fd_sc_hd__buf_1 _38373_ (.A(_16706_),
    .X(_16707_));
 sky130_fd_sc_hd__nor2_2 _38374_ (.A(_16545_),
    .B(_16624_),
    .Y(_16708_));
 sky130_fd_sc_hd__a21oi_2 _38375_ (.A1(_16704_),
    .A2(_16707_),
    .B1(_16708_),
    .Y(_16709_));
 sky130_fd_sc_hd__nand3_2 _38376_ (.A(_16704_),
    .B(_16708_),
    .C(_16706_),
    .Y(_16710_));
 sky130_vsdinv _38377_ (.A(_16710_),
    .Y(_16711_));
 sky130_fd_sc_hd__nand2_2 _38378_ (.A(_16639_),
    .B(_16636_),
    .Y(_16712_));
 sky130_fd_sc_hd__o21bai_2 _38379_ (.A1(_16709_),
    .A2(_16711_),
    .B1_N(_16712_),
    .Y(_16713_));
 sky130_fd_sc_hd__o2bb2ai_2 _38380_ (.A1_N(_16707_),
    .A2_N(_16704_),
    .B1(_16545_),
    .B2(_16624_),
    .Y(_16714_));
 sky130_fd_sc_hd__nand3_2 _38381_ (.A(_16714_),
    .B(_16710_),
    .C(_16712_),
    .Y(_16715_));
 sky130_fd_sc_hd__nand2_2 _38382_ (.A(_16713_),
    .B(_16715_),
    .Y(_16716_));
 sky130_fd_sc_hd__nor2_2 _38383_ (.A(_16646_),
    .B(_16551_),
    .Y(_16717_));
 sky130_fd_sc_hd__nand2_2 _38384_ (.A(_16561_),
    .B(_16717_),
    .Y(_16718_));
 sky130_fd_sc_hd__a21boi_2 _38385_ (.A1(_16550_),
    .A2(_16645_),
    .B1_N(_16642_),
    .Y(_16719_));
 sky130_vsdinv _38386_ (.A(_16719_),
    .Y(_16720_));
 sky130_fd_sc_hd__nand2_2 _38387_ (.A(_16718_),
    .B(_16720_),
    .Y(_16721_));
 sky130_fd_sc_hd__xnor2_2 _38388_ (.A(_16716_),
    .B(_16721_),
    .Y(_02681_));
 sky130_vsdinv _38389_ (.A(_16715_),
    .Y(_16722_));
 sky130_fd_sc_hd__a21oi_2 _38390_ (.A1(_16695_),
    .A2(_16691_),
    .B1(_16693_),
    .Y(_16723_));
 sky130_fd_sc_hd__o21ai_2 _38391_ (.A1(_16699_),
    .A2(_16723_),
    .B1(_16697_),
    .Y(_16724_));
 sky130_fd_sc_hd__nor2_2 _38392_ (.A(_16526_),
    .B(_16687_),
    .Y(_16725_));
 sky130_fd_sc_hd__o21ba_2 _38393_ (.A1(_16608_),
    .A2(_16688_),
    .B1_N(_16725_),
    .X(_16726_));
 sky130_fd_sc_hd__nand2_2 _38394_ (.A(_16724_),
    .B(_16726_),
    .Y(_16727_));
 sky130_fd_sc_hd__nand3b_2 _38395_ (.A_N(_16726_),
    .B(_16701_),
    .C(_16697_),
    .Y(_16728_));
 sky130_fd_sc_hd__nand2_2 _38396_ (.A(_16727_),
    .B(_16728_),
    .Y(_16729_));
 sky130_fd_sc_hd__and2b_2 _38397_ (.A_N(_14955_),
    .B(_15134_),
    .X(_16730_));
 sky130_fd_sc_hd__a21oi_2 _38398_ (.A1(_15136_),
    .A2(_14955_),
    .B1(_16730_),
    .Y(_16731_));
 sky130_fd_sc_hd__nand2_2 _38399_ (.A(_16729_),
    .B(_16731_),
    .Y(_16732_));
 sky130_fd_sc_hd__nand3b_2 _38400_ (.A_N(_16731_),
    .B(_16727_),
    .C(_16728_),
    .Y(_16733_));
 sky130_fd_sc_hd__nand2_2 _38401_ (.A(_16698_),
    .B(_16040_),
    .Y(_16734_));
 sky130_fd_sc_hd__a21o_2 _38402_ (.A1(_16732_),
    .A2(_16733_),
    .B1(_16734_),
    .X(_16735_));
 sky130_fd_sc_hd__nand3_2 _38403_ (.A(_16732_),
    .B(_16734_),
    .C(_16733_),
    .Y(_16736_));
 sky130_fd_sc_hd__nand2_2 _38404_ (.A(_16735_),
    .B(_16736_),
    .Y(_16737_));
 sky130_vsdinv _38405_ (.A(_15880_),
    .Y(_16738_));
 sky130_fd_sc_hd__mux2_2 _38406_ (.A0(_15873_),
    .A1(_16738_),
    .S(_14849_),
    .X(_16739_));
 sky130_fd_sc_hd__nor2_2 _38407_ (.A(_16516_),
    .B(_16650_),
    .Y(_16740_));
 sky130_fd_sc_hd__o21bai_2 _38408_ (.A1(_16515_),
    .A2(_16651_),
    .B1_N(_16740_),
    .Y(_16741_));
 sky130_fd_sc_hd__xnor2_2 _38409_ (.A(_16739_),
    .B(_16741_),
    .Y(_16742_));
 sky130_fd_sc_hd__a21o_2 _38410_ (.A1(_16679_),
    .A2(_16680_),
    .B1(_16682_),
    .X(_16743_));
 sky130_fd_sc_hd__mux2_2 _38411_ (.A0(_16104_),
    .A1(_16102_),
    .S(_15995_),
    .X(_16744_));
 sky130_fd_sc_hd__nor2_2 _38412_ (.A(_16418_),
    .B(_16655_),
    .Y(_16745_));
 sky130_fd_sc_hd__o21bai_2 _38413_ (.A1(_16505_),
    .A2(_16656_),
    .B1_N(_16745_),
    .Y(_16746_));
 sky130_fd_sc_hd__xor2_2 _38414_ (.A(_16744_),
    .B(_16746_),
    .X(_16747_));
 sky130_fd_sc_hd__and2_2 _38415_ (.A(_16677_),
    .B(_16659_),
    .X(_16748_));
 sky130_fd_sc_hd__o21bai_2 _38416_ (.A1(_16657_),
    .A2(_16678_),
    .B1_N(_16748_),
    .Y(_16749_));
 sky130_fd_sc_hd__and2_2 _38417_ (.A(_16387_),
    .B(_18698_),
    .X(_16750_));
 sky130_fd_sc_hd__and2_2 _38418_ (.A(_16673_),
    .B(_16668_),
    .X(_16751_));
 sky130_fd_sc_hd__a21oi_2 _38419_ (.A1(_16674_),
    .A2(_16664_),
    .B1(_16751_),
    .Y(_16752_));
 sky130_fd_sc_hd__xor2_2 _38420_ (.A(_16750_),
    .B(_16752_),
    .X(_16753_));
 sky130_fd_sc_hd__xnor2_2 _38421_ (.A(_16669_),
    .B(_16664_),
    .Y(_16754_));
 sky130_fd_sc_hd__and2b_2 _38422_ (.A_N(_19137_),
    .B(_11291_),
    .X(_16755_));
 sky130_fd_sc_hd__xor2_2 _38423_ (.A(_16755_),
    .B(_16663_),
    .X(_16756_));
 sky130_fd_sc_hd__xor2_2 _38424_ (.A(_16754_),
    .B(_16756_),
    .X(_16757_));
 sky130_fd_sc_hd__xor2_2 _38425_ (.A(_16753_),
    .B(_16757_),
    .X(_16758_));
 sky130_fd_sc_hd__nor2_2 _38426_ (.A(_16563_),
    .B(_16662_),
    .Y(_16759_));
 sky130_fd_sc_hd__a21oi_2 _38427_ (.A1(_16564_),
    .A2(_16661_),
    .B1(_16759_),
    .Y(_16760_));
 sky130_fd_sc_hd__nor3_2 _38428_ (.A(_10916_),
    .B(_16973_),
    .C(_16670_),
    .Y(_16761_));
 sky130_fd_sc_hd__a21o_2 _38429_ (.A1(_16672_),
    .A2(_16669_),
    .B1(_16761_),
    .X(_16762_));
 sky130_fd_sc_hd__nand2_2 _38430_ (.A(_16675_),
    .B(_16666_),
    .Y(_16763_));
 sky130_fd_sc_hd__o21ai_2 _38431_ (.A1(_16663_),
    .A2(_16676_),
    .B1(_16763_),
    .Y(_16764_));
 sky130_fd_sc_hd__xor2_2 _38432_ (.A(_16762_),
    .B(_16764_),
    .X(_16765_));
 sky130_fd_sc_hd__xor2_2 _38433_ (.A(_16760_),
    .B(_16765_),
    .X(_16766_));
 sky130_fd_sc_hd__xor2_2 _38434_ (.A(_16758_),
    .B(_16766_),
    .X(_16767_));
 sky130_fd_sc_hd__xor2_2 _38435_ (.A(_16749_),
    .B(_16767_),
    .X(_16768_));
 sky130_fd_sc_hd__xor2_2 _38436_ (.A(_16747_),
    .B(_16768_),
    .X(_16769_));
 sky130_fd_sc_hd__xor2_2 _38437_ (.A(_16743_),
    .B(_16769_),
    .X(_16770_));
 sky130_fd_sc_hd__nor2_2 _38438_ (.A(_16742_),
    .B(_16770_),
    .Y(_16771_));
 sky130_fd_sc_hd__and2_2 _38439_ (.A(_16770_),
    .B(_16742_),
    .X(_16772_));
 sky130_fd_sc_hd__a21oi_2 _38440_ (.A1(_16686_),
    .A2(_16689_),
    .B1(_16684_),
    .Y(_16773_));
 sky130_fd_sc_hd__o21a_2 _38441_ (.A1(_16771_),
    .A2(_16772_),
    .B1(_16773_),
    .X(_16774_));
 sky130_fd_sc_hd__nor3_2 _38442_ (.A(_16773_),
    .B(_16771_),
    .C(_16772_),
    .Y(_16775_));
 sky130_vsdinv _38443_ (.A(_16708_),
    .Y(_16776_));
 sky130_fd_sc_hd__a21oi_2 _38444_ (.A1(_16705_),
    .A2(_16701_),
    .B1(_16703_),
    .Y(_16777_));
 sky130_fd_sc_hd__o221ai_2 _38445_ (.A1(_16774_),
    .A2(_16775_),
    .B1(_16776_),
    .B2(_16777_),
    .C1(_16707_),
    .Y(_16778_));
 sky130_fd_sc_hd__o21ai_2 _38446_ (.A1(_16776_),
    .A2(_16777_),
    .B1(_16707_),
    .Y(_16779_));
 sky130_fd_sc_hd__nor2_2 _38447_ (.A(_16775_),
    .B(_16774_),
    .Y(_16780_));
 sky130_fd_sc_hd__nand2_2 _38448_ (.A(_16779_),
    .B(_16780_),
    .Y(_16781_));
 sky130_fd_sc_hd__nand3_2 _38449_ (.A(_16737_),
    .B(_16778_),
    .C(_16781_),
    .Y(_16782_));
 sky130_fd_sc_hd__nand2_2 _38450_ (.A(_16781_),
    .B(_16778_),
    .Y(_16783_));
 sky130_fd_sc_hd__nand3_2 _38451_ (.A(_16783_),
    .B(_16735_),
    .C(_16736_),
    .Y(_16784_));
 sky130_fd_sc_hd__nand2_2 _38452_ (.A(_16782_),
    .B(_16784_),
    .Y(_16785_));
 sky130_fd_sc_hd__a21oi_2 _38453_ (.A1(_16718_),
    .A2(_16720_),
    .B1(_16716_),
    .Y(_16786_));
 sky130_fd_sc_hd__nor3_2 _38454_ (.A(_16722_),
    .B(_16785_),
    .C(_16786_),
    .Y(_16787_));
 sky130_vsdinv _38455_ (.A(_16716_),
    .Y(_16788_));
 sky130_fd_sc_hd__nand2_2 _38456_ (.A(_16721_),
    .B(_16788_),
    .Y(_16789_));
 sky130_vsdinv _38457_ (.A(_16785_),
    .Y(_16790_));
 sky130_fd_sc_hd__a21oi_2 _38458_ (.A1(_16789_),
    .A2(_16715_),
    .B1(_16790_),
    .Y(_16791_));
 sky130_fd_sc_hd__nor2_2 _38459_ (.A(_16787_),
    .B(_16791_),
    .Y(_02682_));
 sky130_fd_sc_hd__nand2_2 _38460_ (.A(_05627_),
    .B(_05618_),
    .Y(_16792_));
 sky130_fd_sc_hd__o21bai_2 _38461_ (.A1(_05487_),
    .A2(_05488_),
    .B1_N(_05486_),
    .Y(_16793_));
 sky130_fd_sc_hd__xnor2_2 _38462_ (.A(_16792_),
    .B(_16793_),
    .Y(_02628_));
 sky130_fd_sc_hd__and4_2 _38463_ (.A(_02321_),
    .B(_02318_),
    .C(_05247_),
    .D(_19124_),
    .X(_00050_));
 sky130_fd_sc_hd__nor3b_2 _38464_ (.A(_05168_),
    .B(_18527_),
    .C_N(_00066_),
    .Y(_00068_));
 sky130_fd_sc_hd__nor2b_2 _38465_ (.A(_05168_),
    .B_N(_00084_),
    .Y(_00085_));
 sky130_fd_sc_hd__nor2b_2 _38466_ (.A(_05168_),
    .B_N(_00094_),
    .Y(_00095_));
 sky130_fd_sc_hd__o21a_2 _38467_ (.A1(instr_sra),
    .A2(instr_srai),
    .B1(_16958_),
    .X(_00216_));
 sky130_fd_sc_hd__o21a_2 _38468_ (.A1(_04292_),
    .A2(_17044_),
    .B1(_00321_),
    .X(_16794_));
 sky130_fd_sc_hd__o211ai_2 _38469_ (.A1(_17038_),
    .A2(_17403_),
    .B1(_19773_),
    .C1(_00321_),
    .Y(_16795_));
 sky130_fd_sc_hd__o211a_2 _38470_ (.A1(_16936_),
    .A2(_16794_),
    .B1(_17998_),
    .C1(_16795_),
    .X(_04072_));
 sky130_fd_sc_hd__conb_1 _38471_ (.LO(mem_addr[0]));
 sky130_fd_sc_hd__conb_1 _38472_ (.LO(mem_addr[1]));
 sky130_fd_sc_hd__conb_1 _38473_ (.LO(mem_la_addr[0]));
 sky130_fd_sc_hd__conb_1 _38474_ (.LO(mem_la_addr[1]));
 sky130_fd_sc_hd__conb_1 _38475_ (.LO(trace_data[0]));
 sky130_fd_sc_hd__conb_1 _38476_ (.LO(trace_data[1]));
 sky130_fd_sc_hd__conb_1 _38477_ (.LO(trace_data[2]));
 sky130_fd_sc_hd__conb_1 _38478_ (.LO(trace_data[3]));
 sky130_fd_sc_hd__conb_1 _38479_ (.LO(trace_data[4]));
 sky130_fd_sc_hd__conb_1 _38480_ (.LO(trace_data[5]));
 sky130_fd_sc_hd__conb_1 _38481_ (.LO(trace_data[6]));
 sky130_fd_sc_hd__conb_1 _38482_ (.LO(trace_data[7]));
 sky130_fd_sc_hd__conb_1 _38483_ (.LO(trace_data[8]));
 sky130_fd_sc_hd__conb_1 _38484_ (.LO(trace_data[9]));
 sky130_fd_sc_hd__conb_1 _38485_ (.LO(trace_data[10]));
 sky130_fd_sc_hd__conb_1 _38486_ (.LO(trace_data[11]));
 sky130_fd_sc_hd__conb_1 _38487_ (.LO(trace_data[12]));
 sky130_fd_sc_hd__conb_1 _38488_ (.LO(trace_data[13]));
 sky130_fd_sc_hd__conb_1 _38489_ (.LO(trace_data[14]));
 sky130_fd_sc_hd__conb_1 _38490_ (.LO(trace_data[15]));
 sky130_fd_sc_hd__conb_1 _38491_ (.LO(trace_data[16]));
 sky130_fd_sc_hd__conb_1 _38492_ (.LO(trace_data[17]));
 sky130_fd_sc_hd__conb_1 _38493_ (.LO(trace_data[18]));
 sky130_fd_sc_hd__conb_1 _38494_ (.LO(trace_data[19]));
 sky130_fd_sc_hd__conb_1 _38495_ (.LO(trace_data[20]));
 sky130_fd_sc_hd__conb_1 _38496_ (.LO(trace_data[21]));
 sky130_fd_sc_hd__conb_1 _38497_ (.LO(trace_data[22]));
 sky130_fd_sc_hd__conb_1 _38498_ (.LO(trace_data[23]));
 sky130_fd_sc_hd__conb_1 _38499_ (.LO(trace_data[24]));
 sky130_fd_sc_hd__conb_1 _38500_ (.LO(trace_data[25]));
 sky130_fd_sc_hd__conb_1 _38501_ (.LO(trace_data[26]));
 sky130_fd_sc_hd__conb_1 _38502_ (.LO(trace_data[27]));
 sky130_fd_sc_hd__conb_1 _38503_ (.LO(trace_data[28]));
 sky130_fd_sc_hd__conb_1 _38504_ (.LO(trace_data[29]));
 sky130_fd_sc_hd__conb_1 _38505_ (.LO(trace_data[30]));
 sky130_fd_sc_hd__conb_1 _38506_ (.LO(trace_data[31]));
 sky130_fd_sc_hd__conb_1 _38507_ (.LO(trace_data[32]));
 sky130_fd_sc_hd__conb_1 _38508_ (.LO(trace_data[33]));
 sky130_fd_sc_hd__conb_1 _38509_ (.LO(trace_data[34]));
 sky130_fd_sc_hd__conb_1 _38510_ (.LO(trace_data[35]));
 sky130_fd_sc_hd__conb_1 _38511_ (.LO(trace_valid));
 sky130_fd_sc_hd__conb_1 _38512_ (.LO(_00313_));
 sky130_fd_sc_hd__buf_2 _38513_ (.A(mem_la_wdata[0]),
    .X(pcpi_rs2[0]));
 sky130_fd_sc_hd__buf_2 _38514_ (.A(mem_la_wdata[1]),
    .X(pcpi_rs2[1]));
 sky130_fd_sc_hd__buf_2 _38515_ (.A(mem_la_wdata[2]),
    .X(pcpi_rs2[2]));
 sky130_fd_sc_hd__buf_2 _38516_ (.A(mem_la_wdata[3]),
    .X(pcpi_rs2[3]));
 sky130_fd_sc_hd__buf_2 _38517_ (.A(mem_la_wdata[4]),
    .X(pcpi_rs2[4]));
 sky130_fd_sc_hd__buf_2 _38518_ (.A(mem_la_wdata[5]),
    .X(pcpi_rs2[5]));
 sky130_fd_sc_hd__buf_2 _38519_ (.A(mem_la_wdata[6]),
    .X(pcpi_rs2[6]));
 sky130_fd_sc_hd__buf_2 _38520_ (.A(mem_la_wdata[7]),
    .X(pcpi_rs2[7]));
 sky130_fd_sc_hd__mux2_1 _38521_ (.A0(decoder_trigger),
    .A1(_02410_),
    .S(_00309_),
    .X(_19782_));
 sky130_fd_sc_hd__mux2_1 _38522_ (.A0(\reg_out[2] ),
    .A1(\reg_next_pc[2] ),
    .S(_02183_),
    .X(_02184_));
 sky130_fd_sc_hd__mux2_1 _38523_ (.A0(_02184_),
    .A1(pcpi_rs1[2]),
    .S(_00301_),
    .X(mem_la_addr[2]));
 sky130_fd_sc_hd__mux2_1 _38524_ (.A0(\reg_out[3] ),
    .A1(\reg_next_pc[3] ),
    .S(_02183_),
    .X(_02185_));
 sky130_fd_sc_hd__mux2_1 _38525_ (.A0(_02185_),
    .A1(pcpi_rs1[3]),
    .S(_00301_),
    .X(mem_la_addr[3]));
 sky130_fd_sc_hd__mux2_1 _38526_ (.A0(\reg_out[4] ),
    .A1(\reg_next_pc[4] ),
    .S(_02183_),
    .X(_02186_));
 sky130_fd_sc_hd__mux2_1 _38527_ (.A0(_02186_),
    .A1(pcpi_rs1[4]),
    .S(_00301_),
    .X(mem_la_addr[4]));
 sky130_fd_sc_hd__mux2_1 _38528_ (.A0(\reg_out[5] ),
    .A1(\reg_next_pc[5] ),
    .S(_02183_),
    .X(_02187_));
 sky130_fd_sc_hd__mux2_1 _38529_ (.A0(_02187_),
    .A1(pcpi_rs1[5]),
    .S(_00301_),
    .X(mem_la_addr[5]));
 sky130_fd_sc_hd__mux2_1 _38530_ (.A0(\reg_out[6] ),
    .A1(\reg_next_pc[6] ),
    .S(_02183_),
    .X(_02188_));
 sky130_fd_sc_hd__mux2_1 _38531_ (.A0(_02188_),
    .A1(pcpi_rs1[6]),
    .S(_00301_),
    .X(mem_la_addr[6]));
 sky130_fd_sc_hd__mux2_1 _38532_ (.A0(\reg_out[7] ),
    .A1(\reg_next_pc[7] ),
    .S(_02183_),
    .X(_02189_));
 sky130_fd_sc_hd__mux2_1 _38533_ (.A0(_02189_),
    .A1(pcpi_rs1[7]),
    .S(_00301_),
    .X(mem_la_addr[7]));
 sky130_fd_sc_hd__mux2_1 _38534_ (.A0(\reg_out[8] ),
    .A1(\reg_next_pc[8] ),
    .S(_02183_),
    .X(_02190_));
 sky130_fd_sc_hd__mux2_1 _38535_ (.A0(_02190_),
    .A1(pcpi_rs1[8]),
    .S(_00301_),
    .X(mem_la_addr[8]));
 sky130_fd_sc_hd__mux2_1 _38536_ (.A0(\reg_out[9] ),
    .A1(\reg_next_pc[9] ),
    .S(_02183_),
    .X(_02191_));
 sky130_fd_sc_hd__mux2_1 _38537_ (.A0(_02191_),
    .A1(pcpi_rs1[9]),
    .S(_00301_),
    .X(mem_la_addr[9]));
 sky130_fd_sc_hd__mux2_1 _38538_ (.A0(\reg_out[10] ),
    .A1(\reg_next_pc[10] ),
    .S(_02183_),
    .X(_02192_));
 sky130_fd_sc_hd__mux2_1 _38539_ (.A0(_02192_),
    .A1(pcpi_rs1[10]),
    .S(_00301_),
    .X(mem_la_addr[10]));
 sky130_fd_sc_hd__mux2_1 _38540_ (.A0(\reg_out[11] ),
    .A1(\reg_next_pc[11] ),
    .S(_02183_),
    .X(_02193_));
 sky130_fd_sc_hd__mux2_1 _38541_ (.A0(_02193_),
    .A1(pcpi_rs1[11]),
    .S(_00301_),
    .X(mem_la_addr[11]));
 sky130_fd_sc_hd__mux2_1 _38542_ (.A0(\reg_out[12] ),
    .A1(\reg_next_pc[12] ),
    .S(_02183_),
    .X(_02194_));
 sky130_fd_sc_hd__mux2_1 _38543_ (.A0(_02194_),
    .A1(pcpi_rs1[12]),
    .S(_00301_),
    .X(mem_la_addr[12]));
 sky130_fd_sc_hd__mux2_1 _38544_ (.A0(\reg_out[13] ),
    .A1(\reg_next_pc[13] ),
    .S(_02183_),
    .X(_02195_));
 sky130_fd_sc_hd__mux2_1 _38545_ (.A0(_02195_),
    .A1(pcpi_rs1[13]),
    .S(_00301_),
    .X(mem_la_addr[13]));
 sky130_fd_sc_hd__mux2_1 _38546_ (.A0(\reg_out[14] ),
    .A1(\reg_next_pc[14] ),
    .S(_02183_),
    .X(_02196_));
 sky130_fd_sc_hd__mux2_1 _38547_ (.A0(_02196_),
    .A1(pcpi_rs1[14]),
    .S(_00301_),
    .X(mem_la_addr[14]));
 sky130_fd_sc_hd__mux2_1 _38548_ (.A0(\reg_out[15] ),
    .A1(\reg_next_pc[15] ),
    .S(_02183_),
    .X(_02197_));
 sky130_fd_sc_hd__mux2_1 _38549_ (.A0(_02197_),
    .A1(pcpi_rs1[15]),
    .S(_00301_),
    .X(mem_la_addr[15]));
 sky130_fd_sc_hd__mux2_1 _38550_ (.A0(\reg_out[16] ),
    .A1(\reg_next_pc[16] ),
    .S(_02183_),
    .X(_02198_));
 sky130_fd_sc_hd__mux2_1 _38551_ (.A0(_02198_),
    .A1(pcpi_rs1[16]),
    .S(_00301_),
    .X(mem_la_addr[16]));
 sky130_fd_sc_hd__mux2_1 _38552_ (.A0(\reg_out[17] ),
    .A1(\reg_next_pc[17] ),
    .S(_02183_),
    .X(_02199_));
 sky130_fd_sc_hd__mux2_1 _38553_ (.A0(_02199_),
    .A1(pcpi_rs1[17]),
    .S(_00301_),
    .X(mem_la_addr[17]));
 sky130_fd_sc_hd__mux2_1 _38554_ (.A0(\reg_out[18] ),
    .A1(\reg_next_pc[18] ),
    .S(_02183_),
    .X(_02200_));
 sky130_fd_sc_hd__mux2_1 _38555_ (.A0(_02200_),
    .A1(pcpi_rs1[18]),
    .S(_00301_),
    .X(mem_la_addr[18]));
 sky130_fd_sc_hd__mux2_1 _38556_ (.A0(\reg_out[19] ),
    .A1(\reg_next_pc[19] ),
    .S(_02183_),
    .X(_02201_));
 sky130_fd_sc_hd__mux2_1 _38557_ (.A0(_02201_),
    .A1(pcpi_rs1[19]),
    .S(_00301_),
    .X(mem_la_addr[19]));
 sky130_fd_sc_hd__mux2_1 _38558_ (.A0(\reg_out[20] ),
    .A1(\reg_next_pc[20] ),
    .S(_02183_),
    .X(_02202_));
 sky130_fd_sc_hd__mux2_1 _38559_ (.A0(_02202_),
    .A1(pcpi_rs1[20]),
    .S(_00301_),
    .X(mem_la_addr[20]));
 sky130_fd_sc_hd__mux2_1 _38560_ (.A0(\reg_out[21] ),
    .A1(\reg_next_pc[21] ),
    .S(_02183_),
    .X(_02203_));
 sky130_fd_sc_hd__mux2_1 _38561_ (.A0(_02203_),
    .A1(pcpi_rs1[21]),
    .S(_00301_),
    .X(mem_la_addr[21]));
 sky130_fd_sc_hd__mux2_1 _38562_ (.A0(\reg_out[22] ),
    .A1(\reg_next_pc[22] ),
    .S(_02183_),
    .X(_02204_));
 sky130_fd_sc_hd__mux2_1 _38563_ (.A0(_02204_),
    .A1(pcpi_rs1[22]),
    .S(_00301_),
    .X(mem_la_addr[22]));
 sky130_fd_sc_hd__mux2_1 _38564_ (.A0(\reg_out[23] ),
    .A1(\reg_next_pc[23] ),
    .S(_02183_),
    .X(_02205_));
 sky130_fd_sc_hd__mux2_1 _38565_ (.A0(_02205_),
    .A1(pcpi_rs1[23]),
    .S(_00301_),
    .X(mem_la_addr[23]));
 sky130_fd_sc_hd__mux2_1 _38566_ (.A0(\reg_out[24] ),
    .A1(\reg_next_pc[24] ),
    .S(_02183_),
    .X(_02206_));
 sky130_fd_sc_hd__mux2_1 _38567_ (.A0(_02206_),
    .A1(pcpi_rs1[24]),
    .S(_00301_),
    .X(mem_la_addr[24]));
 sky130_fd_sc_hd__mux2_1 _38568_ (.A0(\reg_out[25] ),
    .A1(\reg_next_pc[25] ),
    .S(_02183_),
    .X(_02207_));
 sky130_fd_sc_hd__mux2_1 _38569_ (.A0(_02207_),
    .A1(pcpi_rs1[25]),
    .S(_00301_),
    .X(mem_la_addr[25]));
 sky130_fd_sc_hd__mux2_1 _38570_ (.A0(\reg_out[26] ),
    .A1(\reg_next_pc[26] ),
    .S(_02183_),
    .X(_02208_));
 sky130_fd_sc_hd__mux2_1 _38571_ (.A0(_02208_),
    .A1(pcpi_rs1[26]),
    .S(_00301_),
    .X(mem_la_addr[26]));
 sky130_fd_sc_hd__mux2_1 _38572_ (.A0(\reg_out[27] ),
    .A1(\reg_next_pc[27] ),
    .S(_02183_),
    .X(_02209_));
 sky130_fd_sc_hd__mux2_1 _38573_ (.A0(_02209_),
    .A1(pcpi_rs1[27]),
    .S(_00301_),
    .X(mem_la_addr[27]));
 sky130_fd_sc_hd__mux2_1 _38574_ (.A0(\reg_out[28] ),
    .A1(\reg_next_pc[28] ),
    .S(_02183_),
    .X(_02210_));
 sky130_fd_sc_hd__mux2_1 _38575_ (.A0(_02210_),
    .A1(pcpi_rs1[28]),
    .S(_00301_),
    .X(mem_la_addr[28]));
 sky130_fd_sc_hd__mux2_1 _38576_ (.A0(\reg_out[29] ),
    .A1(\reg_next_pc[29] ),
    .S(_02183_),
    .X(_02211_));
 sky130_fd_sc_hd__mux2_1 _38577_ (.A0(_02211_),
    .A1(pcpi_rs1[29]),
    .S(_00301_),
    .X(mem_la_addr[29]));
 sky130_fd_sc_hd__mux2_1 _38578_ (.A0(\reg_out[30] ),
    .A1(\reg_next_pc[30] ),
    .S(_02183_),
    .X(_02212_));
 sky130_fd_sc_hd__mux2_1 _38579_ (.A0(_02212_),
    .A1(pcpi_rs1[30]),
    .S(_00301_),
    .X(mem_la_addr[30]));
 sky130_fd_sc_hd__mux2_1 _38580_ (.A0(\reg_out[31] ),
    .A1(\reg_next_pc[31] ),
    .S(_02183_),
    .X(_02213_));
 sky130_fd_sc_hd__mux2_1 _38581_ (.A0(_02213_),
    .A1(pcpi_rs1[31]),
    .S(_00301_),
    .X(mem_la_addr[31]));
 sky130_fd_sc_hd__mux2_1 _38582_ (.A0(_02167_),
    .A1(pcpi_rs2[8]),
    .S(_01683_),
    .X(mem_la_wdata[8]));
 sky130_fd_sc_hd__mux2_1 _38583_ (.A0(_02168_),
    .A1(pcpi_rs2[9]),
    .S(_01683_),
    .X(mem_la_wdata[9]));
 sky130_fd_sc_hd__mux2_1 _38584_ (.A0(_02169_),
    .A1(pcpi_rs2[10]),
    .S(_01683_),
    .X(mem_la_wdata[10]));
 sky130_fd_sc_hd__mux2_1 _38585_ (.A0(_02170_),
    .A1(pcpi_rs2[11]),
    .S(_01683_),
    .X(mem_la_wdata[11]));
 sky130_fd_sc_hd__mux2_1 _38586_ (.A0(_02171_),
    .A1(pcpi_rs2[12]),
    .S(_01683_),
    .X(mem_la_wdata[12]));
 sky130_fd_sc_hd__mux2_1 _38587_ (.A0(_02172_),
    .A1(pcpi_rs2[13]),
    .S(_01683_),
    .X(mem_la_wdata[13]));
 sky130_fd_sc_hd__mux2_1 _38588_ (.A0(_02173_),
    .A1(pcpi_rs2[14]),
    .S(_01683_),
    .X(mem_la_wdata[14]));
 sky130_fd_sc_hd__mux2_1 _38589_ (.A0(_02174_),
    .A1(pcpi_rs2[15]),
    .S(_01683_),
    .X(mem_la_wdata[15]));
 sky130_fd_sc_hd__mux2_1 _38590_ (.A0(_02175_),
    .A1(pcpi_rs2[16]),
    .S(_01683_),
    .X(mem_la_wdata[16]));
 sky130_fd_sc_hd__mux2_1 _38591_ (.A0(_02176_),
    .A1(pcpi_rs2[17]),
    .S(_01683_),
    .X(mem_la_wdata[17]));
 sky130_fd_sc_hd__mux2_1 _38592_ (.A0(_02177_),
    .A1(pcpi_rs2[18]),
    .S(_01683_),
    .X(mem_la_wdata[18]));
 sky130_fd_sc_hd__mux2_1 _38593_ (.A0(_02178_),
    .A1(pcpi_rs2[19]),
    .S(_01683_),
    .X(mem_la_wdata[19]));
 sky130_fd_sc_hd__mux2_1 _38594_ (.A0(_02179_),
    .A1(pcpi_rs2[20]),
    .S(_01683_),
    .X(mem_la_wdata[20]));
 sky130_fd_sc_hd__mux2_1 _38595_ (.A0(_02180_),
    .A1(pcpi_rs2[21]),
    .S(_01683_),
    .X(mem_la_wdata[21]));
 sky130_fd_sc_hd__mux2_1 _38596_ (.A0(_02181_),
    .A1(pcpi_rs2[22]),
    .S(_01683_),
    .X(mem_la_wdata[22]));
 sky130_fd_sc_hd__mux2_1 _38597_ (.A0(_02182_),
    .A1(pcpi_rs2[23]),
    .S(_01683_),
    .X(mem_la_wdata[23]));
 sky130_fd_sc_hd__mux2_1 _38598_ (.A0(_02167_),
    .A1(pcpi_rs2[24]),
    .S(_01683_),
    .X(mem_la_wdata[24]));
 sky130_fd_sc_hd__mux2_1 _38599_ (.A0(_02168_),
    .A1(pcpi_rs2[25]),
    .S(_01683_),
    .X(mem_la_wdata[25]));
 sky130_fd_sc_hd__mux2_1 _38600_ (.A0(_02169_),
    .A1(pcpi_rs2[26]),
    .S(_01683_),
    .X(mem_la_wdata[26]));
 sky130_fd_sc_hd__mux2_1 _38601_ (.A0(_02170_),
    .A1(pcpi_rs2[27]),
    .S(_01683_),
    .X(mem_la_wdata[27]));
 sky130_fd_sc_hd__mux2_1 _38602_ (.A0(_02171_),
    .A1(pcpi_rs2[28]),
    .S(_01683_),
    .X(mem_la_wdata[28]));
 sky130_fd_sc_hd__mux2_1 _38603_ (.A0(_02172_),
    .A1(pcpi_rs2[29]),
    .S(_01683_),
    .X(mem_la_wdata[29]));
 sky130_fd_sc_hd__mux2_1 _38604_ (.A0(_02173_),
    .A1(pcpi_rs2[30]),
    .S(_01683_),
    .X(mem_la_wdata[30]));
 sky130_fd_sc_hd__mux2_1 _38605_ (.A0(_02174_),
    .A1(pcpi_rs2[31]),
    .S(_01683_),
    .X(mem_la_wdata[31]));
 sky130_fd_sc_hd__mux2_1 _38606_ (.A0(\mem_rdata_q[7] ),
    .A1(mem_rdata[7]),
    .S(mem_xfer),
    .X(\mem_rdata_latched[7] ));
 sky130_fd_sc_hd__mux2_1 _38607_ (.A0(\mem_rdata_q[8] ),
    .A1(mem_rdata[8]),
    .S(mem_xfer),
    .X(\mem_rdata_latched[8] ));
 sky130_fd_sc_hd__mux2_1 _38608_ (.A0(\mem_rdata_q[9] ),
    .A1(mem_rdata[9]),
    .S(mem_xfer),
    .X(\mem_rdata_latched[9] ));
 sky130_fd_sc_hd__mux2_1 _38609_ (.A0(\mem_rdata_q[10] ),
    .A1(mem_rdata[10]),
    .S(mem_xfer),
    .X(\mem_rdata_latched[10] ));
 sky130_fd_sc_hd__mux2_1 _38610_ (.A0(\mem_rdata_q[11] ),
    .A1(mem_rdata[11]),
    .S(mem_xfer),
    .X(\mem_rdata_latched[11] ));
 sky130_fd_sc_hd__mux2_1 _38611_ (.A0(\mem_rdata_q[12] ),
    .A1(mem_rdata[12]),
    .S(mem_xfer),
    .X(\mem_rdata_latched[12] ));
 sky130_fd_sc_hd__mux2_1 _38612_ (.A0(\mem_rdata_q[13] ),
    .A1(mem_rdata[13]),
    .S(mem_xfer),
    .X(\mem_rdata_latched[13] ));
 sky130_fd_sc_hd__mux2_1 _38613_ (.A0(\mem_rdata_q[14] ),
    .A1(mem_rdata[14]),
    .S(mem_xfer),
    .X(\mem_rdata_latched[14] ));
 sky130_fd_sc_hd__mux2_1 _38614_ (.A0(\mem_rdata_q[15] ),
    .A1(mem_rdata[15]),
    .S(mem_xfer),
    .X(\mem_rdata_latched[15] ));
 sky130_fd_sc_hd__mux2_1 _38615_ (.A0(\mem_rdata_q[16] ),
    .A1(mem_rdata[16]),
    .S(mem_xfer),
    .X(\mem_rdata_latched[16] ));
 sky130_fd_sc_hd__mux2_1 _38616_ (.A0(\mem_rdata_q[17] ),
    .A1(mem_rdata[17]),
    .S(mem_xfer),
    .X(\mem_rdata_latched[17] ));
 sky130_fd_sc_hd__mux2_1 _38617_ (.A0(\mem_rdata_q[18] ),
    .A1(mem_rdata[18]),
    .S(mem_xfer),
    .X(\mem_rdata_latched[18] ));
 sky130_fd_sc_hd__mux2_1 _38618_ (.A0(\mem_rdata_q[19] ),
    .A1(mem_rdata[19]),
    .S(mem_xfer),
    .X(\mem_rdata_latched[19] ));
 sky130_fd_sc_hd__mux2_1 _38619_ (.A0(\mem_rdata_q[20] ),
    .A1(mem_rdata[20]),
    .S(mem_xfer),
    .X(\mem_rdata_latched[20] ));
 sky130_fd_sc_hd__mux2_1 _38620_ (.A0(\mem_rdata_q[21] ),
    .A1(mem_rdata[21]),
    .S(mem_xfer),
    .X(\mem_rdata_latched[21] ));
 sky130_fd_sc_hd__mux2_1 _38621_ (.A0(\mem_rdata_q[22] ),
    .A1(mem_rdata[22]),
    .S(mem_xfer),
    .X(\mem_rdata_latched[22] ));
 sky130_fd_sc_hd__mux2_1 _38622_ (.A0(\mem_rdata_q[23] ),
    .A1(mem_rdata[23]),
    .S(mem_xfer),
    .X(\mem_rdata_latched[23] ));
 sky130_fd_sc_hd__mux2_1 _38623_ (.A0(\mem_rdata_q[24] ),
    .A1(mem_rdata[24]),
    .S(mem_xfer),
    .X(\mem_rdata_latched[24] ));
 sky130_fd_sc_hd__mux2_1 _38624_ (.A0(\mem_rdata_q[25] ),
    .A1(mem_rdata[25]),
    .S(mem_xfer),
    .X(\mem_rdata_latched[25] ));
 sky130_fd_sc_hd__mux2_1 _38625_ (.A0(\mem_rdata_q[26] ),
    .A1(mem_rdata[26]),
    .S(mem_xfer),
    .X(\mem_rdata_latched[26] ));
 sky130_fd_sc_hd__mux2_1 _38626_ (.A0(\mem_rdata_q[27] ),
    .A1(mem_rdata[27]),
    .S(mem_xfer),
    .X(\mem_rdata_latched[27] ));
 sky130_fd_sc_hd__mux2_1 _38627_ (.A0(\mem_rdata_q[28] ),
    .A1(mem_rdata[28]),
    .S(mem_xfer),
    .X(\mem_rdata_latched[28] ));
 sky130_fd_sc_hd__mux2_1 _38628_ (.A0(\mem_rdata_q[29] ),
    .A1(mem_rdata[29]),
    .S(mem_xfer),
    .X(\mem_rdata_latched[29] ));
 sky130_fd_sc_hd__mux2_1 _38629_ (.A0(\mem_rdata_q[30] ),
    .A1(mem_rdata[30]),
    .S(mem_xfer),
    .X(\mem_rdata_latched[30] ));
 sky130_fd_sc_hd__mux2_1 _38630_ (.A0(\mem_rdata_q[31] ),
    .A1(mem_rdata[31]),
    .S(mem_xfer),
    .X(\mem_rdata_latched[31] ));
 sky130_fd_sc_hd__mux2_1 _38631_ (.A0(_02134_),
    .A1(\alu_add_sub[0] ),
    .S(_02133_),
    .X(\alu_out[0] ));
 sky130_fd_sc_hd__mux2_1 _38632_ (.A0(_02135_),
    .A1(\alu_add_sub[1] ),
    .S(_02133_),
    .X(\alu_out[1] ));
 sky130_fd_sc_hd__mux2_1 _38633_ (.A0(_02136_),
    .A1(\alu_add_sub[2] ),
    .S(_02133_),
    .X(\alu_out[2] ));
 sky130_fd_sc_hd__mux2_1 _38634_ (.A0(_02137_),
    .A1(\alu_add_sub[3] ),
    .S(_02133_),
    .X(\alu_out[3] ));
 sky130_fd_sc_hd__mux2_1 _38635_ (.A0(_02138_),
    .A1(\alu_add_sub[4] ),
    .S(_02133_),
    .X(\alu_out[4] ));
 sky130_fd_sc_hd__mux2_1 _38636_ (.A0(_02139_),
    .A1(\alu_add_sub[5] ),
    .S(_02133_),
    .X(\alu_out[5] ));
 sky130_fd_sc_hd__mux2_1 _38637_ (.A0(_02140_),
    .A1(\alu_add_sub[6] ),
    .S(_02133_),
    .X(\alu_out[6] ));
 sky130_fd_sc_hd__mux2_1 _38638_ (.A0(_02141_),
    .A1(\alu_add_sub[7] ),
    .S(_02133_),
    .X(\alu_out[7] ));
 sky130_fd_sc_hd__mux2_1 _38639_ (.A0(_02142_),
    .A1(\alu_add_sub[8] ),
    .S(_02133_),
    .X(\alu_out[8] ));
 sky130_fd_sc_hd__mux2_1 _38640_ (.A0(_02143_),
    .A1(\alu_add_sub[9] ),
    .S(_02133_),
    .X(\alu_out[9] ));
 sky130_fd_sc_hd__mux2_1 _38641_ (.A0(_02144_),
    .A1(\alu_add_sub[10] ),
    .S(_02133_),
    .X(\alu_out[10] ));
 sky130_fd_sc_hd__mux2_1 _38642_ (.A0(_02145_),
    .A1(\alu_add_sub[11] ),
    .S(_02133_),
    .X(\alu_out[11] ));
 sky130_fd_sc_hd__mux2_1 _38643_ (.A0(_02146_),
    .A1(\alu_add_sub[12] ),
    .S(_02133_),
    .X(\alu_out[12] ));
 sky130_fd_sc_hd__mux2_1 _38644_ (.A0(_02147_),
    .A1(\alu_add_sub[13] ),
    .S(_02133_),
    .X(\alu_out[13] ));
 sky130_fd_sc_hd__mux2_1 _38645_ (.A0(_02148_),
    .A1(\alu_add_sub[14] ),
    .S(_02133_),
    .X(\alu_out[14] ));
 sky130_fd_sc_hd__mux2_1 _38646_ (.A0(_02149_),
    .A1(\alu_add_sub[15] ),
    .S(_02133_),
    .X(\alu_out[15] ));
 sky130_fd_sc_hd__mux2_1 _38647_ (.A0(_02150_),
    .A1(\alu_add_sub[16] ),
    .S(_02133_),
    .X(\alu_out[16] ));
 sky130_fd_sc_hd__mux2_1 _38648_ (.A0(_02151_),
    .A1(\alu_add_sub[17] ),
    .S(_02133_),
    .X(\alu_out[17] ));
 sky130_fd_sc_hd__mux2_1 _38649_ (.A0(_02152_),
    .A1(\alu_add_sub[18] ),
    .S(_02133_),
    .X(\alu_out[18] ));
 sky130_fd_sc_hd__mux2_1 _38650_ (.A0(_02153_),
    .A1(\alu_add_sub[19] ),
    .S(_02133_),
    .X(\alu_out[19] ));
 sky130_fd_sc_hd__mux2_1 _38651_ (.A0(_02154_),
    .A1(\alu_add_sub[20] ),
    .S(_02133_),
    .X(\alu_out[20] ));
 sky130_fd_sc_hd__mux2_1 _38652_ (.A0(_02155_),
    .A1(\alu_add_sub[21] ),
    .S(_02133_),
    .X(\alu_out[21] ));
 sky130_fd_sc_hd__mux2_1 _38653_ (.A0(_02156_),
    .A1(\alu_add_sub[22] ),
    .S(_02133_),
    .X(\alu_out[22] ));
 sky130_fd_sc_hd__mux2_1 _38654_ (.A0(_02157_),
    .A1(\alu_add_sub[23] ),
    .S(_02133_),
    .X(\alu_out[23] ));
 sky130_fd_sc_hd__mux2_1 _38655_ (.A0(_02158_),
    .A1(\alu_add_sub[24] ),
    .S(_02133_),
    .X(\alu_out[24] ));
 sky130_fd_sc_hd__mux2_1 _38656_ (.A0(_02159_),
    .A1(\alu_add_sub[25] ),
    .S(_02133_),
    .X(\alu_out[25] ));
 sky130_fd_sc_hd__mux2_1 _38657_ (.A0(_02160_),
    .A1(\alu_add_sub[26] ),
    .S(_02133_),
    .X(\alu_out[26] ));
 sky130_fd_sc_hd__mux2_1 _38658_ (.A0(_02161_),
    .A1(\alu_add_sub[27] ),
    .S(_02133_),
    .X(\alu_out[27] ));
 sky130_fd_sc_hd__mux2_1 _38659_ (.A0(_02162_),
    .A1(\alu_add_sub[28] ),
    .S(_02133_),
    .X(\alu_out[28] ));
 sky130_fd_sc_hd__mux2_1 _38660_ (.A0(_02163_),
    .A1(\alu_add_sub[29] ),
    .S(_02133_),
    .X(\alu_out[29] ));
 sky130_fd_sc_hd__mux2_1 _38661_ (.A0(_02164_),
    .A1(\alu_add_sub[30] ),
    .S(_02133_),
    .X(\alu_out[30] ));
 sky130_fd_sc_hd__mux2_1 _38662_ (.A0(_02165_),
    .A1(\alu_add_sub[31] ),
    .S(_02133_),
    .X(\alu_out[31] ));
 sky130_fd_sc_hd__mux2_1 _38663_ (.A0(_02071_),
    .A1(\reg_next_pc[0] ),
    .S(_02069_),
    .X(\cpuregs_wrdata[0] ));
 sky130_fd_sc_hd__mux2_1 _38664_ (.A0(_02072_),
    .A1(\reg_pc[1] ),
    .S(_02069_),
    .X(\cpuregs_wrdata[1] ));
 sky130_fd_sc_hd__mux2_1 _38665_ (.A0(_02074_),
    .A1(_02073_),
    .S(_02069_),
    .X(\cpuregs_wrdata[2] ));
 sky130_fd_sc_hd__mux2_1 _38666_ (.A0(_02076_),
    .A1(_02075_),
    .S(_02069_),
    .X(\cpuregs_wrdata[3] ));
 sky130_fd_sc_hd__mux2_1 _38667_ (.A0(_02078_),
    .A1(_02077_),
    .S(_02069_),
    .X(\cpuregs_wrdata[4] ));
 sky130_fd_sc_hd__mux2_1 _38668_ (.A0(_02080_),
    .A1(_02079_),
    .S(_02069_),
    .X(\cpuregs_wrdata[5] ));
 sky130_fd_sc_hd__mux2_1 _38669_ (.A0(_02082_),
    .A1(_02081_),
    .S(_02069_),
    .X(\cpuregs_wrdata[6] ));
 sky130_fd_sc_hd__mux2_1 _38670_ (.A0(_02084_),
    .A1(_02083_),
    .S(_02069_),
    .X(\cpuregs_wrdata[7] ));
 sky130_fd_sc_hd__mux2_1 _38671_ (.A0(_02086_),
    .A1(_02085_),
    .S(_02069_),
    .X(\cpuregs_wrdata[8] ));
 sky130_fd_sc_hd__mux2_1 _38672_ (.A0(_02088_),
    .A1(_02087_),
    .S(_02069_),
    .X(\cpuregs_wrdata[9] ));
 sky130_fd_sc_hd__mux2_1 _38673_ (.A0(_02090_),
    .A1(_02089_),
    .S(_02069_),
    .X(\cpuregs_wrdata[10] ));
 sky130_fd_sc_hd__mux2_1 _38674_ (.A0(_02092_),
    .A1(_02091_),
    .S(_02069_),
    .X(\cpuregs_wrdata[11] ));
 sky130_fd_sc_hd__mux2_1 _38675_ (.A0(_02094_),
    .A1(_02093_),
    .S(_02069_),
    .X(\cpuregs_wrdata[12] ));
 sky130_fd_sc_hd__mux2_1 _38676_ (.A0(_02096_),
    .A1(_02095_),
    .S(_02069_),
    .X(\cpuregs_wrdata[13] ));
 sky130_fd_sc_hd__mux2_1 _38677_ (.A0(_02098_),
    .A1(_02097_),
    .S(_02069_),
    .X(\cpuregs_wrdata[14] ));
 sky130_fd_sc_hd__mux2_1 _38678_ (.A0(_02100_),
    .A1(_02099_),
    .S(_02069_),
    .X(\cpuregs_wrdata[15] ));
 sky130_fd_sc_hd__mux2_1 _38679_ (.A0(_02102_),
    .A1(_02101_),
    .S(_02069_),
    .X(\cpuregs_wrdata[16] ));
 sky130_fd_sc_hd__mux2_1 _38680_ (.A0(_02104_),
    .A1(_02103_),
    .S(_02069_),
    .X(\cpuregs_wrdata[17] ));
 sky130_fd_sc_hd__mux2_1 _38681_ (.A0(_02106_),
    .A1(_02105_),
    .S(_02069_),
    .X(\cpuregs_wrdata[18] ));
 sky130_fd_sc_hd__mux2_1 _38682_ (.A0(_02108_),
    .A1(_02107_),
    .S(_02069_),
    .X(\cpuregs_wrdata[19] ));
 sky130_fd_sc_hd__mux2_1 _38683_ (.A0(_02110_),
    .A1(_02109_),
    .S(_02069_),
    .X(\cpuregs_wrdata[20] ));
 sky130_fd_sc_hd__mux2_1 _38684_ (.A0(_02112_),
    .A1(_02111_),
    .S(_02069_),
    .X(\cpuregs_wrdata[21] ));
 sky130_fd_sc_hd__mux2_1 _38685_ (.A0(_02114_),
    .A1(_02113_),
    .S(_02069_),
    .X(\cpuregs_wrdata[22] ));
 sky130_fd_sc_hd__mux2_1 _38686_ (.A0(_02116_),
    .A1(_02115_),
    .S(_02069_),
    .X(\cpuregs_wrdata[23] ));
 sky130_fd_sc_hd__mux2_1 _38687_ (.A0(_02118_),
    .A1(_02117_),
    .S(_02069_),
    .X(\cpuregs_wrdata[24] ));
 sky130_fd_sc_hd__mux2_1 _38688_ (.A0(_02120_),
    .A1(_02119_),
    .S(_02069_),
    .X(\cpuregs_wrdata[25] ));
 sky130_fd_sc_hd__mux2_1 _38689_ (.A0(_02122_),
    .A1(_02121_),
    .S(_02069_),
    .X(\cpuregs_wrdata[26] ));
 sky130_fd_sc_hd__mux2_1 _38690_ (.A0(_02124_),
    .A1(_02123_),
    .S(_02069_),
    .X(\cpuregs_wrdata[27] ));
 sky130_fd_sc_hd__mux2_1 _38691_ (.A0(_02126_),
    .A1(_02125_),
    .S(_02069_),
    .X(\cpuregs_wrdata[28] ));
 sky130_fd_sc_hd__mux2_1 _38692_ (.A0(_02128_),
    .A1(_02127_),
    .S(_02069_),
    .X(\cpuregs_wrdata[29] ));
 sky130_fd_sc_hd__mux2_1 _38693_ (.A0(_02130_),
    .A1(_02129_),
    .S(_02069_),
    .X(\cpuregs_wrdata[30] ));
 sky130_fd_sc_hd__mux2_1 _38694_ (.A0(_02132_),
    .A1(_02131_),
    .S(_02069_),
    .X(\cpuregs_wrdata[31] ));
 sky130_fd_sc_hd__mux2_1 _38695_ (.A0(_02316_),
    .A1(_02317_),
    .S(_00307_),
    .X(_00004_));
 sky130_fd_sc_hd__mux2_1 _38696_ (.A0(_00347_),
    .A1(_19783_),
    .S(_00336_),
    .X(_00348_));
 sky130_fd_sc_hd__mux2_1 _38697_ (.A0(_19783_),
    .A1(_00348_),
    .S(resetn),
    .X(_00003_));
 sky130_fd_sc_hd__mux2_1 _38698_ (.A0(_02304_),
    .A1(_02305_),
    .S(\irq_state[1] ),
    .X(_02306_));
 sky130_fd_sc_hd__mux2_1 _38699_ (.A0(_02306_),
    .A1(_02304_),
    .S(_02217_),
    .X(_00008_));
 sky130_fd_sc_hd__mux2_1 _38700_ (.A0(_02214_),
    .A1(_02215_),
    .S(\irq_state[1] ),
    .X(_02216_));
 sky130_fd_sc_hd__mux2_1 _38701_ (.A0(_02216_),
    .A1(_02214_),
    .S(_02217_),
    .X(_00031_));
 sky130_fd_sc_hd__mux2_1 _38702_ (.A0(_02218_),
    .A1(_02219_),
    .S(\irq_state[1] ),
    .X(_02220_));
 sky130_fd_sc_hd__mux2_1 _38703_ (.A0(_02220_),
    .A1(_02218_),
    .S(_02217_),
    .X(_00032_));
 sky130_fd_sc_hd__mux2_1 _38704_ (.A0(_02221_),
    .A1(_02222_),
    .S(\irq_state[1] ),
    .X(_02223_));
 sky130_fd_sc_hd__mux2_1 _38705_ (.A0(_02223_),
    .A1(_02221_),
    .S(_02217_),
    .X(_00033_));
 sky130_fd_sc_hd__mux2_1 _38706_ (.A0(_02224_),
    .A1(_02225_),
    .S(\irq_state[1] ),
    .X(_02226_));
 sky130_fd_sc_hd__mux2_1 _38707_ (.A0(_02226_),
    .A1(_02224_),
    .S(_02217_),
    .X(_00034_));
 sky130_fd_sc_hd__mux2_1 _38708_ (.A0(_02227_),
    .A1(_02228_),
    .S(\irq_state[1] ),
    .X(_02229_));
 sky130_fd_sc_hd__mux2_1 _38709_ (.A0(_02229_),
    .A1(_02227_),
    .S(_02217_),
    .X(_00035_));
 sky130_fd_sc_hd__mux2_1 _38710_ (.A0(_02230_),
    .A1(_02231_),
    .S(\irq_state[1] ),
    .X(_02232_));
 sky130_fd_sc_hd__mux2_1 _38711_ (.A0(_02232_),
    .A1(_02230_),
    .S(_02217_),
    .X(_00036_));
 sky130_fd_sc_hd__mux2_1 _38712_ (.A0(_02233_),
    .A1(_02234_),
    .S(\irq_state[1] ),
    .X(_02235_));
 sky130_fd_sc_hd__mux2_1 _38713_ (.A0(_02235_),
    .A1(_02233_),
    .S(_02217_),
    .X(_00037_));
 sky130_fd_sc_hd__mux2_1 _38714_ (.A0(_02236_),
    .A1(_02237_),
    .S(\irq_state[1] ),
    .X(_02238_));
 sky130_fd_sc_hd__mux2_1 _38715_ (.A0(_02238_),
    .A1(_02236_),
    .S(_02217_),
    .X(_00009_));
 sky130_fd_sc_hd__mux2_1 _38716_ (.A0(_02239_),
    .A1(_02240_),
    .S(\irq_state[1] ),
    .X(_02241_));
 sky130_fd_sc_hd__mux2_1 _38717_ (.A0(_02241_),
    .A1(_02239_),
    .S(_02217_),
    .X(_00010_));
 sky130_fd_sc_hd__mux2_1 _38718_ (.A0(_02242_),
    .A1(_02243_),
    .S(\irq_state[1] ),
    .X(_02244_));
 sky130_fd_sc_hd__mux2_1 _38719_ (.A0(_02244_),
    .A1(_02242_),
    .S(_02217_),
    .X(_00011_));
 sky130_fd_sc_hd__mux2_1 _38720_ (.A0(_02245_),
    .A1(_02246_),
    .S(\irq_state[1] ),
    .X(_02247_));
 sky130_fd_sc_hd__mux2_1 _38721_ (.A0(_02247_),
    .A1(_02245_),
    .S(_02217_),
    .X(_00012_));
 sky130_fd_sc_hd__mux2_1 _38722_ (.A0(_02248_),
    .A1(_02249_),
    .S(\irq_state[1] ),
    .X(_02250_));
 sky130_fd_sc_hd__mux2_1 _38723_ (.A0(_02250_),
    .A1(_02248_),
    .S(_02217_),
    .X(_00013_));
 sky130_fd_sc_hd__mux2_1 _38724_ (.A0(_02251_),
    .A1(_02252_),
    .S(\irq_state[1] ),
    .X(_02253_));
 sky130_fd_sc_hd__mux2_1 _38725_ (.A0(_02253_),
    .A1(_02251_),
    .S(_02217_),
    .X(_00014_));
 sky130_fd_sc_hd__mux2_1 _38726_ (.A0(_02254_),
    .A1(_02255_),
    .S(\irq_state[1] ),
    .X(_02256_));
 sky130_fd_sc_hd__mux2_1 _38727_ (.A0(_02256_),
    .A1(_02254_),
    .S(_02217_),
    .X(_00015_));
 sky130_fd_sc_hd__mux2_1 _38728_ (.A0(_02257_),
    .A1(_02258_),
    .S(\irq_state[1] ),
    .X(_02259_));
 sky130_fd_sc_hd__mux2_1 _38729_ (.A0(_02259_),
    .A1(_02257_),
    .S(_02217_),
    .X(_00016_));
 sky130_fd_sc_hd__mux2_1 _38730_ (.A0(_02260_),
    .A1(_02261_),
    .S(\irq_state[1] ),
    .X(_02262_));
 sky130_fd_sc_hd__mux2_1 _38731_ (.A0(_02262_),
    .A1(_02260_),
    .S(_02217_),
    .X(_00017_));
 sky130_fd_sc_hd__mux2_1 _38732_ (.A0(_02263_),
    .A1(_02264_),
    .S(\irq_state[1] ),
    .X(_02265_));
 sky130_fd_sc_hd__mux2_1 _38733_ (.A0(_02265_),
    .A1(_02263_),
    .S(_02217_),
    .X(_00018_));
 sky130_fd_sc_hd__mux2_1 _38734_ (.A0(_02266_),
    .A1(_02267_),
    .S(\irq_state[1] ),
    .X(_02268_));
 sky130_fd_sc_hd__mux2_1 _38735_ (.A0(_02268_),
    .A1(_02266_),
    .S(_02217_),
    .X(_00019_));
 sky130_fd_sc_hd__mux2_1 _38736_ (.A0(_02269_),
    .A1(_02270_),
    .S(\irq_state[1] ),
    .X(_02271_));
 sky130_fd_sc_hd__mux2_1 _38737_ (.A0(_02271_),
    .A1(_02269_),
    .S(_02217_),
    .X(_00020_));
 sky130_fd_sc_hd__mux2_1 _38738_ (.A0(_02272_),
    .A1(_02273_),
    .S(\irq_state[1] ),
    .X(_02274_));
 sky130_fd_sc_hd__mux2_1 _38739_ (.A0(_02274_),
    .A1(_02272_),
    .S(_02217_),
    .X(_00021_));
 sky130_fd_sc_hd__mux2_1 _38740_ (.A0(_02275_),
    .A1(_02276_),
    .S(\irq_state[1] ),
    .X(_02277_));
 sky130_fd_sc_hd__mux2_1 _38741_ (.A0(_02277_),
    .A1(_02275_),
    .S(_02217_),
    .X(_00022_));
 sky130_fd_sc_hd__mux2_1 _38742_ (.A0(_02278_),
    .A1(_02279_),
    .S(\irq_state[1] ),
    .X(_02280_));
 sky130_fd_sc_hd__mux2_1 _38743_ (.A0(_02280_),
    .A1(_02278_),
    .S(_02217_),
    .X(_00023_));
 sky130_fd_sc_hd__mux2_1 _38744_ (.A0(_02281_),
    .A1(_02282_),
    .S(\irq_state[1] ),
    .X(_02283_));
 sky130_fd_sc_hd__mux2_1 _38745_ (.A0(_02283_),
    .A1(_02281_),
    .S(_02217_),
    .X(_00024_));
 sky130_fd_sc_hd__mux2_1 _38746_ (.A0(_02284_),
    .A1(_02285_),
    .S(\irq_state[1] ),
    .X(_02286_));
 sky130_fd_sc_hd__mux2_1 _38747_ (.A0(_02286_),
    .A1(_02284_),
    .S(_02217_),
    .X(_00025_));
 sky130_fd_sc_hd__mux2_1 _38748_ (.A0(_02287_),
    .A1(_02288_),
    .S(\irq_state[1] ),
    .X(_02289_));
 sky130_fd_sc_hd__mux2_1 _38749_ (.A0(_02289_),
    .A1(_02287_),
    .S(_02217_),
    .X(_00026_));
 sky130_fd_sc_hd__mux2_1 _38750_ (.A0(_02290_),
    .A1(_02291_),
    .S(\irq_state[1] ),
    .X(_02292_));
 sky130_fd_sc_hd__mux2_1 _38751_ (.A0(_02292_),
    .A1(_02290_),
    .S(_02217_),
    .X(_00027_));
 sky130_fd_sc_hd__mux2_1 _38752_ (.A0(_02293_),
    .A1(_02294_),
    .S(\irq_state[1] ),
    .X(_02295_));
 sky130_fd_sc_hd__mux2_1 _38753_ (.A0(_02295_),
    .A1(_02293_),
    .S(_02217_),
    .X(_00028_));
 sky130_fd_sc_hd__mux2_1 _38754_ (.A0(_02296_),
    .A1(_02297_),
    .S(\irq_state[1] ),
    .X(_02298_));
 sky130_fd_sc_hd__mux2_1 _38755_ (.A0(_02298_),
    .A1(_02296_),
    .S(_02217_),
    .X(_00029_));
 sky130_fd_sc_hd__mux2_1 _38756_ (.A0(_02299_),
    .A1(_02300_),
    .S(\irq_state[1] ),
    .X(_02301_));
 sky130_fd_sc_hd__mux2_1 _38757_ (.A0(_02301_),
    .A1(_02299_),
    .S(_02217_),
    .X(_00030_));
 sky130_fd_sc_hd__mux2_1 _38758_ (.A0(_01467_),
    .A1(\reg_next_pc[1] ),
    .S(_00292_),
    .X(_02590_));
 sky130_fd_sc_hd__mux2_1 _38759_ (.A0(_00295_),
    .A1(\reg_next_pc[2] ),
    .S(_00292_),
    .X(_02560_));
 sky130_fd_sc_hd__mux2_1 _38760_ (.A0(_01470_),
    .A1(\reg_next_pc[3] ),
    .S(_00292_),
    .X(_02571_));
 sky130_fd_sc_hd__mux2_1 _38761_ (.A0(_01478_),
    .A1(\reg_next_pc[5] ),
    .S(_00292_),
    .X(_02583_));
 sky130_fd_sc_hd__mux2_1 _38762_ (.A0(_01481_),
    .A1(\reg_next_pc[6] ),
    .S(_00292_),
    .X(_02584_));
 sky130_fd_sc_hd__mux2_1 _38763_ (.A0(_01484_),
    .A1(\reg_next_pc[7] ),
    .S(_00292_),
    .X(_02585_));
 sky130_fd_sc_hd__mux2_1 _38764_ (.A0(_01487_),
    .A1(\reg_next_pc[8] ),
    .S(_00292_),
    .X(_02586_));
 sky130_fd_sc_hd__mux2_1 _38765_ (.A0(_01490_),
    .A1(\reg_next_pc[9] ),
    .S(_00292_),
    .X(_02587_));
 sky130_fd_sc_hd__mux2_1 _38766_ (.A0(_01493_),
    .A1(\reg_next_pc[10] ),
    .S(_00292_),
    .X(_02588_));
 sky130_fd_sc_hd__mux2_1 _38767_ (.A0(_01496_),
    .A1(\reg_next_pc[11] ),
    .S(_00292_),
    .X(_02589_));
 sky130_fd_sc_hd__mux2_1 _38768_ (.A0(_01499_),
    .A1(\reg_next_pc[12] ),
    .S(_00292_),
    .X(_02561_));
 sky130_fd_sc_hd__mux2_1 _38769_ (.A0(_01502_),
    .A1(\reg_next_pc[13] ),
    .S(_00292_),
    .X(_02562_));
 sky130_fd_sc_hd__mux2_1 _38770_ (.A0(_01505_),
    .A1(\reg_next_pc[14] ),
    .S(_00292_),
    .X(_02563_));
 sky130_fd_sc_hd__mux2_1 _38771_ (.A0(_01508_),
    .A1(\reg_next_pc[15] ),
    .S(_00292_),
    .X(_02564_));
 sky130_fd_sc_hd__mux2_1 _38772_ (.A0(_01511_),
    .A1(\reg_next_pc[16] ),
    .S(_00292_),
    .X(_02565_));
 sky130_fd_sc_hd__mux2_1 _38773_ (.A0(_01514_),
    .A1(\reg_next_pc[17] ),
    .S(_00292_),
    .X(_02566_));
 sky130_fd_sc_hd__mux2_1 _38774_ (.A0(_01517_),
    .A1(\reg_next_pc[18] ),
    .S(_00292_),
    .X(_02567_));
 sky130_fd_sc_hd__mux2_1 _38775_ (.A0(_01520_),
    .A1(\reg_next_pc[19] ),
    .S(_00292_),
    .X(_02568_));
 sky130_fd_sc_hd__mux2_1 _38776_ (.A0(_01523_),
    .A1(\reg_next_pc[20] ),
    .S(_00292_),
    .X(_02569_));
 sky130_fd_sc_hd__mux2_1 _38777_ (.A0(_01526_),
    .A1(\reg_next_pc[21] ),
    .S(_00292_),
    .X(_02570_));
 sky130_fd_sc_hd__mux2_1 _38778_ (.A0(_01529_),
    .A1(\reg_next_pc[22] ),
    .S(_00292_),
    .X(_02572_));
 sky130_fd_sc_hd__mux2_1 _38779_ (.A0(_01532_),
    .A1(\reg_next_pc[23] ),
    .S(_00292_),
    .X(_02573_));
 sky130_fd_sc_hd__mux2_1 _38780_ (.A0(_01535_),
    .A1(\reg_next_pc[24] ),
    .S(_00292_),
    .X(_02574_));
 sky130_fd_sc_hd__mux2_1 _38781_ (.A0(_01538_),
    .A1(\reg_next_pc[25] ),
    .S(_00292_),
    .X(_02575_));
 sky130_fd_sc_hd__mux2_1 _38782_ (.A0(_01541_),
    .A1(\reg_next_pc[26] ),
    .S(_00292_),
    .X(_02576_));
 sky130_fd_sc_hd__mux2_1 _38783_ (.A0(_01544_),
    .A1(\reg_next_pc[27] ),
    .S(_00292_),
    .X(_02577_));
 sky130_fd_sc_hd__mux2_1 _38784_ (.A0(_01547_),
    .A1(\reg_next_pc[28] ),
    .S(_00292_),
    .X(_02578_));
 sky130_fd_sc_hd__mux2_1 _38785_ (.A0(_01550_),
    .A1(\reg_next_pc[29] ),
    .S(_00292_),
    .X(_02579_));
 sky130_fd_sc_hd__mux2_1 _38786_ (.A0(_01553_),
    .A1(\reg_next_pc[30] ),
    .S(_00292_),
    .X(_02580_));
 sky130_fd_sc_hd__mux2_1 _38787_ (.A0(_01556_),
    .A1(\reg_next_pc[31] ),
    .S(_00292_),
    .X(_02581_));
 sky130_fd_sc_hd__mux2_1 _38788_ (.A0(_00057_),
    .A1(_00064_),
    .S(mem_la_wdata[3]),
    .X(_00065_));
 sky130_fd_sc_hd__mux2_1 _38789_ (.A0(_00065_),
    .A1(_02543_),
    .S(mem_la_wdata[4]),
    .X(_19819_));
 sky130_fd_sc_hd__mux2_1 _38790_ (.A0(_00075_),
    .A1(_00082_),
    .S(mem_la_wdata[3]),
    .X(_00083_));
 sky130_fd_sc_hd__mux2_1 _38791_ (.A0(_00083_),
    .A1(_02544_),
    .S(mem_la_wdata[4]),
    .X(_19820_));
 sky130_fd_sc_hd__mux2_1 _38792_ (.A0(_00089_),
    .A1(_00092_),
    .S(mem_la_wdata[3]),
    .X(_00093_));
 sky130_fd_sc_hd__mux2_1 _38793_ (.A0(_00093_),
    .A1(_02545_),
    .S(mem_la_wdata[4]),
    .X(_19821_));
 sky130_fd_sc_hd__mux2_1 _38794_ (.A0(_00099_),
    .A1(_00102_),
    .S(mem_la_wdata[3]),
    .X(_00103_));
 sky130_fd_sc_hd__mux2_1 _38795_ (.A0(_00103_),
    .A1(_02546_),
    .S(mem_la_wdata[4]),
    .X(_19822_));
 sky130_fd_sc_hd__mux2_1 _38796_ (.A0(_00107_),
    .A1(_00108_),
    .S(mem_la_wdata[3]),
    .X(_00109_));
 sky130_fd_sc_hd__mux2_1 _38797_ (.A0(_00109_),
    .A1(_02547_),
    .S(mem_la_wdata[4]),
    .X(_19823_));
 sky130_fd_sc_hd__mux2_1 _38798_ (.A0(_00113_),
    .A1(_00114_),
    .S(mem_la_wdata[3]),
    .X(_00115_));
 sky130_fd_sc_hd__mux2_1 _38799_ (.A0(_00115_),
    .A1(_02548_),
    .S(mem_la_wdata[4]),
    .X(_19824_));
 sky130_fd_sc_hd__mux2_1 _38800_ (.A0(_00119_),
    .A1(_00120_),
    .S(mem_la_wdata[3]),
    .X(_00121_));
 sky130_fd_sc_hd__mux2_1 _38801_ (.A0(_00121_),
    .A1(_02549_),
    .S(mem_la_wdata[4]),
    .X(_19825_));
 sky130_fd_sc_hd__mux2_1 _38802_ (.A0(_00125_),
    .A1(_00126_),
    .S(mem_la_wdata[3]),
    .X(_00127_));
 sky130_fd_sc_hd__mux2_1 _38803_ (.A0(_00127_),
    .A1(_02550_),
    .S(mem_la_wdata[4]),
    .X(_19826_));
 sky130_fd_sc_hd__mux2_1 _38804_ (.A0(_00129_),
    .A1(_00106_),
    .S(mem_la_wdata[2]),
    .X(_00130_));
 sky130_fd_sc_hd__mux2_1 _38805_ (.A0(_00130_),
    .A1(_00057_),
    .S(mem_la_wdata[3]),
    .X(_00131_));
 sky130_fd_sc_hd__mux2_1 _38806_ (.A0(_00131_),
    .A1(_02551_),
    .S(mem_la_wdata[4]),
    .X(_19827_));
 sky130_fd_sc_hd__mux2_1 _38807_ (.A0(_00133_),
    .A1(_00112_),
    .S(mem_la_wdata[2]),
    .X(_00134_));
 sky130_fd_sc_hd__mux2_1 _38808_ (.A0(_00134_),
    .A1(_00075_),
    .S(mem_la_wdata[3]),
    .X(_00135_));
 sky130_fd_sc_hd__mux2_1 _38809_ (.A0(_00135_),
    .A1(_02552_),
    .S(mem_la_wdata[4]),
    .X(_19828_));
 sky130_fd_sc_hd__mux2_1 _38810_ (.A0(_00137_),
    .A1(_00118_),
    .S(mem_la_wdata[2]),
    .X(_00138_));
 sky130_fd_sc_hd__mux2_1 _38811_ (.A0(_00138_),
    .A1(_00089_),
    .S(mem_la_wdata[3]),
    .X(_00139_));
 sky130_fd_sc_hd__mux2_1 _38812_ (.A0(_00139_),
    .A1(_02553_),
    .S(mem_la_wdata[4]),
    .X(_19829_));
 sky130_fd_sc_hd__mux2_1 _38813_ (.A0(_00141_),
    .A1(_00124_),
    .S(mem_la_wdata[2]),
    .X(_00142_));
 sky130_fd_sc_hd__mux2_1 _38814_ (.A0(_00142_),
    .A1(_00099_),
    .S(mem_la_wdata[3]),
    .X(_00143_));
 sky130_fd_sc_hd__mux2_1 _38815_ (.A0(_00143_),
    .A1(_02554_),
    .S(mem_la_wdata[4]),
    .X(_19830_));
 sky130_fd_sc_hd__mux2_1 _38816_ (.A0(_00144_),
    .A1(_00136_),
    .S(mem_la_wdata[1]),
    .X(_00145_));
 sky130_fd_sc_hd__mux2_1 _38817_ (.A0(_00145_),
    .A1(_00129_),
    .S(mem_la_wdata[2]),
    .X(_00146_));
 sky130_fd_sc_hd__mux2_1 _38818_ (.A0(_00146_),
    .A1(_00107_),
    .S(mem_la_wdata[3]),
    .X(_00147_));
 sky130_fd_sc_hd__mux2_1 _38819_ (.A0(_00147_),
    .A1(_02555_),
    .S(mem_la_wdata[4]),
    .X(_19831_));
 sky130_fd_sc_hd__mux2_1 _38820_ (.A0(_00148_),
    .A1(_00140_),
    .S(mem_la_wdata[1]),
    .X(_00149_));
 sky130_fd_sc_hd__mux2_1 _38821_ (.A0(_00149_),
    .A1(_00133_),
    .S(mem_la_wdata[2]),
    .X(_00150_));
 sky130_fd_sc_hd__mux2_1 _38822_ (.A0(_00150_),
    .A1(_00113_),
    .S(mem_la_wdata[3]),
    .X(_00151_));
 sky130_fd_sc_hd__mux2_1 _38823_ (.A0(_00151_),
    .A1(_02556_),
    .S(mem_la_wdata[4]),
    .X(_19832_));
 sky130_fd_sc_hd__mux2_1 _38824_ (.A0(pcpi_rs1[30]),
    .A1(pcpi_rs1[29]),
    .S(mem_la_wdata[0]),
    .X(_00152_));
 sky130_fd_sc_hd__mux2_1 _38825_ (.A0(_00152_),
    .A1(_00144_),
    .S(mem_la_wdata[1]),
    .X(_00153_));
 sky130_fd_sc_hd__mux2_1 _38826_ (.A0(_00153_),
    .A1(_00137_),
    .S(mem_la_wdata[2]),
    .X(_00154_));
 sky130_fd_sc_hd__mux2_1 _38827_ (.A0(_00154_),
    .A1(_00119_),
    .S(mem_la_wdata[3]),
    .X(_00155_));
 sky130_fd_sc_hd__mux2_1 _38828_ (.A0(_00155_),
    .A1(_02557_),
    .S(mem_la_wdata[4]),
    .X(_19833_));
 sky130_fd_sc_hd__mux2_1 _38829_ (.A0(pcpi_rs1[31]),
    .A1(pcpi_rs1[30]),
    .S(mem_la_wdata[0]),
    .X(_00156_));
 sky130_fd_sc_hd__mux2_1 _38830_ (.A0(_00156_),
    .A1(_00148_),
    .S(mem_la_wdata[1]),
    .X(_00157_));
 sky130_fd_sc_hd__mux2_1 _38831_ (.A0(_00157_),
    .A1(_00141_),
    .S(mem_la_wdata[2]),
    .X(_00158_));
 sky130_fd_sc_hd__mux2_1 _38832_ (.A0(_00158_),
    .A1(_00125_),
    .S(mem_la_wdata[3]),
    .X(_00159_));
 sky130_fd_sc_hd__mux2_1 _38833_ (.A0(_00159_),
    .A1(_02558_),
    .S(mem_la_wdata[4]),
    .X(_19834_));
 sky130_fd_sc_hd__mux2_1 _38834_ (.A0(pcpi_rs1[0]),
    .A1(pcpi_rs1[1]),
    .S(mem_la_wdata[0]),
    .X(_00160_));
 sky130_fd_sc_hd__mux2_1 _38835_ (.A0(_00160_),
    .A1(_00161_),
    .S(mem_la_wdata[1]),
    .X(_00162_));
 sky130_fd_sc_hd__mux2_1 _38836_ (.A0(_00162_),
    .A1(_00165_),
    .S(mem_la_wdata[2]),
    .X(_00166_));
 sky130_fd_sc_hd__mux2_1 _38837_ (.A0(_00166_),
    .A1(_00173_),
    .S(mem_la_wdata[3]),
    .X(_00174_));
 sky130_fd_sc_hd__mux2_1 _38838_ (.A0(_00174_),
    .A1(_00189_),
    .S(mem_la_wdata[4]),
    .X(_19835_));
 sky130_fd_sc_hd__mux2_1 _38839_ (.A0(pcpi_rs1[1]),
    .A1(pcpi_rs1[2]),
    .S(mem_la_wdata[0]),
    .X(_00190_));
 sky130_fd_sc_hd__mux2_1 _38840_ (.A0(_00190_),
    .A1(_00191_),
    .S(mem_la_wdata[1]),
    .X(_00192_));
 sky130_fd_sc_hd__mux2_1 _38841_ (.A0(_00192_),
    .A1(_00195_),
    .S(mem_la_wdata[2]),
    .X(_00196_));
 sky130_fd_sc_hd__mux2_1 _38842_ (.A0(_00196_),
    .A1(_00203_),
    .S(mem_la_wdata[3]),
    .X(_00204_));
 sky130_fd_sc_hd__mux2_1 _38843_ (.A0(_00204_),
    .A1(_00220_),
    .S(mem_la_wdata[4]),
    .X(_19846_));
 sky130_fd_sc_hd__mux2_1 _38844_ (.A0(_00161_),
    .A1(_00163_),
    .S(mem_la_wdata[1]),
    .X(_00221_));
 sky130_fd_sc_hd__mux2_1 _38845_ (.A0(_00221_),
    .A1(_00222_),
    .S(mem_la_wdata[2]),
    .X(_00223_));
 sky130_fd_sc_hd__mux2_1 _38846_ (.A0(_00223_),
    .A1(_00226_),
    .S(mem_la_wdata[3]),
    .X(_00227_));
 sky130_fd_sc_hd__mux2_1 _38847_ (.A0(_00227_),
    .A1(_00234_),
    .S(mem_la_wdata[4]),
    .X(_19857_));
 sky130_fd_sc_hd__mux2_1 _38848_ (.A0(_00191_),
    .A1(_00193_),
    .S(mem_la_wdata[1]),
    .X(_00235_));
 sky130_fd_sc_hd__mux2_1 _38849_ (.A0(_00235_),
    .A1(_00236_),
    .S(mem_la_wdata[2]),
    .X(_00237_));
 sky130_fd_sc_hd__mux2_1 _38850_ (.A0(_00237_),
    .A1(_00240_),
    .S(mem_la_wdata[3]),
    .X(_00241_));
 sky130_fd_sc_hd__mux2_1 _38851_ (.A0(_00241_),
    .A1(_00248_),
    .S(mem_la_wdata[4]),
    .X(_19860_));
 sky130_fd_sc_hd__mux2_1 _38852_ (.A0(_00165_),
    .A1(_00169_),
    .S(mem_la_wdata[2]),
    .X(_00249_));
 sky130_fd_sc_hd__mux2_1 _38853_ (.A0(_00249_),
    .A1(_00250_),
    .S(mem_la_wdata[3]),
    .X(_00251_));
 sky130_fd_sc_hd__mux2_1 _38854_ (.A0(_00251_),
    .A1(_00254_),
    .S(mem_la_wdata[4]),
    .X(_19861_));
 sky130_fd_sc_hd__mux2_1 _38855_ (.A0(_00195_),
    .A1(_00199_),
    .S(mem_la_wdata[2]),
    .X(_00255_));
 sky130_fd_sc_hd__mux2_1 _38856_ (.A0(_00255_),
    .A1(_00256_),
    .S(mem_la_wdata[3]),
    .X(_00257_));
 sky130_fd_sc_hd__mux2_1 _38857_ (.A0(_00257_),
    .A1(_00260_),
    .S(mem_la_wdata[4]),
    .X(_19862_));
 sky130_fd_sc_hd__mux2_1 _38858_ (.A0(_00222_),
    .A1(_00224_),
    .S(mem_la_wdata[2]),
    .X(_00261_));
 sky130_fd_sc_hd__mux2_1 _38859_ (.A0(_00261_),
    .A1(_00262_),
    .S(mem_la_wdata[3]),
    .X(_00263_));
 sky130_fd_sc_hd__mux2_1 _38860_ (.A0(_00263_),
    .A1(_00266_),
    .S(mem_la_wdata[4]),
    .X(_19863_));
 sky130_fd_sc_hd__mux2_1 _38861_ (.A0(_00236_),
    .A1(_00238_),
    .S(mem_la_wdata[2]),
    .X(_00267_));
 sky130_fd_sc_hd__mux2_1 _38862_ (.A0(_00267_),
    .A1(_00268_),
    .S(mem_la_wdata[3]),
    .X(_00269_));
 sky130_fd_sc_hd__mux2_1 _38863_ (.A0(_00269_),
    .A1(_00272_),
    .S(mem_la_wdata[4]),
    .X(_19864_));
 sky130_fd_sc_hd__mux2_1 _38864_ (.A0(_00173_),
    .A1(_00181_),
    .S(mem_la_wdata[3]),
    .X(_00273_));
 sky130_fd_sc_hd__mux2_1 _38865_ (.A0(_00273_),
    .A1(_00274_),
    .S(mem_la_wdata[4]),
    .X(_19865_));
 sky130_fd_sc_hd__mux2_1 _38866_ (.A0(_00203_),
    .A1(_00211_),
    .S(mem_la_wdata[3]),
    .X(_00275_));
 sky130_fd_sc_hd__mux2_1 _38867_ (.A0(_00275_),
    .A1(_00276_),
    .S(mem_la_wdata[4]),
    .X(_19866_));
 sky130_fd_sc_hd__mux2_1 _38868_ (.A0(_00226_),
    .A1(_00230_),
    .S(mem_la_wdata[3]),
    .X(_00277_));
 sky130_fd_sc_hd__mux2_1 _38869_ (.A0(_00277_),
    .A1(_00278_),
    .S(mem_la_wdata[4]),
    .X(_19836_));
 sky130_fd_sc_hd__mux2_1 _38870_ (.A0(_00240_),
    .A1(_00244_),
    .S(mem_la_wdata[3]),
    .X(_00279_));
 sky130_fd_sc_hd__mux2_1 _38871_ (.A0(_00279_),
    .A1(_00280_),
    .S(mem_la_wdata[4]),
    .X(_19837_));
 sky130_fd_sc_hd__mux2_1 _38872_ (.A0(_00250_),
    .A1(_00252_),
    .S(mem_la_wdata[3]),
    .X(_00281_));
 sky130_fd_sc_hd__mux2_1 _38873_ (.A0(_00281_),
    .A1(_00282_),
    .S(mem_la_wdata[4]),
    .X(_19838_));
 sky130_fd_sc_hd__mux2_1 _38874_ (.A0(_00256_),
    .A1(_00258_),
    .S(mem_la_wdata[3]),
    .X(_00283_));
 sky130_fd_sc_hd__mux2_1 _38875_ (.A0(_00283_),
    .A1(_00284_),
    .S(mem_la_wdata[4]),
    .X(_19839_));
 sky130_fd_sc_hd__mux2_1 _38876_ (.A0(_00262_),
    .A1(_00264_),
    .S(mem_la_wdata[3]),
    .X(_00285_));
 sky130_fd_sc_hd__mux2_1 _38877_ (.A0(_00285_),
    .A1(_00286_),
    .S(mem_la_wdata[4]),
    .X(_19840_));
 sky130_fd_sc_hd__mux2_1 _38878_ (.A0(_00268_),
    .A1(_00270_),
    .S(mem_la_wdata[3]),
    .X(_00287_));
 sky130_fd_sc_hd__mux2_1 _38879_ (.A0(_00287_),
    .A1(_00288_),
    .S(mem_la_wdata[4]),
    .X(_19841_));
 sky130_fd_sc_hd__mux2_1 _38880_ (.A0(_00189_),
    .A1(_00216_),
    .S(mem_la_wdata[4]),
    .X(_19842_));
 sky130_fd_sc_hd__mux2_1 _38881_ (.A0(_00220_),
    .A1(_00216_),
    .S(mem_la_wdata[4]),
    .X(_19843_));
 sky130_fd_sc_hd__mux2_1 _38882_ (.A0(_00234_),
    .A1(_00216_),
    .S(mem_la_wdata[4]),
    .X(_19844_));
 sky130_fd_sc_hd__mux2_1 _38883_ (.A0(_00248_),
    .A1(_00216_),
    .S(mem_la_wdata[4]),
    .X(_19845_));
 sky130_fd_sc_hd__mux2_1 _38884_ (.A0(_00254_),
    .A1(_00216_),
    .S(mem_la_wdata[4]),
    .X(_19847_));
 sky130_fd_sc_hd__mux2_1 _38885_ (.A0(_00260_),
    .A1(_00216_),
    .S(mem_la_wdata[4]),
    .X(_19848_));
 sky130_fd_sc_hd__mux2_1 _38886_ (.A0(_00266_),
    .A1(_00216_),
    .S(mem_la_wdata[4]),
    .X(_19849_));
 sky130_fd_sc_hd__mux2_1 _38887_ (.A0(_00272_),
    .A1(_00216_),
    .S(mem_la_wdata[4]),
    .X(_19850_));
 sky130_fd_sc_hd__mux2_1 _38888_ (.A0(_00274_),
    .A1(_00216_),
    .S(mem_la_wdata[4]),
    .X(_19851_));
 sky130_fd_sc_hd__mux2_1 _38889_ (.A0(_00276_),
    .A1(_00216_),
    .S(mem_la_wdata[4]),
    .X(_19852_));
 sky130_fd_sc_hd__mux2_1 _38890_ (.A0(_00278_),
    .A1(_00216_),
    .S(mem_la_wdata[4]),
    .X(_19853_));
 sky130_fd_sc_hd__mux2_1 _38891_ (.A0(_00280_),
    .A1(_00216_),
    .S(mem_la_wdata[4]),
    .X(_19854_));
 sky130_fd_sc_hd__mux2_1 _38892_ (.A0(_00282_),
    .A1(_00216_),
    .S(mem_la_wdata[4]),
    .X(_19855_));
 sky130_fd_sc_hd__mux2_1 _38893_ (.A0(_00284_),
    .A1(_00216_),
    .S(mem_la_wdata[4]),
    .X(_19856_));
 sky130_fd_sc_hd__mux2_1 _38894_ (.A0(_00286_),
    .A1(_00216_),
    .S(mem_la_wdata[4]),
    .X(_19858_));
 sky130_fd_sc_hd__mux2_1 _38895_ (.A0(_00288_),
    .A1(_00216_),
    .S(mem_la_wdata[4]),
    .X(_19859_));
 sky130_fd_sc_hd__mux2_1 _38896_ (.A0(_01697_),
    .A1(_01698_),
    .S(\irq_state[1] ),
    .X(_01699_));
 sky130_fd_sc_hd__mux2_1 _38897_ (.A0(_01705_),
    .A1(_01699_),
    .S(_01700_),
    .X(_19818_));
 sky130_fd_sc_hd__mux2_1 _38898_ (.A0(_01720_),
    .A1(\irq_pending[0] ),
    .S(_01706_),
    .X(_19784_));
 sky130_fd_sc_hd__mux2_1 _38899_ (.A0(_01733_),
    .A1(\irq_pending[1] ),
    .S(_01706_),
    .X(_19795_));
 sky130_fd_sc_hd__mux2_1 _38900_ (.A0(_01746_),
    .A1(\irq_pending[2] ),
    .S(_01706_),
    .X(_19806_));
 sky130_fd_sc_hd__mux2_1 _38901_ (.A0(_01759_),
    .A1(\irq_pending[3] ),
    .S(_01706_),
    .X(_19809_));
 sky130_fd_sc_hd__mux2_1 _38902_ (.A0(_01772_),
    .A1(\irq_pending[4] ),
    .S(_01706_),
    .X(_19810_));
 sky130_fd_sc_hd__mux2_1 _38903_ (.A0(_01785_),
    .A1(\irq_pending[5] ),
    .S(_01706_),
    .X(_19811_));
 sky130_fd_sc_hd__mux2_1 _38904_ (.A0(_01798_),
    .A1(\irq_pending[6] ),
    .S(_01706_),
    .X(_19812_));
 sky130_fd_sc_hd__mux2_1 _38905_ (.A0(_01811_),
    .A1(\irq_pending[7] ),
    .S(_01706_),
    .X(_19813_));
 sky130_fd_sc_hd__mux2_1 _38906_ (.A0(_01825_),
    .A1(\irq_pending[8] ),
    .S(_01706_),
    .X(_19814_));
 sky130_fd_sc_hd__mux2_1 _38907_ (.A0(_01838_),
    .A1(\irq_pending[9] ),
    .S(_01706_),
    .X(_19815_));
 sky130_fd_sc_hd__mux2_1 _38908_ (.A0(_01851_),
    .A1(\irq_pending[10] ),
    .S(_01706_),
    .X(_19785_));
 sky130_fd_sc_hd__mux2_1 _38909_ (.A0(_01864_),
    .A1(\irq_pending[11] ),
    .S(_01706_),
    .X(_19786_));
 sky130_fd_sc_hd__mux2_1 _38910_ (.A0(_01877_),
    .A1(\irq_pending[12] ),
    .S(_01706_),
    .X(_19787_));
 sky130_fd_sc_hd__mux2_1 _38911_ (.A0(_01890_),
    .A1(\irq_pending[13] ),
    .S(_01706_),
    .X(_19788_));
 sky130_fd_sc_hd__mux2_1 _38912_ (.A0(_01903_),
    .A1(\irq_pending[14] ),
    .S(_01706_),
    .X(_19789_));
 sky130_fd_sc_hd__mux2_1 _38913_ (.A0(_01916_),
    .A1(\irq_pending[15] ),
    .S(_01706_),
    .X(_19790_));
 sky130_fd_sc_hd__mux2_1 _38914_ (.A0(_01925_),
    .A1(\irq_pending[16] ),
    .S(_01706_),
    .X(_19791_));
 sky130_fd_sc_hd__mux2_1 _38915_ (.A0(_01934_),
    .A1(\irq_pending[17] ),
    .S(_01706_),
    .X(_19792_));
 sky130_fd_sc_hd__mux2_1 _38916_ (.A0(_01943_),
    .A1(\irq_pending[18] ),
    .S(_01706_),
    .X(_19793_));
 sky130_fd_sc_hd__mux2_1 _38917_ (.A0(_01952_),
    .A1(\irq_pending[19] ),
    .S(_01706_),
    .X(_19794_));
 sky130_fd_sc_hd__mux2_1 _38918_ (.A0(_01961_),
    .A1(\irq_pending[20] ),
    .S(_01706_),
    .X(_19796_));
 sky130_fd_sc_hd__mux2_1 _38919_ (.A0(_01970_),
    .A1(\irq_pending[21] ),
    .S(_01706_),
    .X(_19797_));
 sky130_fd_sc_hd__mux2_1 _38920_ (.A0(_01979_),
    .A1(\irq_pending[22] ),
    .S(_01706_),
    .X(_19798_));
 sky130_fd_sc_hd__mux2_1 _38921_ (.A0(_01988_),
    .A1(\irq_pending[23] ),
    .S(_01706_),
    .X(_19799_));
 sky130_fd_sc_hd__mux2_1 _38922_ (.A0(_01997_),
    .A1(\irq_pending[24] ),
    .S(_01706_),
    .X(_19800_));
 sky130_fd_sc_hd__mux2_1 _38923_ (.A0(_02006_),
    .A1(\irq_pending[25] ),
    .S(_01706_),
    .X(_19801_));
 sky130_fd_sc_hd__mux2_1 _38924_ (.A0(_02015_),
    .A1(\irq_pending[26] ),
    .S(_01706_),
    .X(_19802_));
 sky130_fd_sc_hd__mux2_1 _38925_ (.A0(_02024_),
    .A1(\irq_pending[27] ),
    .S(_01706_),
    .X(_19803_));
 sky130_fd_sc_hd__mux2_1 _38926_ (.A0(_02033_),
    .A1(\irq_pending[28] ),
    .S(_01706_),
    .X(_19804_));
 sky130_fd_sc_hd__mux2_1 _38927_ (.A0(_02042_),
    .A1(\irq_pending[29] ),
    .S(_01706_),
    .X(_19805_));
 sky130_fd_sc_hd__mux2_1 _38928_ (.A0(_02051_),
    .A1(\irq_pending[30] ),
    .S(_01706_),
    .X(_19807_));
 sky130_fd_sc_hd__mux2_1 _38929_ (.A0(_02060_),
    .A1(\irq_pending[31] ),
    .S(_01706_),
    .X(_19808_));
 sky130_fd_sc_hd__mux2_1 _38930_ (.A0(_02061_),
    .A1(\cpu_state[2] ),
    .S(_02542_),
    .X(_19779_));
 sky130_fd_sc_hd__mux2_1 _38931_ (.A0(\decoded_rd[0] ),
    .A1(\irq_state[0] ),
    .S(_00308_),
    .X(_19778_));
 sky130_fd_sc_hd__mux2_1 _38932_ (.A0(_02062_),
    .A1(_02065_),
    .S(_02542_),
    .X(_19816_));
 sky130_fd_sc_hd__mux2_1 _38933_ (.A0(_02068_),
    .A1(_02066_),
    .S(_02067_),
    .X(_19817_));
 sky130_fd_sc_hd__mux2_1 _38934_ (.A0(_02166_),
    .A1(_00291_),
    .S(_00290_),
    .X(_19780_));
 sky130_fd_sc_hd__mux2_1 _38935_ (.A0(_02166_),
    .A1(mem_do_wdata),
    .S(_00290_),
    .X(_19781_));
 sky130_fd_sc_hd__mux2_1 _38936_ (.A0(_00271_),
    .A1(_00216_),
    .S(mem_la_wdata[3]),
    .X(_00288_));
 sky130_fd_sc_hd__mux2_1 _38937_ (.A0(_00265_),
    .A1(_00216_),
    .S(mem_la_wdata[3]),
    .X(_00286_));
 sky130_fd_sc_hd__mux2_1 _38938_ (.A0(_00259_),
    .A1(_00216_),
    .S(mem_la_wdata[3]),
    .X(_00284_));
 sky130_fd_sc_hd__mux2_1 _38939_ (.A0(_00253_),
    .A1(_00216_),
    .S(mem_la_wdata[3]),
    .X(_00282_));
 sky130_fd_sc_hd__mux2_1 _38940_ (.A0(_00247_),
    .A1(_00216_),
    .S(mem_la_wdata[3]),
    .X(_00280_));
 sky130_fd_sc_hd__mux2_1 _38941_ (.A0(_00233_),
    .A1(_00216_),
    .S(mem_la_wdata[3]),
    .X(_00278_));
 sky130_fd_sc_hd__mux2_1 _38942_ (.A0(_00219_),
    .A1(_00216_),
    .S(mem_la_wdata[3]),
    .X(_00276_));
 sky130_fd_sc_hd__mux2_1 _38943_ (.A0(_00188_),
    .A1(_00216_),
    .S(mem_la_wdata[3]),
    .X(_00274_));
 sky130_fd_sc_hd__mux2_1 _38944_ (.A0(_00270_),
    .A1(_00271_),
    .S(mem_la_wdata[3]),
    .X(_00272_));
 sky130_fd_sc_hd__mux2_1 _38945_ (.A0(_00246_),
    .A1(_00216_),
    .S(mem_la_wdata[2]),
    .X(_00271_));
 sky130_fd_sc_hd__mux2_1 _38946_ (.A0(_00243_),
    .A1(_00245_),
    .S(mem_la_wdata[2]),
    .X(_00270_));
 sky130_fd_sc_hd__mux2_1 _38947_ (.A0(_00239_),
    .A1(_00242_),
    .S(mem_la_wdata[2]),
    .X(_00268_));
 sky130_fd_sc_hd__mux2_1 _38948_ (.A0(_00264_),
    .A1(_00265_),
    .S(mem_la_wdata[3]),
    .X(_00266_));
 sky130_fd_sc_hd__mux2_1 _38949_ (.A0(_00232_),
    .A1(_00216_),
    .S(mem_la_wdata[2]),
    .X(_00265_));
 sky130_fd_sc_hd__mux2_1 _38950_ (.A0(_00229_),
    .A1(_00231_),
    .S(mem_la_wdata[2]),
    .X(_00264_));
 sky130_fd_sc_hd__mux2_1 _38951_ (.A0(_00225_),
    .A1(_00228_),
    .S(mem_la_wdata[2]),
    .X(_00262_));
 sky130_fd_sc_hd__mux2_1 _38952_ (.A0(_00258_),
    .A1(_00259_),
    .S(mem_la_wdata[3]),
    .X(_00260_));
 sky130_fd_sc_hd__mux2_1 _38953_ (.A0(_00218_),
    .A1(_00216_),
    .S(mem_la_wdata[2]),
    .X(_00259_));
 sky130_fd_sc_hd__mux2_1 _38954_ (.A0(_00210_),
    .A1(_00214_),
    .S(mem_la_wdata[2]),
    .X(_00258_));
 sky130_fd_sc_hd__mux2_1 _38955_ (.A0(_00202_),
    .A1(_00207_),
    .S(mem_la_wdata[2]),
    .X(_00256_));
 sky130_fd_sc_hd__mux2_1 _38956_ (.A0(_00252_),
    .A1(_00253_),
    .S(mem_la_wdata[3]),
    .X(_00254_));
 sky130_fd_sc_hd__mux2_1 _38957_ (.A0(_00187_),
    .A1(_00216_),
    .S(mem_la_wdata[2]),
    .X(_00253_));
 sky130_fd_sc_hd__mux2_1 _38958_ (.A0(_00180_),
    .A1(_00184_),
    .S(mem_la_wdata[2]),
    .X(_00252_));
 sky130_fd_sc_hd__mux2_1 _38959_ (.A0(_00172_),
    .A1(_00177_),
    .S(mem_la_wdata[2]),
    .X(_00250_));
 sky130_fd_sc_hd__mux2_1 _38960_ (.A0(_00244_),
    .A1(_00247_),
    .S(mem_la_wdata[3]),
    .X(_00248_));
 sky130_fd_sc_hd__mux2_1 _38961_ (.A0(_00245_),
    .A1(_00246_),
    .S(mem_la_wdata[2]),
    .X(_00247_));
 sky130_fd_sc_hd__mux2_1 _38962_ (.A0(_00217_),
    .A1(_00216_),
    .S(mem_la_wdata[1]),
    .X(_00246_));
 sky130_fd_sc_hd__mux2_1 _38963_ (.A0(_00213_),
    .A1(_00215_),
    .S(mem_la_wdata[1]),
    .X(_00245_));
 sky130_fd_sc_hd__mux2_1 _38964_ (.A0(_00242_),
    .A1(_00243_),
    .S(mem_la_wdata[2]),
    .X(_00244_));
 sky130_fd_sc_hd__mux2_1 _38965_ (.A0(_00209_),
    .A1(_00212_),
    .S(mem_la_wdata[1]),
    .X(_00243_));
 sky130_fd_sc_hd__mux2_1 _38966_ (.A0(_00206_),
    .A1(_00208_),
    .S(mem_la_wdata[1]),
    .X(_00242_));
 sky130_fd_sc_hd__mux2_1 _38967_ (.A0(_00238_),
    .A1(_00239_),
    .S(mem_la_wdata[2]),
    .X(_00240_));
 sky130_fd_sc_hd__mux2_1 _38968_ (.A0(_00201_),
    .A1(_00205_),
    .S(mem_la_wdata[1]),
    .X(_00239_));
 sky130_fd_sc_hd__mux2_1 _38969_ (.A0(_00198_),
    .A1(_00200_),
    .S(mem_la_wdata[1]),
    .X(_00238_));
 sky130_fd_sc_hd__mux2_1 _38970_ (.A0(_00194_),
    .A1(_00197_),
    .S(mem_la_wdata[1]),
    .X(_00236_));
 sky130_fd_sc_hd__mux2_1 _38971_ (.A0(_00230_),
    .A1(_00233_),
    .S(mem_la_wdata[3]),
    .X(_00234_));
 sky130_fd_sc_hd__mux2_1 _38972_ (.A0(_00231_),
    .A1(_00232_),
    .S(mem_la_wdata[2]),
    .X(_00233_));
 sky130_fd_sc_hd__mux2_1 _38973_ (.A0(_00186_),
    .A1(_00216_),
    .S(mem_la_wdata[1]),
    .X(_00232_));
 sky130_fd_sc_hd__mux2_1 _38974_ (.A0(_00183_),
    .A1(_00185_),
    .S(mem_la_wdata[1]),
    .X(_00231_));
 sky130_fd_sc_hd__mux2_1 _38975_ (.A0(_00228_),
    .A1(_00229_),
    .S(mem_la_wdata[2]),
    .X(_00230_));
 sky130_fd_sc_hd__mux2_1 _38976_ (.A0(_00179_),
    .A1(_00182_),
    .S(mem_la_wdata[1]),
    .X(_00229_));
 sky130_fd_sc_hd__mux2_1 _38977_ (.A0(_00176_),
    .A1(_00178_),
    .S(mem_la_wdata[1]),
    .X(_00228_));
 sky130_fd_sc_hd__mux2_1 _38978_ (.A0(_00224_),
    .A1(_00225_),
    .S(mem_la_wdata[2]),
    .X(_00226_));
 sky130_fd_sc_hd__mux2_1 _38979_ (.A0(_00171_),
    .A1(_00175_),
    .S(mem_la_wdata[1]),
    .X(_00225_));
 sky130_fd_sc_hd__mux2_1 _38980_ (.A0(_00168_),
    .A1(_00170_),
    .S(mem_la_wdata[1]),
    .X(_00224_));
 sky130_fd_sc_hd__mux2_1 _38981_ (.A0(_00164_),
    .A1(_00167_),
    .S(mem_la_wdata[1]),
    .X(_00222_));
 sky130_fd_sc_hd__mux2_1 _38982_ (.A0(_00211_),
    .A1(_00219_),
    .S(mem_la_wdata[3]),
    .X(_00220_));
 sky130_fd_sc_hd__mux2_1 _38983_ (.A0(_00214_),
    .A1(_00218_),
    .S(mem_la_wdata[2]),
    .X(_00219_));
 sky130_fd_sc_hd__mux2_1 _38984_ (.A0(_00215_),
    .A1(_00217_),
    .S(mem_la_wdata[1]),
    .X(_00218_));
 sky130_fd_sc_hd__mux2_1 _38985_ (.A0(pcpi_rs1[31]),
    .A1(_00216_),
    .S(mem_la_wdata[0]),
    .X(_00217_));
 sky130_fd_sc_hd__mux2_1 _38986_ (.A0(pcpi_rs1[29]),
    .A1(pcpi_rs1[30]),
    .S(mem_la_wdata[0]),
    .X(_00215_));
 sky130_fd_sc_hd__mux2_1 _38987_ (.A0(_00212_),
    .A1(_00213_),
    .S(mem_la_wdata[1]),
    .X(_00214_));
 sky130_fd_sc_hd__mux2_1 _38988_ (.A0(pcpi_rs1[27]),
    .A1(pcpi_rs1[28]),
    .S(mem_la_wdata[0]),
    .X(_00213_));
 sky130_fd_sc_hd__mux2_1 _38989_ (.A0(pcpi_rs1[25]),
    .A1(pcpi_rs1[26]),
    .S(mem_la_wdata[0]),
    .X(_00212_));
 sky130_fd_sc_hd__mux2_1 _38990_ (.A0(_00207_),
    .A1(_00210_),
    .S(mem_la_wdata[2]),
    .X(_00211_));
 sky130_fd_sc_hd__mux2_1 _38991_ (.A0(_00208_),
    .A1(_00209_),
    .S(mem_la_wdata[1]),
    .X(_00210_));
 sky130_fd_sc_hd__mux2_1 _38992_ (.A0(pcpi_rs1[23]),
    .A1(pcpi_rs1[24]),
    .S(mem_la_wdata[0]),
    .X(_00209_));
 sky130_fd_sc_hd__mux2_1 _38993_ (.A0(pcpi_rs1[21]),
    .A1(pcpi_rs1[22]),
    .S(mem_la_wdata[0]),
    .X(_00208_));
 sky130_fd_sc_hd__mux2_1 _38994_ (.A0(_00205_),
    .A1(_00206_),
    .S(mem_la_wdata[1]),
    .X(_00207_));
 sky130_fd_sc_hd__mux2_1 _38995_ (.A0(pcpi_rs1[19]),
    .A1(pcpi_rs1[20]),
    .S(mem_la_wdata[0]),
    .X(_00206_));
 sky130_fd_sc_hd__mux2_1 _38996_ (.A0(pcpi_rs1[17]),
    .A1(pcpi_rs1[18]),
    .S(mem_la_wdata[0]),
    .X(_00205_));
 sky130_fd_sc_hd__mux2_1 _38997_ (.A0(_00199_),
    .A1(_00202_),
    .S(mem_la_wdata[2]),
    .X(_00203_));
 sky130_fd_sc_hd__mux2_1 _38998_ (.A0(_00200_),
    .A1(_00201_),
    .S(mem_la_wdata[1]),
    .X(_00202_));
 sky130_fd_sc_hd__mux2_1 _38999_ (.A0(pcpi_rs1[15]),
    .A1(pcpi_rs1[16]),
    .S(mem_la_wdata[0]),
    .X(_00201_));
 sky130_fd_sc_hd__mux2_1 _39000_ (.A0(pcpi_rs1[13]),
    .A1(pcpi_rs1[14]),
    .S(mem_la_wdata[0]),
    .X(_00200_));
 sky130_fd_sc_hd__mux2_1 _39001_ (.A0(_00197_),
    .A1(_00198_),
    .S(mem_la_wdata[1]),
    .X(_00199_));
 sky130_fd_sc_hd__mux2_1 _39002_ (.A0(pcpi_rs1[11]),
    .A1(pcpi_rs1[12]),
    .S(mem_la_wdata[0]),
    .X(_00198_));
 sky130_fd_sc_hd__mux2_1 _39003_ (.A0(pcpi_rs1[9]),
    .A1(pcpi_rs1[10]),
    .S(mem_la_wdata[0]),
    .X(_00197_));
 sky130_fd_sc_hd__mux2_1 _39004_ (.A0(_00193_),
    .A1(_00194_),
    .S(mem_la_wdata[1]),
    .X(_00195_));
 sky130_fd_sc_hd__mux2_1 _39005_ (.A0(pcpi_rs1[7]),
    .A1(pcpi_rs1[8]),
    .S(mem_la_wdata[0]),
    .X(_00194_));
 sky130_fd_sc_hd__mux2_1 _39006_ (.A0(pcpi_rs1[5]),
    .A1(pcpi_rs1[6]),
    .S(mem_la_wdata[0]),
    .X(_00193_));
 sky130_fd_sc_hd__mux2_1 _39007_ (.A0(pcpi_rs1[3]),
    .A1(pcpi_rs1[4]),
    .S(mem_la_wdata[0]),
    .X(_00191_));
 sky130_fd_sc_hd__mux2_1 _39008_ (.A0(_00181_),
    .A1(_00188_),
    .S(mem_la_wdata[3]),
    .X(_00189_));
 sky130_fd_sc_hd__mux2_1 _39009_ (.A0(_00184_),
    .A1(_00187_),
    .S(mem_la_wdata[2]),
    .X(_00188_));
 sky130_fd_sc_hd__mux2_1 _39010_ (.A0(_00185_),
    .A1(_00186_),
    .S(mem_la_wdata[1]),
    .X(_00187_));
 sky130_fd_sc_hd__mux2_1 _39011_ (.A0(pcpi_rs1[30]),
    .A1(pcpi_rs1[31]),
    .S(mem_la_wdata[0]),
    .X(_00186_));
 sky130_fd_sc_hd__mux2_1 _39012_ (.A0(pcpi_rs1[28]),
    .A1(pcpi_rs1[29]),
    .S(mem_la_wdata[0]),
    .X(_00185_));
 sky130_fd_sc_hd__mux2_1 _39013_ (.A0(_00182_),
    .A1(_00183_),
    .S(mem_la_wdata[1]),
    .X(_00184_));
 sky130_fd_sc_hd__mux2_1 _39014_ (.A0(pcpi_rs1[26]),
    .A1(pcpi_rs1[27]),
    .S(mem_la_wdata[0]),
    .X(_00183_));
 sky130_fd_sc_hd__mux2_1 _39015_ (.A0(pcpi_rs1[24]),
    .A1(pcpi_rs1[25]),
    .S(mem_la_wdata[0]),
    .X(_00182_));
 sky130_fd_sc_hd__mux2_1 _39016_ (.A0(_00177_),
    .A1(_00180_),
    .S(mem_la_wdata[2]),
    .X(_00181_));
 sky130_fd_sc_hd__mux2_1 _39017_ (.A0(_00178_),
    .A1(_00179_),
    .S(mem_la_wdata[1]),
    .X(_00180_));
 sky130_fd_sc_hd__mux2_1 _39018_ (.A0(pcpi_rs1[22]),
    .A1(pcpi_rs1[23]),
    .S(mem_la_wdata[0]),
    .X(_00179_));
 sky130_fd_sc_hd__mux2_1 _39019_ (.A0(pcpi_rs1[20]),
    .A1(pcpi_rs1[21]),
    .S(mem_la_wdata[0]),
    .X(_00178_));
 sky130_fd_sc_hd__mux2_1 _39020_ (.A0(_00175_),
    .A1(_00176_),
    .S(mem_la_wdata[1]),
    .X(_00177_));
 sky130_fd_sc_hd__mux2_1 _39021_ (.A0(pcpi_rs1[18]),
    .A1(pcpi_rs1[19]),
    .S(mem_la_wdata[0]),
    .X(_00176_));
 sky130_fd_sc_hd__mux2_1 _39022_ (.A0(pcpi_rs1[16]),
    .A1(pcpi_rs1[17]),
    .S(mem_la_wdata[0]),
    .X(_00175_));
 sky130_fd_sc_hd__mux2_1 _39023_ (.A0(_00169_),
    .A1(_00172_),
    .S(mem_la_wdata[2]),
    .X(_00173_));
 sky130_fd_sc_hd__mux2_1 _39024_ (.A0(_00170_),
    .A1(_00171_),
    .S(mem_la_wdata[1]),
    .X(_00172_));
 sky130_fd_sc_hd__mux2_1 _39025_ (.A0(pcpi_rs1[14]),
    .A1(pcpi_rs1[15]),
    .S(mem_la_wdata[0]),
    .X(_00171_));
 sky130_fd_sc_hd__mux2_1 _39026_ (.A0(pcpi_rs1[12]),
    .A1(pcpi_rs1[13]),
    .S(mem_la_wdata[0]),
    .X(_00170_));
 sky130_fd_sc_hd__mux2_1 _39027_ (.A0(_00167_),
    .A1(_00168_),
    .S(mem_la_wdata[1]),
    .X(_00169_));
 sky130_fd_sc_hd__mux2_1 _39028_ (.A0(pcpi_rs1[10]),
    .A1(pcpi_rs1[11]),
    .S(mem_la_wdata[0]),
    .X(_00168_));
 sky130_fd_sc_hd__mux2_1 _39029_ (.A0(pcpi_rs1[8]),
    .A1(pcpi_rs1[9]),
    .S(mem_la_wdata[0]),
    .X(_00167_));
 sky130_fd_sc_hd__mux2_1 _39030_ (.A0(_00163_),
    .A1(_00164_),
    .S(mem_la_wdata[1]),
    .X(_00165_));
 sky130_fd_sc_hd__mux2_1 _39031_ (.A0(pcpi_rs1[6]),
    .A1(pcpi_rs1[7]),
    .S(mem_la_wdata[0]),
    .X(_00164_));
 sky130_fd_sc_hd__mux2_1 _39032_ (.A0(pcpi_rs1[4]),
    .A1(pcpi_rs1[5]),
    .S(mem_la_wdata[0]),
    .X(_00163_));
 sky130_fd_sc_hd__mux2_1 _39033_ (.A0(pcpi_rs1[2]),
    .A1(pcpi_rs1[3]),
    .S(mem_la_wdata[0]),
    .X(_00161_));
 sky130_fd_sc_hd__mux2_1 _39034_ (.A0(pcpi_rs1[29]),
    .A1(pcpi_rs1[28]),
    .S(mem_la_wdata[0]),
    .X(_00148_));
 sky130_fd_sc_hd__mux2_1 _39035_ (.A0(pcpi_rs1[28]),
    .A1(pcpi_rs1[27]),
    .S(mem_la_wdata[0]),
    .X(_00144_));
 sky130_fd_sc_hd__mux2_1 _39036_ (.A0(_00140_),
    .A1(_00132_),
    .S(mem_la_wdata[1]),
    .X(_00141_));
 sky130_fd_sc_hd__mux2_1 _39037_ (.A0(pcpi_rs1[27]),
    .A1(pcpi_rs1[26]),
    .S(mem_la_wdata[0]),
    .X(_00140_));
 sky130_fd_sc_hd__mux2_1 _39038_ (.A0(_00136_),
    .A1(_00128_),
    .S(mem_la_wdata[1]),
    .X(_00137_));
 sky130_fd_sc_hd__mux2_1 _39039_ (.A0(pcpi_rs1[26]),
    .A1(pcpi_rs1[25]),
    .S(mem_la_wdata[0]),
    .X(_00136_));
 sky130_fd_sc_hd__mux2_1 _39040_ (.A0(_00132_),
    .A1(_00123_),
    .S(mem_la_wdata[1]),
    .X(_00133_));
 sky130_fd_sc_hd__mux2_1 _39041_ (.A0(pcpi_rs1[25]),
    .A1(pcpi_rs1[24]),
    .S(mem_la_wdata[0]),
    .X(_00132_));
 sky130_fd_sc_hd__mux2_1 _39042_ (.A0(_00128_),
    .A1(_00117_),
    .S(mem_la_wdata[1]),
    .X(_00129_));
 sky130_fd_sc_hd__mux2_1 _39043_ (.A0(pcpi_rs1[24]),
    .A1(pcpi_rs1[23]),
    .S(mem_la_wdata[0]),
    .X(_00128_));
 sky130_fd_sc_hd__mux2_1 _39044_ (.A0(_00098_),
    .A1(_00100_),
    .S(mem_la_wdata[2]),
    .X(_00126_));
 sky130_fd_sc_hd__mux2_1 _39045_ (.A0(_00124_),
    .A1(_00097_),
    .S(mem_la_wdata[2]),
    .X(_00125_));
 sky130_fd_sc_hd__mux2_1 _39046_ (.A0(_00123_),
    .A1(_00111_),
    .S(mem_la_wdata[1]),
    .X(_00124_));
 sky130_fd_sc_hd__mux2_1 _39047_ (.A0(pcpi_rs1[23]),
    .A1(pcpi_rs1[22]),
    .S(mem_la_wdata[0]),
    .X(_00123_));
 sky130_fd_sc_hd__mux2_1 _39048_ (.A0(_00101_),
    .A1(_00094_),
    .S(mem_la_wdata[2]),
    .X(_00122_));
 sky130_fd_sc_hd__mux2_1 _39049_ (.A0(_00088_),
    .A1(_00090_),
    .S(mem_la_wdata[2]),
    .X(_00120_));
 sky130_fd_sc_hd__mux2_1 _39050_ (.A0(_00118_),
    .A1(_00087_),
    .S(mem_la_wdata[2]),
    .X(_00119_));
 sky130_fd_sc_hd__mux2_1 _39051_ (.A0(_00117_),
    .A1(_00105_),
    .S(mem_la_wdata[1]),
    .X(_00118_));
 sky130_fd_sc_hd__mux2_1 _39052_ (.A0(pcpi_rs1[22]),
    .A1(pcpi_rs1[21]),
    .S(mem_la_wdata[0]),
    .X(_00117_));
 sky130_fd_sc_hd__mux2_1 _39053_ (.A0(_00091_),
    .A1(_00084_),
    .S(mem_la_wdata[2]),
    .X(_00116_));
 sky130_fd_sc_hd__mux2_1 _39054_ (.A0(_00074_),
    .A1(_00078_),
    .S(mem_la_wdata[2]),
    .X(_00114_));
 sky130_fd_sc_hd__mux2_1 _39055_ (.A0(_00112_),
    .A1(_00071_),
    .S(mem_la_wdata[2]),
    .X(_00113_));
 sky130_fd_sc_hd__mux2_1 _39056_ (.A0(_00111_),
    .A1(_00096_),
    .S(mem_la_wdata[1]),
    .X(_00112_));
 sky130_fd_sc_hd__mux2_1 _39057_ (.A0(pcpi_rs1[21]),
    .A1(pcpi_rs1[20]),
    .S(mem_la_wdata[0]),
    .X(_00111_));
 sky130_fd_sc_hd__mux2_1 _39058_ (.A0(_00081_),
    .A1(_00067_),
    .S(mem_la_wdata[2]),
    .X(_00110_));
 sky130_fd_sc_hd__mux2_1 _39059_ (.A0(_00056_),
    .A1(_00060_),
    .S(mem_la_wdata[2]),
    .X(_00108_));
 sky130_fd_sc_hd__mux2_1 _39060_ (.A0(_00106_),
    .A1(_00053_),
    .S(mem_la_wdata[2]),
    .X(_00107_));
 sky130_fd_sc_hd__mux2_1 _39061_ (.A0(_00105_),
    .A1(_00086_),
    .S(mem_la_wdata[1]),
    .X(_00106_));
 sky130_fd_sc_hd__mux2_1 _39062_ (.A0(pcpi_rs1[20]),
    .A1(pcpi_rs1[19]),
    .S(mem_la_wdata[0]),
    .X(_00105_));
 sky130_fd_sc_hd__mux2_1 _39063_ (.A0(_00063_),
    .A1(_00049_),
    .S(mem_la_wdata[2]),
    .X(_00104_));
 sky130_fd_sc_hd__mux2_1 _39064_ (.A0(_00100_),
    .A1(_00101_),
    .S(mem_la_wdata[2]),
    .X(_00102_));
 sky130_fd_sc_hd__mux2_1 _39065_ (.A0(_00077_),
    .A1(_00079_),
    .S(mem_la_wdata[1]),
    .X(_00101_));
 sky130_fd_sc_hd__mux2_1 _39066_ (.A0(_00073_),
    .A1(_00076_),
    .S(mem_la_wdata[1]),
    .X(_00100_));
 sky130_fd_sc_hd__mux2_1 _39067_ (.A0(_00097_),
    .A1(_00098_),
    .S(mem_la_wdata[2]),
    .X(_00099_));
 sky130_fd_sc_hd__mux2_1 _39068_ (.A0(_00070_),
    .A1(_00072_),
    .S(mem_la_wdata[1]),
    .X(_00098_));
 sky130_fd_sc_hd__mux2_1 _39069_ (.A0(_00096_),
    .A1(_00069_),
    .S(mem_la_wdata[1]),
    .X(_00097_));
 sky130_fd_sc_hd__mux2_1 _39070_ (.A0(pcpi_rs1[19]),
    .A1(pcpi_rs1[18]),
    .S(mem_la_wdata[0]),
    .X(_00096_));
 sky130_fd_sc_hd__mux2_1 _39071_ (.A0(_00080_),
    .A1(_00066_),
    .S(mem_la_wdata[1]),
    .X(_00094_));
 sky130_fd_sc_hd__mux2_1 _39072_ (.A0(_00090_),
    .A1(_00091_),
    .S(mem_la_wdata[2]),
    .X(_00092_));
 sky130_fd_sc_hd__mux2_1 _39073_ (.A0(_00059_),
    .A1(_00061_),
    .S(mem_la_wdata[1]),
    .X(_00091_));
 sky130_fd_sc_hd__mux2_1 _39074_ (.A0(_00055_),
    .A1(_00058_),
    .S(mem_la_wdata[1]),
    .X(_00090_));
 sky130_fd_sc_hd__mux2_1 _39075_ (.A0(_00087_),
    .A1(_00088_),
    .S(mem_la_wdata[2]),
    .X(_00089_));
 sky130_fd_sc_hd__mux2_1 _39076_ (.A0(_00052_),
    .A1(_00054_),
    .S(mem_la_wdata[1]),
    .X(_00088_));
 sky130_fd_sc_hd__mux2_1 _39077_ (.A0(_00086_),
    .A1(_00051_),
    .S(mem_la_wdata[1]),
    .X(_00087_));
 sky130_fd_sc_hd__mux2_1 _39078_ (.A0(pcpi_rs1[18]),
    .A1(pcpi_rs1[17]),
    .S(mem_la_wdata[0]),
    .X(_00086_));
 sky130_fd_sc_hd__mux2_1 _39079_ (.A0(_00062_),
    .A1(_00048_),
    .S(mem_la_wdata[1]),
    .X(_00084_));
 sky130_fd_sc_hd__mux2_1 _39080_ (.A0(_00078_),
    .A1(_00081_),
    .S(mem_la_wdata[2]),
    .X(_00082_));
 sky130_fd_sc_hd__mux2_1 _39081_ (.A0(_00079_),
    .A1(_00080_),
    .S(mem_la_wdata[1]),
    .X(_00081_));
 sky130_fd_sc_hd__mux2_1 _39082_ (.A0(pcpi_rs1[3]),
    .A1(pcpi_rs1[2]),
    .S(mem_la_wdata[0]),
    .X(_00080_));
 sky130_fd_sc_hd__mux2_1 _39083_ (.A0(pcpi_rs1[5]),
    .A1(pcpi_rs1[4]),
    .S(mem_la_wdata[0]),
    .X(_00079_));
 sky130_fd_sc_hd__mux2_1 _39084_ (.A0(_00076_),
    .A1(_00077_),
    .S(mem_la_wdata[1]),
    .X(_00078_));
 sky130_fd_sc_hd__mux2_1 _39085_ (.A0(pcpi_rs1[7]),
    .A1(pcpi_rs1[6]),
    .S(mem_la_wdata[0]),
    .X(_00077_));
 sky130_fd_sc_hd__mux2_1 _39086_ (.A0(pcpi_rs1[9]),
    .A1(pcpi_rs1[8]),
    .S(mem_la_wdata[0]),
    .X(_00076_));
 sky130_fd_sc_hd__mux2_1 _39087_ (.A0(_00071_),
    .A1(_00074_),
    .S(mem_la_wdata[2]),
    .X(_00075_));
 sky130_fd_sc_hd__mux2_1 _39088_ (.A0(_00072_),
    .A1(_00073_),
    .S(mem_la_wdata[1]),
    .X(_00074_));
 sky130_fd_sc_hd__mux2_1 _39089_ (.A0(pcpi_rs1[11]),
    .A1(pcpi_rs1[10]),
    .S(mem_la_wdata[0]),
    .X(_00073_));
 sky130_fd_sc_hd__mux2_1 _39090_ (.A0(pcpi_rs1[13]),
    .A1(pcpi_rs1[12]),
    .S(mem_la_wdata[0]),
    .X(_00072_));
 sky130_fd_sc_hd__mux2_1 _39091_ (.A0(_00069_),
    .A1(_00070_),
    .S(mem_la_wdata[1]),
    .X(_00071_));
 sky130_fd_sc_hd__mux2_1 _39092_ (.A0(pcpi_rs1[15]),
    .A1(pcpi_rs1[14]),
    .S(mem_la_wdata[0]),
    .X(_00070_));
 sky130_fd_sc_hd__mux2_1 _39093_ (.A0(pcpi_rs1[17]),
    .A1(pcpi_rs1[16]),
    .S(mem_la_wdata[0]),
    .X(_00069_));
 sky130_fd_sc_hd__mux2_1 _39094_ (.A0(pcpi_rs1[1]),
    .A1(pcpi_rs1[0]),
    .S(mem_la_wdata[0]),
    .X(_00066_));
 sky130_fd_sc_hd__mux2_1 _39095_ (.A0(_00060_),
    .A1(_00063_),
    .S(mem_la_wdata[2]),
    .X(_00064_));
 sky130_fd_sc_hd__mux2_1 _39096_ (.A0(_00061_),
    .A1(_00062_),
    .S(mem_la_wdata[1]),
    .X(_00063_));
 sky130_fd_sc_hd__mux2_1 _39097_ (.A0(pcpi_rs1[2]),
    .A1(pcpi_rs1[1]),
    .S(mem_la_wdata[0]),
    .X(_00062_));
 sky130_fd_sc_hd__mux2_1 _39098_ (.A0(pcpi_rs1[4]),
    .A1(pcpi_rs1[3]),
    .S(mem_la_wdata[0]),
    .X(_00061_));
 sky130_fd_sc_hd__mux2_1 _39099_ (.A0(_00058_),
    .A1(_00059_),
    .S(mem_la_wdata[1]),
    .X(_00060_));
 sky130_fd_sc_hd__mux2_1 _39100_ (.A0(pcpi_rs1[6]),
    .A1(pcpi_rs1[5]),
    .S(mem_la_wdata[0]),
    .X(_00059_));
 sky130_fd_sc_hd__mux2_1 _39101_ (.A0(pcpi_rs1[8]),
    .A1(pcpi_rs1[7]),
    .S(mem_la_wdata[0]),
    .X(_00058_));
 sky130_fd_sc_hd__mux2_1 _39102_ (.A0(_00053_),
    .A1(_00056_),
    .S(mem_la_wdata[2]),
    .X(_00057_));
 sky130_fd_sc_hd__mux2_1 _39103_ (.A0(_00054_),
    .A1(_00055_),
    .S(mem_la_wdata[1]),
    .X(_00056_));
 sky130_fd_sc_hd__mux2_1 _39104_ (.A0(pcpi_rs1[10]),
    .A1(pcpi_rs1[9]),
    .S(mem_la_wdata[0]),
    .X(_00055_));
 sky130_fd_sc_hd__mux2_1 _39105_ (.A0(pcpi_rs1[12]),
    .A1(pcpi_rs1[11]),
    .S(mem_la_wdata[0]),
    .X(_00054_));
 sky130_fd_sc_hd__mux2_1 _39106_ (.A0(_00051_),
    .A1(_00052_),
    .S(mem_la_wdata[1]),
    .X(_00053_));
 sky130_fd_sc_hd__mux2_1 _39107_ (.A0(pcpi_rs1[14]),
    .A1(pcpi_rs1[13]),
    .S(mem_la_wdata[0]),
    .X(_00052_));
 sky130_fd_sc_hd__mux2_1 _39108_ (.A0(pcpi_rs1[16]),
    .A1(pcpi_rs1[15]),
    .S(mem_la_wdata[0]),
    .X(_00051_));
 sky130_fd_sc_hd__mux2_1 _39109_ (.A0(_02408_),
    .A1(pcpi_rs2[31]),
    .S(instr_sub),
    .X(_02409_));
 sky130_fd_sc_hd__mux2_1 _39110_ (.A0(_02406_),
    .A1(_02405_),
    .S(instr_sub),
    .X(_02407_));
 sky130_fd_sc_hd__mux2_1 _39111_ (.A0(_02403_),
    .A1(_02402_),
    .S(instr_sub),
    .X(_02404_));
 sky130_fd_sc_hd__mux2_1 _39112_ (.A0(_02400_),
    .A1(_02399_),
    .S(instr_sub),
    .X(_02401_));
 sky130_fd_sc_hd__mux2_1 _39113_ (.A0(_02397_),
    .A1(_02396_),
    .S(instr_sub),
    .X(_02398_));
 sky130_fd_sc_hd__mux2_1 _39114_ (.A0(_02394_),
    .A1(_02393_),
    .S(instr_sub),
    .X(_02395_));
 sky130_fd_sc_hd__mux2_1 _39115_ (.A0(_02391_),
    .A1(_02390_),
    .S(instr_sub),
    .X(_02392_));
 sky130_fd_sc_hd__mux2_1 _39116_ (.A0(_02388_),
    .A1(_02387_),
    .S(instr_sub),
    .X(_02389_));
 sky130_fd_sc_hd__mux2_1 _39117_ (.A0(_02385_),
    .A1(_02384_),
    .S(instr_sub),
    .X(_02386_));
 sky130_fd_sc_hd__mux2_1 _39118_ (.A0(_02382_),
    .A1(_02381_),
    .S(instr_sub),
    .X(_02383_));
 sky130_fd_sc_hd__mux2_1 _39119_ (.A0(_02379_),
    .A1(_02378_),
    .S(instr_sub),
    .X(_02380_));
 sky130_fd_sc_hd__mux2_1 _39120_ (.A0(_02376_),
    .A1(_02375_),
    .S(instr_sub),
    .X(_02377_));
 sky130_fd_sc_hd__mux2_1 _39121_ (.A0(_02373_),
    .A1(_02372_),
    .S(instr_sub),
    .X(_02374_));
 sky130_fd_sc_hd__mux2_1 _39122_ (.A0(_02370_),
    .A1(_02369_),
    .S(instr_sub),
    .X(_02371_));
 sky130_fd_sc_hd__mux2_1 _39123_ (.A0(_02367_),
    .A1(_02366_),
    .S(instr_sub),
    .X(_02368_));
 sky130_fd_sc_hd__mux2_1 _39124_ (.A0(_02364_),
    .A1(_02363_),
    .S(instr_sub),
    .X(_02365_));
 sky130_fd_sc_hd__mux2_1 _39125_ (.A0(_02361_),
    .A1(_02360_),
    .S(instr_sub),
    .X(_02362_));
 sky130_fd_sc_hd__mux2_1 _39126_ (.A0(_02358_),
    .A1(_02357_),
    .S(instr_sub),
    .X(_02359_));
 sky130_fd_sc_hd__mux2_1 _39127_ (.A0(_02355_),
    .A1(_02354_),
    .S(instr_sub),
    .X(_02356_));
 sky130_fd_sc_hd__mux2_1 _39128_ (.A0(_02352_),
    .A1(_02351_),
    .S(instr_sub),
    .X(_02353_));
 sky130_fd_sc_hd__mux2_1 _39129_ (.A0(_02349_),
    .A1(_02348_),
    .S(instr_sub),
    .X(_02350_));
 sky130_fd_sc_hd__mux2_1 _39130_ (.A0(_02346_),
    .A1(_02345_),
    .S(instr_sub),
    .X(_02347_));
 sky130_fd_sc_hd__mux2_1 _39131_ (.A0(_02343_),
    .A1(_02342_),
    .S(instr_sub),
    .X(_02344_));
 sky130_fd_sc_hd__mux2_1 _39132_ (.A0(_02340_),
    .A1(_02339_),
    .S(instr_sub),
    .X(_02341_));
 sky130_fd_sc_hd__mux2_1 _39133_ (.A0(_02337_),
    .A1(_02336_),
    .S(instr_sub),
    .X(_02338_));
 sky130_fd_sc_hd__mux2_1 _39134_ (.A0(_02334_),
    .A1(_02333_),
    .S(instr_sub),
    .X(_02335_));
 sky130_fd_sc_hd__mux2_1 _39135_ (.A0(_02331_),
    .A1(_02330_),
    .S(instr_sub),
    .X(_02332_));
 sky130_fd_sc_hd__mux2_1 _39136_ (.A0(_02328_),
    .A1(_02327_),
    .S(instr_sub),
    .X(_02329_));
 sky130_fd_sc_hd__mux2_1 _39137_ (.A0(_02325_),
    .A1(_02324_),
    .S(instr_sub),
    .X(_02326_));
 sky130_fd_sc_hd__mux2_1 _39138_ (.A0(_02322_),
    .A1(_02321_),
    .S(instr_sub),
    .X(_02323_));
 sky130_fd_sc_hd__mux2_1 _39139_ (.A0(_02319_),
    .A1(_02318_),
    .S(instr_sub),
    .X(_02320_));
 sky130_fd_sc_hd__mux2_1 _39140_ (.A0(_02313_),
    .A1(_02314_),
    .S(_00306_),
    .X(_02315_));
 sky130_fd_sc_hd__mux2_1 _39141_ (.A0(_02311_),
    .A1(_02315_),
    .S(_00303_),
    .X(_02316_));
 sky130_fd_sc_hd__mux2_1 _39142_ (.A0(_02311_),
    .A1(_02312_),
    .S(_00305_),
    .X(_02313_));
 sky130_fd_sc_hd__mux2_1 _39143_ (.A0(_02307_),
    .A1(_02308_),
    .S(\irq_state[1] ),
    .X(_02309_));
 sky130_fd_sc_hd__mux2_1 _39144_ (.A0(_02309_),
    .A1(_02307_),
    .S(_02217_),
    .X(_02310_));
 sky130_fd_sc_hd__mux2_1 _39145_ (.A0(_02302_),
    .A1(\irq_pending[0] ),
    .S(_01208_),
    .X(_02303_));
 sky130_fd_sc_hd__mux2_1 _39146_ (.A0(\reg_out[0] ),
    .A1(\alu_out_q[0] ),
    .S(latched_stalu),
    .X(_02070_));
 sky130_fd_sc_hd__mux2_1 _39147_ (.A0(_02063_),
    .A1(_00343_),
    .S(is_beq_bne_blt_bge_bltu_bgeu),
    .X(_02064_));
 sky130_fd_sc_hd__mux2_1 _39148_ (.A0(_02056_),
    .A1(_02055_),
    .S(_01714_),
    .X(_02057_));
 sky130_fd_sc_hd__mux2_1 _39149_ (.A0(_02058_),
    .A1(_02057_),
    .S(_01717_),
    .X(_02059_));
 sky130_fd_sc_hd__mux2_1 _39150_ (.A0(\pcpi_mul.rd[31] ),
    .A1(\pcpi_mul.rd[63] ),
    .S(\pcpi_mul.shift_out ),
    .X(_02054_));
 sky130_fd_sc_hd__mux2_1 _39151_ (.A0(_01908_),
    .A1(_02052_),
    .S(_01816_),
    .X(_02053_));
 sky130_fd_sc_hd__mux2_1 _39152_ (.A0(_02047_),
    .A1(_02046_),
    .S(_01714_),
    .X(_02048_));
 sky130_fd_sc_hd__mux2_1 _39153_ (.A0(_02049_),
    .A1(_02048_),
    .S(_01717_),
    .X(_02050_));
 sky130_fd_sc_hd__mux2_1 _39154_ (.A0(\pcpi_mul.rd[30] ),
    .A1(\pcpi_mul.rd[62] ),
    .S(\pcpi_mul.shift_out ),
    .X(_02045_));
 sky130_fd_sc_hd__mux2_1 _39155_ (.A0(_01908_),
    .A1(_02043_),
    .S(_01816_),
    .X(_02044_));
 sky130_fd_sc_hd__mux2_1 _39156_ (.A0(_02038_),
    .A1(_02037_),
    .S(_01714_),
    .X(_02039_));
 sky130_fd_sc_hd__mux2_1 _39157_ (.A0(_02040_),
    .A1(_02039_),
    .S(_01717_),
    .X(_02041_));
 sky130_fd_sc_hd__mux2_1 _39158_ (.A0(\pcpi_mul.rd[29] ),
    .A1(\pcpi_mul.rd[61] ),
    .S(\pcpi_mul.shift_out ),
    .X(_02036_));
 sky130_fd_sc_hd__mux2_1 _39159_ (.A0(_01908_),
    .A1(_02034_),
    .S(_01816_),
    .X(_02035_));
 sky130_fd_sc_hd__mux2_1 _39160_ (.A0(_02029_),
    .A1(_02028_),
    .S(_01714_),
    .X(_02030_));
 sky130_fd_sc_hd__mux2_1 _39161_ (.A0(_02031_),
    .A1(_02030_),
    .S(_01717_),
    .X(_02032_));
 sky130_fd_sc_hd__mux2_1 _39162_ (.A0(\pcpi_mul.rd[28] ),
    .A1(\pcpi_mul.rd[60] ),
    .S(\pcpi_mul.shift_out ),
    .X(_02027_));
 sky130_fd_sc_hd__mux2_1 _39163_ (.A0(_01908_),
    .A1(_02025_),
    .S(_01816_),
    .X(_02026_));
 sky130_fd_sc_hd__mux2_1 _39164_ (.A0(_02020_),
    .A1(_02019_),
    .S(_01714_),
    .X(_02021_));
 sky130_fd_sc_hd__mux2_1 _39165_ (.A0(_02022_),
    .A1(_02021_),
    .S(_01717_),
    .X(_02023_));
 sky130_fd_sc_hd__mux2_1 _39166_ (.A0(\pcpi_mul.rd[27] ),
    .A1(\pcpi_mul.rd[59] ),
    .S(\pcpi_mul.shift_out ),
    .X(_02018_));
 sky130_fd_sc_hd__mux2_1 _39167_ (.A0(_01908_),
    .A1(_02016_),
    .S(_01816_),
    .X(_02017_));
 sky130_fd_sc_hd__mux2_1 _39168_ (.A0(_02011_),
    .A1(_02010_),
    .S(_01714_),
    .X(_02012_));
 sky130_fd_sc_hd__mux2_1 _39169_ (.A0(_02013_),
    .A1(_02012_),
    .S(_01717_),
    .X(_02014_));
 sky130_fd_sc_hd__mux2_1 _39170_ (.A0(\pcpi_mul.rd[26] ),
    .A1(\pcpi_mul.rd[58] ),
    .S(\pcpi_mul.shift_out ),
    .X(_02009_));
 sky130_fd_sc_hd__mux2_1 _39171_ (.A0(_01908_),
    .A1(_02007_),
    .S(_01816_),
    .X(_02008_));
 sky130_fd_sc_hd__mux2_1 _39172_ (.A0(_02002_),
    .A1(_02001_),
    .S(_01714_),
    .X(_02003_));
 sky130_fd_sc_hd__mux2_1 _39173_ (.A0(_02004_),
    .A1(_02003_),
    .S(_01717_),
    .X(_02005_));
 sky130_fd_sc_hd__mux2_1 _39174_ (.A0(\pcpi_mul.rd[25] ),
    .A1(\pcpi_mul.rd[57] ),
    .S(\pcpi_mul.shift_out ),
    .X(_02000_));
 sky130_fd_sc_hd__mux2_1 _39175_ (.A0(_01908_),
    .A1(_01998_),
    .S(_01816_),
    .X(_01999_));
 sky130_fd_sc_hd__mux2_1 _39176_ (.A0(_01993_),
    .A1(_01992_),
    .S(_01714_),
    .X(_01994_));
 sky130_fd_sc_hd__mux2_1 _39177_ (.A0(_01995_),
    .A1(_01994_),
    .S(_01717_),
    .X(_01996_));
 sky130_fd_sc_hd__mux2_1 _39178_ (.A0(\pcpi_mul.rd[24] ),
    .A1(\pcpi_mul.rd[56] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01991_));
 sky130_fd_sc_hd__mux2_1 _39179_ (.A0(_01908_),
    .A1(_01989_),
    .S(_01816_),
    .X(_01990_));
 sky130_fd_sc_hd__mux2_1 _39180_ (.A0(_01984_),
    .A1(_01983_),
    .S(_01714_),
    .X(_01985_));
 sky130_fd_sc_hd__mux2_1 _39181_ (.A0(_01986_),
    .A1(_01985_),
    .S(_01717_),
    .X(_01987_));
 sky130_fd_sc_hd__mux2_1 _39182_ (.A0(\pcpi_mul.rd[23] ),
    .A1(\pcpi_mul.rd[55] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01982_));
 sky130_fd_sc_hd__mux2_1 _39183_ (.A0(_01908_),
    .A1(_01980_),
    .S(_01816_),
    .X(_01981_));
 sky130_fd_sc_hd__mux2_1 _39184_ (.A0(_01975_),
    .A1(_01974_),
    .S(_01714_),
    .X(_01976_));
 sky130_fd_sc_hd__mux2_1 _39185_ (.A0(_01977_),
    .A1(_01976_),
    .S(_01717_),
    .X(_01978_));
 sky130_fd_sc_hd__mux2_1 _39186_ (.A0(\pcpi_mul.rd[22] ),
    .A1(\pcpi_mul.rd[54] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01973_));
 sky130_fd_sc_hd__mux2_1 _39187_ (.A0(_01908_),
    .A1(_01971_),
    .S(_01816_),
    .X(_01972_));
 sky130_fd_sc_hd__mux2_1 _39188_ (.A0(_01966_),
    .A1(_01965_),
    .S(_01714_),
    .X(_01967_));
 sky130_fd_sc_hd__mux2_1 _39189_ (.A0(_01968_),
    .A1(_01967_),
    .S(_01717_),
    .X(_01969_));
 sky130_fd_sc_hd__mux2_1 _39190_ (.A0(\pcpi_mul.rd[21] ),
    .A1(\pcpi_mul.rd[53] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01964_));
 sky130_fd_sc_hd__mux2_1 _39191_ (.A0(_01908_),
    .A1(_01962_),
    .S(_01816_),
    .X(_01963_));
 sky130_fd_sc_hd__mux2_1 _39192_ (.A0(_01957_),
    .A1(_01956_),
    .S(_01714_),
    .X(_01958_));
 sky130_fd_sc_hd__mux2_1 _39193_ (.A0(_01959_),
    .A1(_01958_),
    .S(_01717_),
    .X(_01960_));
 sky130_fd_sc_hd__mux2_1 _39194_ (.A0(\pcpi_mul.rd[20] ),
    .A1(\pcpi_mul.rd[52] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01955_));
 sky130_fd_sc_hd__mux2_1 _39195_ (.A0(_01908_),
    .A1(_01953_),
    .S(_01816_),
    .X(_01954_));
 sky130_fd_sc_hd__mux2_1 _39196_ (.A0(_01948_),
    .A1(_01947_),
    .S(_01714_),
    .X(_01949_));
 sky130_fd_sc_hd__mux2_1 _39197_ (.A0(_01950_),
    .A1(_01949_),
    .S(_01717_),
    .X(_01951_));
 sky130_fd_sc_hd__mux2_1 _39198_ (.A0(\pcpi_mul.rd[19] ),
    .A1(\pcpi_mul.rd[51] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01946_));
 sky130_fd_sc_hd__mux2_1 _39199_ (.A0(_01908_),
    .A1(_01944_),
    .S(_01816_),
    .X(_01945_));
 sky130_fd_sc_hd__mux2_1 _39200_ (.A0(_01939_),
    .A1(_01938_),
    .S(_01714_),
    .X(_01940_));
 sky130_fd_sc_hd__mux2_1 _39201_ (.A0(_01941_),
    .A1(_01940_),
    .S(_01717_),
    .X(_01942_));
 sky130_fd_sc_hd__mux2_1 _39202_ (.A0(\pcpi_mul.rd[18] ),
    .A1(\pcpi_mul.rd[50] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01937_));
 sky130_fd_sc_hd__mux2_1 _39203_ (.A0(_01908_),
    .A1(_01935_),
    .S(_01816_),
    .X(_01936_));
 sky130_fd_sc_hd__mux2_1 _39204_ (.A0(_01930_),
    .A1(_01929_),
    .S(_01714_),
    .X(_01931_));
 sky130_fd_sc_hd__mux2_1 _39205_ (.A0(_01932_),
    .A1(_01931_),
    .S(_01717_),
    .X(_01933_));
 sky130_fd_sc_hd__mux2_1 _39206_ (.A0(\pcpi_mul.rd[17] ),
    .A1(\pcpi_mul.rd[49] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01928_));
 sky130_fd_sc_hd__mux2_1 _39207_ (.A0(_01908_),
    .A1(_01926_),
    .S(_01816_),
    .X(_01927_));
 sky130_fd_sc_hd__mux2_1 _39208_ (.A0(_01921_),
    .A1(_01920_),
    .S(_01714_),
    .X(_01922_));
 sky130_fd_sc_hd__mux2_1 _39209_ (.A0(_01923_),
    .A1(_01922_),
    .S(_01717_),
    .X(_01924_));
 sky130_fd_sc_hd__mux2_1 _39210_ (.A0(\pcpi_mul.rd[16] ),
    .A1(\pcpi_mul.rd[48] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01919_));
 sky130_fd_sc_hd__mux2_1 _39211_ (.A0(_01908_),
    .A1(_01917_),
    .S(_01816_),
    .X(_01918_));
 sky130_fd_sc_hd__mux2_1 _39212_ (.A0(_01912_),
    .A1(_01911_),
    .S(_01714_),
    .X(_01913_));
 sky130_fd_sc_hd__mux2_1 _39213_ (.A0(_01914_),
    .A1(_01913_),
    .S(_01717_),
    .X(_01915_));
 sky130_fd_sc_hd__mux2_1 _39214_ (.A0(\pcpi_mul.rd[15] ),
    .A1(\pcpi_mul.rd[47] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01910_));
 sky130_fd_sc_hd__mux2_1 _39215_ (.A0(_01908_),
    .A1(_01907_),
    .S(_01816_),
    .X(_01909_));
 sky130_fd_sc_hd__mux2_1 _39216_ (.A0(_01906_),
    .A1(_01904_),
    .S(_01683_),
    .X(_01907_));
 sky130_fd_sc_hd__mux2_1 _39217_ (.A0(mem_rdata[15]),
    .A1(mem_rdata[31]),
    .S(pcpi_rs1[1]),
    .X(_01905_));
 sky130_fd_sc_hd__mux2_1 _39218_ (.A0(_01899_),
    .A1(_01898_),
    .S(_01714_),
    .X(_01900_));
 sky130_fd_sc_hd__mux2_1 _39219_ (.A0(_01901_),
    .A1(_01900_),
    .S(_01717_),
    .X(_01902_));
 sky130_fd_sc_hd__mux2_1 _39220_ (.A0(\pcpi_mul.rd[14] ),
    .A1(\pcpi_mul.rd[46] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01897_));
 sky130_fd_sc_hd__mux2_1 _39221_ (.A0(_01895_),
    .A1(_01894_),
    .S(_01816_),
    .X(_01896_));
 sky130_fd_sc_hd__mux2_1 _39222_ (.A0(_01893_),
    .A1(_01891_),
    .S(_01683_),
    .X(_01894_));
 sky130_fd_sc_hd__mux2_1 _39223_ (.A0(mem_rdata[14]),
    .A1(mem_rdata[30]),
    .S(pcpi_rs1[1]),
    .X(_01892_));
 sky130_fd_sc_hd__mux2_1 _39224_ (.A0(_01886_),
    .A1(_01885_),
    .S(_01714_),
    .X(_01887_));
 sky130_fd_sc_hd__mux2_1 _39225_ (.A0(_01888_),
    .A1(_01887_),
    .S(_01717_),
    .X(_01889_));
 sky130_fd_sc_hd__mux2_1 _39226_ (.A0(\pcpi_mul.rd[13] ),
    .A1(\pcpi_mul.rd[45] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01884_));
 sky130_fd_sc_hd__mux2_1 _39227_ (.A0(_01882_),
    .A1(_01881_),
    .S(_01816_),
    .X(_01883_));
 sky130_fd_sc_hd__mux2_1 _39228_ (.A0(_01880_),
    .A1(_01878_),
    .S(_01683_),
    .X(_01881_));
 sky130_fd_sc_hd__mux2_1 _39229_ (.A0(mem_rdata[13]),
    .A1(mem_rdata[29]),
    .S(pcpi_rs1[1]),
    .X(_01879_));
 sky130_fd_sc_hd__mux2_1 _39230_ (.A0(_01873_),
    .A1(_01872_),
    .S(_01714_),
    .X(_01874_));
 sky130_fd_sc_hd__mux2_1 _39231_ (.A0(_01875_),
    .A1(_01874_),
    .S(_01717_),
    .X(_01876_));
 sky130_fd_sc_hd__mux2_1 _39232_ (.A0(\pcpi_mul.rd[12] ),
    .A1(\pcpi_mul.rd[44] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01871_));
 sky130_fd_sc_hd__mux2_1 _39233_ (.A0(_01869_),
    .A1(_01868_),
    .S(_01816_),
    .X(_01870_));
 sky130_fd_sc_hd__mux2_1 _39234_ (.A0(_01867_),
    .A1(_01865_),
    .S(_01683_),
    .X(_01868_));
 sky130_fd_sc_hd__mux2_1 _39235_ (.A0(mem_rdata[12]),
    .A1(mem_rdata[28]),
    .S(pcpi_rs1[1]),
    .X(_01866_));
 sky130_fd_sc_hd__mux2_1 _39236_ (.A0(_01860_),
    .A1(_01859_),
    .S(_01714_),
    .X(_01861_));
 sky130_fd_sc_hd__mux2_1 _39237_ (.A0(_01862_),
    .A1(_01861_),
    .S(_01717_),
    .X(_01863_));
 sky130_fd_sc_hd__mux2_1 _39238_ (.A0(\pcpi_mul.rd[11] ),
    .A1(\pcpi_mul.rd[43] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01858_));
 sky130_fd_sc_hd__mux2_1 _39239_ (.A0(_01856_),
    .A1(_01855_),
    .S(_01816_),
    .X(_01857_));
 sky130_fd_sc_hd__mux2_1 _39240_ (.A0(_01854_),
    .A1(_01852_),
    .S(_01683_),
    .X(_01855_));
 sky130_fd_sc_hd__mux2_1 _39241_ (.A0(mem_rdata[11]),
    .A1(mem_rdata[27]),
    .S(pcpi_rs1[1]),
    .X(_01853_));
 sky130_fd_sc_hd__mux2_1 _39242_ (.A0(_01847_),
    .A1(_01846_),
    .S(_01714_),
    .X(_01848_));
 sky130_fd_sc_hd__mux2_1 _39243_ (.A0(_01849_),
    .A1(_01848_),
    .S(_01717_),
    .X(_01850_));
 sky130_fd_sc_hd__mux2_1 _39244_ (.A0(\pcpi_mul.rd[10] ),
    .A1(\pcpi_mul.rd[42] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01845_));
 sky130_fd_sc_hd__mux2_1 _39245_ (.A0(_01843_),
    .A1(_01842_),
    .S(_01816_),
    .X(_01844_));
 sky130_fd_sc_hd__mux2_1 _39246_ (.A0(_01841_),
    .A1(_01839_),
    .S(_01683_),
    .X(_01842_));
 sky130_fd_sc_hd__mux2_1 _39247_ (.A0(mem_rdata[10]),
    .A1(mem_rdata[26]),
    .S(pcpi_rs1[1]),
    .X(_01840_));
 sky130_fd_sc_hd__mux2_1 _39248_ (.A0(_01834_),
    .A1(_01833_),
    .S(_01714_),
    .X(_01835_));
 sky130_fd_sc_hd__mux2_1 _39249_ (.A0(_01836_),
    .A1(_01835_),
    .S(_01717_),
    .X(_01837_));
 sky130_fd_sc_hd__mux2_1 _39250_ (.A0(\pcpi_mul.rd[9] ),
    .A1(\pcpi_mul.rd[41] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01832_));
 sky130_fd_sc_hd__mux2_1 _39251_ (.A0(_01830_),
    .A1(_01829_),
    .S(_01816_),
    .X(_01831_));
 sky130_fd_sc_hd__mux2_1 _39252_ (.A0(_01828_),
    .A1(_01826_),
    .S(_01683_),
    .X(_01829_));
 sky130_fd_sc_hd__mux2_1 _39253_ (.A0(mem_rdata[9]),
    .A1(mem_rdata[25]),
    .S(pcpi_rs1[1]),
    .X(_01827_));
 sky130_fd_sc_hd__mux2_1 _39254_ (.A0(_01821_),
    .A1(_01820_),
    .S(_01714_),
    .X(_01822_));
 sky130_fd_sc_hd__mux2_1 _39255_ (.A0(_01823_),
    .A1(_01822_),
    .S(_01717_),
    .X(_01824_));
 sky130_fd_sc_hd__mux2_1 _39256_ (.A0(\pcpi_mul.rd[8] ),
    .A1(\pcpi_mul.rd[40] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01819_));
 sky130_fd_sc_hd__mux2_1 _39257_ (.A0(_01817_),
    .A1(_01815_),
    .S(_01816_),
    .X(_01818_));
 sky130_fd_sc_hd__mux2_1 _39258_ (.A0(_01814_),
    .A1(_01812_),
    .S(_01683_),
    .X(_01815_));
 sky130_fd_sc_hd__mux2_1 _39259_ (.A0(mem_rdata[8]),
    .A1(mem_rdata[24]),
    .S(pcpi_rs1[1]),
    .X(_01813_));
 sky130_fd_sc_hd__mux2_1 _39260_ (.A0(_01807_),
    .A1(_01806_),
    .S(_01714_),
    .X(_01808_));
 sky130_fd_sc_hd__mux2_1 _39261_ (.A0(_01809_),
    .A1(_01808_),
    .S(_01717_),
    .X(_01810_));
 sky130_fd_sc_hd__mux2_1 _39262_ (.A0(\pcpi_mul.rd[7] ),
    .A1(\pcpi_mul.rd[39] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01805_));
 sky130_fd_sc_hd__mux2_1 _39263_ (.A0(_01803_),
    .A1(_01799_),
    .S(_01683_),
    .X(_01804_));
 sky130_fd_sc_hd__mux2_1 _39264_ (.A0(mem_rdata[7]),
    .A1(mem_rdata[23]),
    .S(pcpi_rs1[1]),
    .X(_01802_));
 sky130_fd_sc_hd__mux2_1 _39265_ (.A0(_01800_),
    .A1(_01799_),
    .S(_00304_),
    .X(_01801_));
 sky130_fd_sc_hd__mux2_1 _39266_ (.A0(_01794_),
    .A1(_01793_),
    .S(_01714_),
    .X(_01795_));
 sky130_fd_sc_hd__mux2_1 _39267_ (.A0(_01796_),
    .A1(_01795_),
    .S(_01717_),
    .X(_01797_));
 sky130_fd_sc_hd__mux2_1 _39268_ (.A0(\pcpi_mul.rd[6] ),
    .A1(\pcpi_mul.rd[38] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01792_));
 sky130_fd_sc_hd__mux2_1 _39269_ (.A0(_01790_),
    .A1(_01786_),
    .S(_01683_),
    .X(_01791_));
 sky130_fd_sc_hd__mux2_1 _39270_ (.A0(mem_rdata[6]),
    .A1(mem_rdata[22]),
    .S(pcpi_rs1[1]),
    .X(_01789_));
 sky130_fd_sc_hd__mux2_1 _39271_ (.A0(_01787_),
    .A1(_01786_),
    .S(_00304_),
    .X(_01788_));
 sky130_fd_sc_hd__mux2_1 _39272_ (.A0(_01781_),
    .A1(_01780_),
    .S(_01714_),
    .X(_01782_));
 sky130_fd_sc_hd__mux2_1 _39273_ (.A0(_01783_),
    .A1(_01782_),
    .S(_01717_),
    .X(_01784_));
 sky130_fd_sc_hd__mux2_1 _39274_ (.A0(\pcpi_mul.rd[5] ),
    .A1(\pcpi_mul.rd[37] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01779_));
 sky130_fd_sc_hd__mux2_1 _39275_ (.A0(_01777_),
    .A1(_01773_),
    .S(_01683_),
    .X(_01778_));
 sky130_fd_sc_hd__mux2_1 _39276_ (.A0(mem_rdata[5]),
    .A1(mem_rdata[21]),
    .S(pcpi_rs1[1]),
    .X(_01776_));
 sky130_fd_sc_hd__mux2_1 _39277_ (.A0(_01774_),
    .A1(_01773_),
    .S(_00304_),
    .X(_01775_));
 sky130_fd_sc_hd__mux2_1 _39278_ (.A0(_01768_),
    .A1(_01767_),
    .S(_01714_),
    .X(_01769_));
 sky130_fd_sc_hd__mux2_1 _39279_ (.A0(_01770_),
    .A1(_01769_),
    .S(_01717_),
    .X(_01771_));
 sky130_fd_sc_hd__mux2_1 _39280_ (.A0(\pcpi_mul.rd[4] ),
    .A1(\pcpi_mul.rd[36] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01766_));
 sky130_fd_sc_hd__mux2_1 _39281_ (.A0(_01764_),
    .A1(_01760_),
    .S(_01683_),
    .X(_01765_));
 sky130_fd_sc_hd__mux2_1 _39282_ (.A0(mem_rdata[4]),
    .A1(mem_rdata[20]),
    .S(pcpi_rs1[1]),
    .X(_01763_));
 sky130_fd_sc_hd__mux2_1 _39283_ (.A0(_01761_),
    .A1(_01760_),
    .S(_00304_),
    .X(_01762_));
 sky130_fd_sc_hd__mux2_1 _39284_ (.A0(_01755_),
    .A1(_01754_),
    .S(_01714_),
    .X(_01756_));
 sky130_fd_sc_hd__mux2_1 _39285_ (.A0(_01757_),
    .A1(_01756_),
    .S(_01717_),
    .X(_01758_));
 sky130_fd_sc_hd__mux2_1 _39286_ (.A0(\pcpi_mul.rd[3] ),
    .A1(\pcpi_mul.rd[35] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01753_));
 sky130_fd_sc_hd__mux2_1 _39287_ (.A0(_01751_),
    .A1(_01747_),
    .S(_01683_),
    .X(_01752_));
 sky130_fd_sc_hd__mux2_1 _39288_ (.A0(mem_rdata[3]),
    .A1(mem_rdata[19]),
    .S(pcpi_rs1[1]),
    .X(_01750_));
 sky130_fd_sc_hd__mux2_1 _39289_ (.A0(_01748_),
    .A1(_01747_),
    .S(_00304_),
    .X(_01749_));
 sky130_fd_sc_hd__mux2_1 _39290_ (.A0(_01742_),
    .A1(_01741_),
    .S(_01714_),
    .X(_01743_));
 sky130_fd_sc_hd__mux2_1 _39291_ (.A0(_01744_),
    .A1(_01743_),
    .S(_01717_),
    .X(_01745_));
 sky130_fd_sc_hd__mux2_1 _39292_ (.A0(\pcpi_mul.rd[2] ),
    .A1(\pcpi_mul.rd[34] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01740_));
 sky130_fd_sc_hd__mux2_1 _39293_ (.A0(_01738_),
    .A1(_01734_),
    .S(_01683_),
    .X(_01739_));
 sky130_fd_sc_hd__mux2_1 _39294_ (.A0(mem_rdata[2]),
    .A1(mem_rdata[18]),
    .S(pcpi_rs1[1]),
    .X(_01737_));
 sky130_fd_sc_hd__mux2_1 _39295_ (.A0(_01735_),
    .A1(_01734_),
    .S(_00304_),
    .X(_01736_));
 sky130_fd_sc_hd__mux2_1 _39296_ (.A0(_01729_),
    .A1(_01728_),
    .S(_01714_),
    .X(_01730_));
 sky130_fd_sc_hd__mux2_1 _39297_ (.A0(_01731_),
    .A1(_01730_),
    .S(_01717_),
    .X(_01732_));
 sky130_fd_sc_hd__mux2_1 _39298_ (.A0(\pcpi_mul.rd[1] ),
    .A1(\pcpi_mul.rd[33] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01727_));
 sky130_fd_sc_hd__mux2_1 _39299_ (.A0(_01725_),
    .A1(_01721_),
    .S(_01683_),
    .X(_01726_));
 sky130_fd_sc_hd__mux2_1 _39300_ (.A0(mem_rdata[1]),
    .A1(mem_rdata[17]),
    .S(pcpi_rs1[1]),
    .X(_01724_));
 sky130_fd_sc_hd__mux2_1 _39301_ (.A0(_01722_),
    .A1(_01721_),
    .S(_00304_),
    .X(_01723_));
 sky130_fd_sc_hd__mux2_1 _39302_ (.A0(_01715_),
    .A1(_02559_),
    .S(_01714_),
    .X(_01716_));
 sky130_fd_sc_hd__mux2_1 _39303_ (.A0(_01718_),
    .A1(_01716_),
    .S(_01717_),
    .X(_01719_));
 sky130_fd_sc_hd__mux2_1 _39304_ (.A0(\pcpi_mul.rd[0] ),
    .A1(\pcpi_mul.rd[32] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01713_));
 sky130_fd_sc_hd__mux2_1 _39305_ (.A0(_01711_),
    .A1(_01707_),
    .S(_01683_),
    .X(_01712_));
 sky130_fd_sc_hd__mux2_1 _39306_ (.A0(mem_rdata[0]),
    .A1(mem_rdata[16]),
    .S(pcpi_rs1[1]),
    .X(_01710_));
 sky130_fd_sc_hd__mux2_1 _39307_ (.A0(_01708_),
    .A1(_01707_),
    .S(_00304_),
    .X(_01709_));
 sky130_fd_sc_hd__mux2_1 _39308_ (.A0(_01701_),
    .A1(_01696_),
    .S(_00311_),
    .X(_01702_));
 sky130_fd_sc_hd__mux2_1 _39309_ (.A0(_01702_),
    .A1(_01696_),
    .S(\pcpi_mul.active[1] ),
    .X(_01703_));
 sky130_fd_sc_hd__mux2_1 _39310_ (.A0(_01696_),
    .A1(_01703_),
    .S(_00310_),
    .X(_01704_));
 sky130_fd_sc_hd__mux2_1 _39311_ (.A0(_01693_),
    .A1(mem_wstrb[3]),
    .S(_00316_),
    .X(_01694_));
 sky130_fd_sc_hd__mux2_1 _39312_ (.A0(_01690_),
    .A1(mem_wstrb[2]),
    .S(_00316_),
    .X(_01691_));
 sky130_fd_sc_hd__mux2_1 _39313_ (.A0(_01687_),
    .A1(mem_wstrb[1]),
    .S(_00316_),
    .X(_01688_));
 sky130_fd_sc_hd__mux2_1 _39314_ (.A0(_01684_),
    .A1(mem_wstrb[0]),
    .S(_00316_),
    .X(_01685_));
 sky130_fd_sc_hd__mux2_1 _39315_ (.A0(\reg_next_pc[31] ),
    .A1(_01554_),
    .S(latched_store),
    .X(_01555_));
 sky130_fd_sc_hd__mux2_1 _39316_ (.A0(\reg_out[31] ),
    .A1(\alu_out_q[31] ),
    .S(latched_stalu),
    .X(_01554_));
 sky130_fd_sc_hd__mux2_1 _39317_ (.A0(\reg_next_pc[30] ),
    .A1(_01551_),
    .S(latched_store),
    .X(_01552_));
 sky130_fd_sc_hd__mux2_1 _39318_ (.A0(\reg_out[30] ),
    .A1(\alu_out_q[30] ),
    .S(latched_stalu),
    .X(_01551_));
 sky130_fd_sc_hd__mux2_1 _39319_ (.A0(\reg_next_pc[29] ),
    .A1(_01548_),
    .S(latched_store),
    .X(_01549_));
 sky130_fd_sc_hd__mux2_1 _39320_ (.A0(\reg_out[29] ),
    .A1(\alu_out_q[29] ),
    .S(latched_stalu),
    .X(_01548_));
 sky130_fd_sc_hd__mux2_1 _39321_ (.A0(\reg_next_pc[28] ),
    .A1(_01545_),
    .S(latched_store),
    .X(_01546_));
 sky130_fd_sc_hd__mux2_1 _39322_ (.A0(\reg_out[28] ),
    .A1(\alu_out_q[28] ),
    .S(latched_stalu),
    .X(_01545_));
 sky130_fd_sc_hd__mux2_1 _39323_ (.A0(\reg_next_pc[27] ),
    .A1(_01542_),
    .S(latched_store),
    .X(_01543_));
 sky130_fd_sc_hd__mux2_1 _39324_ (.A0(\reg_out[27] ),
    .A1(\alu_out_q[27] ),
    .S(latched_stalu),
    .X(_01542_));
 sky130_fd_sc_hd__mux2_1 _39325_ (.A0(\reg_next_pc[26] ),
    .A1(_01539_),
    .S(latched_store),
    .X(_01540_));
 sky130_fd_sc_hd__mux2_1 _39326_ (.A0(\reg_out[26] ),
    .A1(\alu_out_q[26] ),
    .S(latched_stalu),
    .X(_01539_));
 sky130_fd_sc_hd__mux2_1 _39327_ (.A0(\reg_next_pc[25] ),
    .A1(_01536_),
    .S(latched_store),
    .X(_01537_));
 sky130_fd_sc_hd__mux2_1 _39328_ (.A0(\reg_out[25] ),
    .A1(\alu_out_q[25] ),
    .S(latched_stalu),
    .X(_01536_));
 sky130_fd_sc_hd__mux2_1 _39329_ (.A0(\reg_next_pc[24] ),
    .A1(_01533_),
    .S(latched_store),
    .X(_01534_));
 sky130_fd_sc_hd__mux2_1 _39330_ (.A0(\reg_out[24] ),
    .A1(\alu_out_q[24] ),
    .S(latched_stalu),
    .X(_01533_));
 sky130_fd_sc_hd__mux2_1 _39331_ (.A0(\reg_next_pc[23] ),
    .A1(_01530_),
    .S(latched_store),
    .X(_01531_));
 sky130_fd_sc_hd__mux2_1 _39332_ (.A0(\reg_out[23] ),
    .A1(\alu_out_q[23] ),
    .S(latched_stalu),
    .X(_01530_));
 sky130_fd_sc_hd__mux2_1 _39333_ (.A0(\reg_next_pc[22] ),
    .A1(_01527_),
    .S(latched_store),
    .X(_01528_));
 sky130_fd_sc_hd__mux2_1 _39334_ (.A0(\reg_out[22] ),
    .A1(\alu_out_q[22] ),
    .S(latched_stalu),
    .X(_01527_));
 sky130_fd_sc_hd__mux2_1 _39335_ (.A0(\reg_next_pc[21] ),
    .A1(_01524_),
    .S(latched_store),
    .X(_01525_));
 sky130_fd_sc_hd__mux2_1 _39336_ (.A0(\reg_out[21] ),
    .A1(\alu_out_q[21] ),
    .S(latched_stalu),
    .X(_01524_));
 sky130_fd_sc_hd__mux2_1 _39337_ (.A0(\reg_next_pc[20] ),
    .A1(_01521_),
    .S(latched_store),
    .X(_01522_));
 sky130_fd_sc_hd__mux2_1 _39338_ (.A0(\reg_out[20] ),
    .A1(\alu_out_q[20] ),
    .S(latched_stalu),
    .X(_01521_));
 sky130_fd_sc_hd__mux2_1 _39339_ (.A0(\reg_next_pc[19] ),
    .A1(_01518_),
    .S(latched_store),
    .X(_01519_));
 sky130_fd_sc_hd__mux2_1 _39340_ (.A0(\reg_out[19] ),
    .A1(\alu_out_q[19] ),
    .S(latched_stalu),
    .X(_01518_));
 sky130_fd_sc_hd__mux2_1 _39341_ (.A0(\reg_next_pc[18] ),
    .A1(_01515_),
    .S(latched_store),
    .X(_01516_));
 sky130_fd_sc_hd__mux2_1 _39342_ (.A0(\reg_out[18] ),
    .A1(\alu_out_q[18] ),
    .S(latched_stalu),
    .X(_01515_));
 sky130_fd_sc_hd__mux2_1 _39343_ (.A0(\reg_next_pc[17] ),
    .A1(_01512_),
    .S(latched_store),
    .X(_01513_));
 sky130_fd_sc_hd__mux2_1 _39344_ (.A0(\reg_out[17] ),
    .A1(\alu_out_q[17] ),
    .S(latched_stalu),
    .X(_01512_));
 sky130_fd_sc_hd__mux2_1 _39345_ (.A0(\reg_next_pc[16] ),
    .A1(_01509_),
    .S(latched_store),
    .X(_01510_));
 sky130_fd_sc_hd__mux2_1 _39346_ (.A0(\reg_out[16] ),
    .A1(\alu_out_q[16] ),
    .S(latched_stalu),
    .X(_01509_));
 sky130_fd_sc_hd__mux2_1 _39347_ (.A0(\reg_next_pc[15] ),
    .A1(_01506_),
    .S(latched_store),
    .X(_01507_));
 sky130_fd_sc_hd__mux2_1 _39348_ (.A0(\reg_out[15] ),
    .A1(\alu_out_q[15] ),
    .S(latched_stalu),
    .X(_01506_));
 sky130_fd_sc_hd__mux2_1 _39349_ (.A0(\reg_next_pc[14] ),
    .A1(_01503_),
    .S(latched_store),
    .X(_01504_));
 sky130_fd_sc_hd__mux2_1 _39350_ (.A0(\reg_out[14] ),
    .A1(\alu_out_q[14] ),
    .S(latched_stalu),
    .X(_01503_));
 sky130_fd_sc_hd__mux2_1 _39351_ (.A0(\reg_next_pc[13] ),
    .A1(_01500_),
    .S(latched_store),
    .X(_01501_));
 sky130_fd_sc_hd__mux2_1 _39352_ (.A0(\reg_out[13] ),
    .A1(\alu_out_q[13] ),
    .S(latched_stalu),
    .X(_01500_));
 sky130_fd_sc_hd__mux2_1 _39353_ (.A0(\reg_next_pc[12] ),
    .A1(_01497_),
    .S(latched_store),
    .X(_01498_));
 sky130_fd_sc_hd__mux2_1 _39354_ (.A0(\reg_out[12] ),
    .A1(\alu_out_q[12] ),
    .S(latched_stalu),
    .X(_01497_));
 sky130_fd_sc_hd__mux2_1 _39355_ (.A0(\reg_next_pc[11] ),
    .A1(_01494_),
    .S(latched_store),
    .X(_01495_));
 sky130_fd_sc_hd__mux2_1 _39356_ (.A0(\reg_out[11] ),
    .A1(\alu_out_q[11] ),
    .S(latched_stalu),
    .X(_01494_));
 sky130_fd_sc_hd__mux2_1 _39357_ (.A0(\reg_next_pc[10] ),
    .A1(_01491_),
    .S(latched_store),
    .X(_01492_));
 sky130_fd_sc_hd__mux2_1 _39358_ (.A0(\reg_out[10] ),
    .A1(\alu_out_q[10] ),
    .S(latched_stalu),
    .X(_01491_));
 sky130_fd_sc_hd__mux2_1 _39359_ (.A0(\reg_next_pc[9] ),
    .A1(_01488_),
    .S(latched_store),
    .X(_01489_));
 sky130_fd_sc_hd__mux2_1 _39360_ (.A0(\reg_out[9] ),
    .A1(\alu_out_q[9] ),
    .S(latched_stalu),
    .X(_01488_));
 sky130_fd_sc_hd__mux2_1 _39361_ (.A0(\reg_next_pc[8] ),
    .A1(_01485_),
    .S(latched_store),
    .X(_01486_));
 sky130_fd_sc_hd__mux2_1 _39362_ (.A0(\reg_out[8] ),
    .A1(\alu_out_q[8] ),
    .S(latched_stalu),
    .X(_01485_));
 sky130_fd_sc_hd__mux2_1 _39363_ (.A0(\reg_next_pc[7] ),
    .A1(_01482_),
    .S(latched_store),
    .X(_01483_));
 sky130_fd_sc_hd__mux2_1 _39364_ (.A0(\reg_out[7] ),
    .A1(\alu_out_q[7] ),
    .S(latched_stalu),
    .X(_01482_));
 sky130_fd_sc_hd__mux2_1 _39365_ (.A0(\reg_next_pc[6] ),
    .A1(_01479_),
    .S(latched_store),
    .X(_01480_));
 sky130_fd_sc_hd__mux2_1 _39366_ (.A0(\reg_out[6] ),
    .A1(\alu_out_q[6] ),
    .S(latched_stalu),
    .X(_01479_));
 sky130_fd_sc_hd__mux2_1 _39367_ (.A0(\reg_next_pc[5] ),
    .A1(_01476_),
    .S(latched_store),
    .X(_01477_));
 sky130_fd_sc_hd__mux2_1 _39368_ (.A0(\reg_out[5] ),
    .A1(\alu_out_q[5] ),
    .S(latched_stalu),
    .X(_01476_));
 sky130_fd_sc_hd__mux2_1 _39369_ (.A0(_01474_),
    .A1(_01471_),
    .S(_00292_),
    .X(_01475_));
 sky130_fd_sc_hd__mux2_1 _39370_ (.A0(\reg_next_pc[4] ),
    .A1(_01472_),
    .S(latched_store),
    .X(_01473_));
 sky130_fd_sc_hd__mux2_1 _39371_ (.A0(\reg_out[4] ),
    .A1(\alu_out_q[4] ),
    .S(latched_stalu),
    .X(_01472_));
 sky130_fd_sc_hd__mux2_1 _39372_ (.A0(\reg_next_pc[3] ),
    .A1(_01468_),
    .S(latched_store),
    .X(_01469_));
 sky130_fd_sc_hd__mux2_1 _39373_ (.A0(\reg_out[3] ),
    .A1(\alu_out_q[3] ),
    .S(latched_stalu),
    .X(_01468_));
 sky130_fd_sc_hd__mux2_1 _39374_ (.A0(\reg_next_pc[1] ),
    .A1(_01465_),
    .S(latched_store),
    .X(_01466_));
 sky130_fd_sc_hd__mux2_1 _39375_ (.A0(\reg_out[1] ),
    .A1(\alu_out_q[1] ),
    .S(latched_stalu),
    .X(_01465_));
 sky130_fd_sc_hd__mux2_1 _39376_ (.A0(_01301_),
    .A1(\timer[31] ),
    .S(_01208_),
    .X(_01302_));
 sky130_fd_sc_hd__mux2_1 _39377_ (.A0(_01298_),
    .A1(\timer[30] ),
    .S(_01208_),
    .X(_01299_));
 sky130_fd_sc_hd__mux2_1 _39378_ (.A0(_01295_),
    .A1(\timer[29] ),
    .S(_01208_),
    .X(_01296_));
 sky130_fd_sc_hd__mux2_1 _39379_ (.A0(_01292_),
    .A1(\timer[28] ),
    .S(_01208_),
    .X(_01293_));
 sky130_fd_sc_hd__mux2_1 _39380_ (.A0(_01289_),
    .A1(\timer[27] ),
    .S(_01208_),
    .X(_01290_));
 sky130_fd_sc_hd__mux2_1 _39381_ (.A0(_01286_),
    .A1(\timer[26] ),
    .S(_01208_),
    .X(_01287_));
 sky130_fd_sc_hd__mux2_1 _39382_ (.A0(_01283_),
    .A1(\timer[25] ),
    .S(_01208_),
    .X(_01284_));
 sky130_fd_sc_hd__mux2_1 _39383_ (.A0(_01280_),
    .A1(\timer[24] ),
    .S(_01208_),
    .X(_01281_));
 sky130_fd_sc_hd__mux2_1 _39384_ (.A0(_01277_),
    .A1(\timer[23] ),
    .S(_01208_),
    .X(_01278_));
 sky130_fd_sc_hd__mux2_1 _39385_ (.A0(_01274_),
    .A1(\timer[22] ),
    .S(_01208_),
    .X(_01275_));
 sky130_fd_sc_hd__mux2_1 _39386_ (.A0(_01271_),
    .A1(\timer[21] ),
    .S(_01208_),
    .X(_01272_));
 sky130_fd_sc_hd__mux2_1 _39387_ (.A0(_01268_),
    .A1(\timer[20] ),
    .S(_01208_),
    .X(_01269_));
 sky130_fd_sc_hd__mux2_1 _39388_ (.A0(_01265_),
    .A1(\timer[19] ),
    .S(_01208_),
    .X(_01266_));
 sky130_fd_sc_hd__mux2_1 _39389_ (.A0(_01262_),
    .A1(\timer[18] ),
    .S(_01208_),
    .X(_01263_));
 sky130_fd_sc_hd__mux2_1 _39390_ (.A0(_01259_),
    .A1(\timer[17] ),
    .S(_01208_),
    .X(_01260_));
 sky130_fd_sc_hd__mux2_1 _39391_ (.A0(_01256_),
    .A1(\timer[16] ),
    .S(_01208_),
    .X(_01257_));
 sky130_fd_sc_hd__mux2_1 _39392_ (.A0(_01253_),
    .A1(\timer[15] ),
    .S(_01208_),
    .X(_01254_));
 sky130_fd_sc_hd__mux2_1 _39393_ (.A0(_01250_),
    .A1(\timer[14] ),
    .S(_01208_),
    .X(_01251_));
 sky130_fd_sc_hd__mux2_1 _39394_ (.A0(_01247_),
    .A1(\timer[13] ),
    .S(_01208_),
    .X(_01248_));
 sky130_fd_sc_hd__mux2_1 _39395_ (.A0(_01244_),
    .A1(\timer[12] ),
    .S(_01208_),
    .X(_01245_));
 sky130_fd_sc_hd__mux2_1 _39396_ (.A0(_01241_),
    .A1(\timer[11] ),
    .S(_01208_),
    .X(_01242_));
 sky130_fd_sc_hd__mux2_1 _39397_ (.A0(_01238_),
    .A1(\timer[10] ),
    .S(_01208_),
    .X(_01239_));
 sky130_fd_sc_hd__mux2_1 _39398_ (.A0(_01235_),
    .A1(\timer[9] ),
    .S(_01208_),
    .X(_01236_));
 sky130_fd_sc_hd__mux2_1 _39399_ (.A0(_01232_),
    .A1(\timer[8] ),
    .S(_01208_),
    .X(_01233_));
 sky130_fd_sc_hd__mux2_1 _39400_ (.A0(_01229_),
    .A1(\timer[7] ),
    .S(_01208_),
    .X(_01230_));
 sky130_fd_sc_hd__mux2_1 _39401_ (.A0(_01226_),
    .A1(\timer[6] ),
    .S(_01208_),
    .X(_01227_));
 sky130_fd_sc_hd__mux2_1 _39402_ (.A0(_01223_),
    .A1(\timer[5] ),
    .S(_01208_),
    .X(_01224_));
 sky130_fd_sc_hd__mux2_1 _39403_ (.A0(_01220_),
    .A1(\timer[4] ),
    .S(_01208_),
    .X(_01221_));
 sky130_fd_sc_hd__mux2_1 _39404_ (.A0(_01217_),
    .A1(\timer[3] ),
    .S(_01208_),
    .X(_01218_));
 sky130_fd_sc_hd__mux2_1 _39405_ (.A0(_01214_),
    .A1(\timer[2] ),
    .S(_01208_),
    .X(_01215_));
 sky130_fd_sc_hd__mux2_1 _39406_ (.A0(_01211_),
    .A1(\timer[1] ),
    .S(_01208_),
    .X(_01212_));
 sky130_fd_sc_hd__mux2_1 _39407_ (.A0(_01206_),
    .A1(_01201_),
    .S(_00368_),
    .X(_01207_));
 sky130_fd_sc_hd__mux2_1 _39408_ (.A0(_01179_),
    .A1(_01174_),
    .S(_00368_),
    .X(_01180_));
 sky130_fd_sc_hd__mux2_1 _39409_ (.A0(_01152_),
    .A1(_01147_),
    .S(_00368_),
    .X(_01153_));
 sky130_fd_sc_hd__mux2_1 _39410_ (.A0(_01125_),
    .A1(_01120_),
    .S(_00368_),
    .X(_01126_));
 sky130_fd_sc_hd__mux2_1 _39411_ (.A0(_01098_),
    .A1(_01093_),
    .S(_00368_),
    .X(_01099_));
 sky130_fd_sc_hd__mux2_1 _39412_ (.A0(_01071_),
    .A1(_01066_),
    .S(_00368_),
    .X(_01072_));
 sky130_fd_sc_hd__mux2_1 _39413_ (.A0(_01044_),
    .A1(_01039_),
    .S(_00368_),
    .X(_01045_));
 sky130_fd_sc_hd__mux2_1 _39414_ (.A0(_01017_),
    .A1(_01012_),
    .S(_00368_),
    .X(_01018_));
 sky130_fd_sc_hd__mux2_1 _39415_ (.A0(_00990_),
    .A1(_00985_),
    .S(_00368_),
    .X(_00991_));
 sky130_fd_sc_hd__mux2_1 _39416_ (.A0(_00963_),
    .A1(_00958_),
    .S(_00368_),
    .X(_00964_));
 sky130_fd_sc_hd__mux2_1 _39417_ (.A0(_00936_),
    .A1(_00931_),
    .S(_00368_),
    .X(_00937_));
 sky130_fd_sc_hd__mux2_1 _39418_ (.A0(_00909_),
    .A1(_00904_),
    .S(_00368_),
    .X(_00910_));
 sky130_fd_sc_hd__mux2_1 _39419_ (.A0(_00882_),
    .A1(_00877_),
    .S(_00368_),
    .X(_00883_));
 sky130_fd_sc_hd__mux2_1 _39420_ (.A0(_00855_),
    .A1(_00850_),
    .S(_00368_),
    .X(_00856_));
 sky130_fd_sc_hd__mux2_1 _39421_ (.A0(_00828_),
    .A1(_00823_),
    .S(_00368_),
    .X(_00829_));
 sky130_fd_sc_hd__mux2_1 _39422_ (.A0(_00801_),
    .A1(_00796_),
    .S(_00368_),
    .X(_00802_));
 sky130_fd_sc_hd__mux2_1 _39423_ (.A0(_00774_),
    .A1(_00769_),
    .S(_00368_),
    .X(_00775_));
 sky130_fd_sc_hd__mux2_1 _39424_ (.A0(_00747_),
    .A1(_00742_),
    .S(_00368_),
    .X(_00748_));
 sky130_fd_sc_hd__mux2_1 _39425_ (.A0(_00720_),
    .A1(_00715_),
    .S(_00368_),
    .X(_00721_));
 sky130_fd_sc_hd__mux2_1 _39426_ (.A0(_00693_),
    .A1(_00688_),
    .S(_00368_),
    .X(_00694_));
 sky130_fd_sc_hd__mux2_1 _39427_ (.A0(_00666_),
    .A1(_00661_),
    .S(_00368_),
    .X(_00667_));
 sky130_fd_sc_hd__mux2_1 _39428_ (.A0(_00639_),
    .A1(_00634_),
    .S(_00368_),
    .X(_00640_));
 sky130_fd_sc_hd__mux2_1 _39429_ (.A0(_00612_),
    .A1(_00607_),
    .S(_00368_),
    .X(_00613_));
 sky130_fd_sc_hd__mux2_1 _39430_ (.A0(_00585_),
    .A1(_00580_),
    .S(_00368_),
    .X(_00586_));
 sky130_fd_sc_hd__mux2_1 _39431_ (.A0(_00558_),
    .A1(_00553_),
    .S(_00368_),
    .X(_00559_));
 sky130_fd_sc_hd__mux2_1 _39432_ (.A0(_00531_),
    .A1(_00526_),
    .S(_00368_),
    .X(_00532_));
 sky130_fd_sc_hd__mux2_1 _39433_ (.A0(_00504_),
    .A1(_00499_),
    .S(_00368_),
    .X(_00505_));
 sky130_fd_sc_hd__mux2_1 _39434_ (.A0(_00477_),
    .A1(_00472_),
    .S(_00368_),
    .X(_00478_));
 sky130_fd_sc_hd__mux2_1 _39435_ (.A0(_00450_),
    .A1(_00445_),
    .S(_00368_),
    .X(_00451_));
 sky130_fd_sc_hd__mux2_1 _39436_ (.A0(_00423_),
    .A1(_00418_),
    .S(_00368_),
    .X(_00424_));
 sky130_fd_sc_hd__mux2_1 _39437_ (.A0(_00396_),
    .A1(_00391_),
    .S(_00368_),
    .X(_00397_));
 sky130_fd_sc_hd__mux2_1 _39438_ (.A0(_00369_),
    .A1(_00365_),
    .S(_00368_),
    .X(_00370_));
 sky130_fd_sc_hd__mux2_1 _39439_ (.A0(_00366_),
    .A1(_00367_),
    .S(\cpu_state[3] ),
    .X(_00368_));
 sky130_fd_sc_hd__mux2_1 _39440_ (.A0(\decoded_rs1[3] ),
    .A1(\decoded_imm_uj[3] ),
    .S(\cpu_state[3] ),
    .X(_00362_));
 sky130_fd_sc_hd__mux2_1 _39441_ (.A0(\decoded_rs1[2] ),
    .A1(\decoded_imm_uj[2] ),
    .S(\cpu_state[3] ),
    .X(_00360_));
 sky130_fd_sc_hd__mux2_1 _39442_ (.A0(\decoded_rs1[1] ),
    .A1(\decoded_imm_uj[1] ),
    .S(\cpu_state[3] ),
    .X(_00358_));
 sky130_fd_sc_hd__mux2_1 _39443_ (.A0(\decoded_rs1[0] ),
    .A1(\decoded_imm_uj[11] ),
    .S(\cpu_state[3] ),
    .X(_00357_));
 sky130_fd_sc_hd__mux2_1 _39444_ (.A0(_00349_),
    .A1(_00323_),
    .S(decoder_trigger),
    .X(_00350_));
 sky130_fd_sc_hd__mux2_1 _39445_ (.A0(_00350_),
    .A1(_00351_),
    .S(_00309_),
    .X(_00352_));
 sky130_fd_sc_hd__mux2_1 _39446_ (.A0(_00352_),
    .A1(_00349_),
    .S(_00308_),
    .X(_00353_));
 sky130_fd_sc_hd__mux2_1 _39447_ (.A0(_00355_),
    .A1(_00353_),
    .S(_00354_),
    .X(_00356_));
 sky130_fd_sc_hd__mux2_1 _39448_ (.A0(_00337_),
    .A1(_00344_),
    .S(is_beq_bne_blt_bge_bltu_bgeu),
    .X(_00345_));
 sky130_fd_sc_hd__mux2_1 _39449_ (.A0(_00345_),
    .A1(_00337_),
    .S(alu_wait),
    .X(_00346_));
 sky130_fd_sc_hd__mux2_1 _39450_ (.A0(_00342_),
    .A1(_00340_),
    .S(_00341_),
    .X(_00343_));
 sky130_fd_sc_hd__mux2_1 _39451_ (.A0(_00338_),
    .A1(_00337_),
    .S(_00296_),
    .X(_00339_));
 sky130_fd_sc_hd__mux2_1 _39452_ (.A0(\mem_rdata_q[12] ),
    .A1(_00334_),
    .S(\mem_rdata_q[13] ),
    .X(_00335_));
 sky130_fd_sc_hd__mux2_1 _39453_ (.A0(\cpu_state[1] ),
    .A1(_00302_),
    .S(\cpu_state[4] ),
    .X(_00333_));
 sky130_fd_sc_hd__mux2_1 _39454_ (.A0(_00322_),
    .A1(_00296_),
    .S(\cpu_state[6] ),
    .X(_00332_));
 sky130_fd_sc_hd__mux2_1 _39455_ (.A0(_00315_),
    .A1(alu_wait),
    .S(\cpu_state[4] ),
    .X(_00331_));
 sky130_fd_sc_hd__mux2_1 _39456_ (.A0(\mem_rdata_q[6] ),
    .A1(mem_rdata[6]),
    .S(mem_xfer),
    .X(_00330_));
 sky130_fd_sc_hd__mux2_1 _39457_ (.A0(\mem_rdata_q[5] ),
    .A1(mem_rdata[5]),
    .S(mem_xfer),
    .X(_00329_));
 sky130_fd_sc_hd__mux2_1 _39458_ (.A0(\mem_rdata_q[4] ),
    .A1(mem_rdata[4]),
    .S(mem_xfer),
    .X(_00328_));
 sky130_fd_sc_hd__mux2_1 _39459_ (.A0(\mem_rdata_q[3] ),
    .A1(mem_rdata[3]),
    .S(mem_xfer),
    .X(_00327_));
 sky130_fd_sc_hd__mux2_1 _39460_ (.A0(\mem_rdata_q[2] ),
    .A1(mem_rdata[2]),
    .S(mem_xfer),
    .X(_00326_));
 sky130_fd_sc_hd__mux2_1 _39461_ (.A0(\mem_rdata_q[1] ),
    .A1(mem_rdata[1]),
    .S(mem_xfer),
    .X(_00325_));
 sky130_fd_sc_hd__mux2_1 _39462_ (.A0(\mem_rdata_q[0] ),
    .A1(mem_rdata[0]),
    .S(mem_xfer),
    .X(_00324_));
 sky130_fd_sc_hd__mux2_1 _39463_ (.A0(\cpu_state[1] ),
    .A1(instr_retirq),
    .S(\cpu_state[2] ),
    .X(_00321_));
 sky130_fd_sc_hd__mux2_1 _39464_ (.A0(_00319_),
    .A1(\cpu_state[5] ),
    .S(_00296_),
    .X(_00320_));
 sky130_fd_sc_hd__mux2_1 _39465_ (.A0(_00317_),
    .A1(\cpu_state[6] ),
    .S(_00296_),
    .X(_00318_));
 sky130_fd_sc_hd__mux2_1 _39466_ (.A0(_00313_),
    .A1(_00312_),
    .S(_00307_),
    .X(_00314_));
 sky130_fd_sc_hd__mux2_1 _39467_ (.A0(_00298_),
    .A1(_00299_),
    .S(_00289_),
    .X(_00300_));
 sky130_fd_sc_hd__mux2_1 _39468_ (.A0(\reg_next_pc[2] ),
    .A1(_00293_),
    .S(latched_store),
    .X(_00294_));
 sky130_fd_sc_hd__mux2_1 _39469_ (.A0(\reg_out[2] ),
    .A1(\alu_out_q[2] ),
    .S(latched_stalu),
    .X(_00293_));
 sky130_fd_sc_hd__mux2_1 _39470_ (.A0(_00126_),
    .A1(_00122_),
    .S(mem_la_wdata[3]),
    .X(_02558_));
 sky130_fd_sc_hd__mux2_1 _39471_ (.A0(_00120_),
    .A1(_00116_),
    .S(mem_la_wdata[3]),
    .X(_02557_));
 sky130_fd_sc_hd__mux2_1 _39472_ (.A0(_00114_),
    .A1(_00110_),
    .S(mem_la_wdata[3]),
    .X(_02556_));
 sky130_fd_sc_hd__mux2_1 _39473_ (.A0(_00108_),
    .A1(_00104_),
    .S(mem_la_wdata[3]),
    .X(_02555_));
 sky130_fd_sc_hd__mux2_1 _39474_ (.A0(_00102_),
    .A1(_00095_),
    .S(mem_la_wdata[3]),
    .X(_02554_));
 sky130_fd_sc_hd__mux2_1 _39475_ (.A0(_00092_),
    .A1(_00085_),
    .S(mem_la_wdata[3]),
    .X(_02553_));
 sky130_fd_sc_hd__mux2_1 _39476_ (.A0(_00082_),
    .A1(_00068_),
    .S(mem_la_wdata[3]),
    .X(_02552_));
 sky130_fd_sc_hd__mux2_1 _39477_ (.A0(_00064_),
    .A1(_00050_),
    .S(mem_la_wdata[3]),
    .X(_02551_));
 sky130_fd_sc_hd__mux2_1 _39478_ (.A0(_01694_),
    .A1(_01695_),
    .S(_00290_),
    .X(_02541_));
 sky130_fd_sc_hd__mux2_1 _39479_ (.A0(_01691_),
    .A1(_01692_),
    .S(_00290_),
    .X(_02540_));
 sky130_fd_sc_hd__mux2_1 _39480_ (.A0(_01688_),
    .A1(_01689_),
    .S(_00290_),
    .X(_02539_));
 sky130_fd_sc_hd__mux2_1 _39481_ (.A0(_01685_),
    .A1(_01686_),
    .S(_00290_),
    .X(_02538_));
 sky130_fd_sc_hd__mux2_1 _39482_ (.A0(_01679_),
    .A1(_01680_),
    .S(instr_jal),
    .X(_01681_));
 sky130_fd_sc_hd__mux2_1 _39483_ (.A0(_01682_),
    .A1(_02581_),
    .S(_00308_),
    .X(_02530_));
 sky130_fd_sc_hd__mux2_1 _39484_ (.A0(_01675_),
    .A1(_01676_),
    .S(instr_jal),
    .X(_01677_));
 sky130_fd_sc_hd__mux2_1 _39485_ (.A0(_01678_),
    .A1(_02580_),
    .S(_00308_),
    .X(_02529_));
 sky130_fd_sc_hd__mux2_1 _39486_ (.A0(_01671_),
    .A1(_01672_),
    .S(instr_jal),
    .X(_01673_));
 sky130_fd_sc_hd__mux2_1 _39487_ (.A0(_01674_),
    .A1(_02579_),
    .S(_00308_),
    .X(_02527_));
 sky130_fd_sc_hd__mux2_1 _39488_ (.A0(_01667_),
    .A1(_01668_),
    .S(instr_jal),
    .X(_01669_));
 sky130_fd_sc_hd__mux2_1 _39489_ (.A0(_01670_),
    .A1(_02578_),
    .S(_00308_),
    .X(_02526_));
 sky130_fd_sc_hd__mux2_1 _39490_ (.A0(_01663_),
    .A1(_01664_),
    .S(instr_jal),
    .X(_01665_));
 sky130_fd_sc_hd__mux2_1 _39491_ (.A0(_01666_),
    .A1(_02577_),
    .S(_00308_),
    .X(_02525_));
 sky130_fd_sc_hd__mux2_1 _39492_ (.A0(_01659_),
    .A1(_01660_),
    .S(instr_jal),
    .X(_01661_));
 sky130_fd_sc_hd__mux2_1 _39493_ (.A0(_01662_),
    .A1(_02576_),
    .S(_00308_),
    .X(_02524_));
 sky130_fd_sc_hd__mux2_1 _39494_ (.A0(_01655_),
    .A1(_01656_),
    .S(instr_jal),
    .X(_01657_));
 sky130_fd_sc_hd__mux2_1 _39495_ (.A0(_01658_),
    .A1(_02575_),
    .S(_00308_),
    .X(_02523_));
 sky130_fd_sc_hd__mux2_1 _39496_ (.A0(_01651_),
    .A1(_01652_),
    .S(instr_jal),
    .X(_01653_));
 sky130_fd_sc_hd__mux2_1 _39497_ (.A0(_01654_),
    .A1(_02574_),
    .S(_00308_),
    .X(_02522_));
 sky130_fd_sc_hd__mux2_1 _39498_ (.A0(_01647_),
    .A1(_01648_),
    .S(instr_jal),
    .X(_01649_));
 sky130_fd_sc_hd__mux2_1 _39499_ (.A0(_01650_),
    .A1(_02573_),
    .S(_00308_),
    .X(_02521_));
 sky130_fd_sc_hd__mux2_1 _39500_ (.A0(_01643_),
    .A1(_01644_),
    .S(instr_jal),
    .X(_01645_));
 sky130_fd_sc_hd__mux2_1 _39501_ (.A0(_01646_),
    .A1(_02572_),
    .S(_00308_),
    .X(_02520_));
 sky130_fd_sc_hd__mux2_1 _39502_ (.A0(_01639_),
    .A1(_01640_),
    .S(instr_jal),
    .X(_01641_));
 sky130_fd_sc_hd__mux2_1 _39503_ (.A0(_01642_),
    .A1(_02570_),
    .S(_00308_),
    .X(_02519_));
 sky130_fd_sc_hd__mux2_1 _39504_ (.A0(_01635_),
    .A1(_01636_),
    .S(instr_jal),
    .X(_01637_));
 sky130_fd_sc_hd__mux2_1 _39505_ (.A0(_01638_),
    .A1(_02569_),
    .S(_00308_),
    .X(_02518_));
 sky130_fd_sc_hd__mux2_1 _39506_ (.A0(_01631_),
    .A1(_01632_),
    .S(instr_jal),
    .X(_01633_));
 sky130_fd_sc_hd__mux2_1 _39507_ (.A0(_01634_),
    .A1(_02568_),
    .S(_00308_),
    .X(_02516_));
 sky130_fd_sc_hd__mux2_1 _39508_ (.A0(_01627_),
    .A1(_01628_),
    .S(instr_jal),
    .X(_01629_));
 sky130_fd_sc_hd__mux2_1 _39509_ (.A0(_01630_),
    .A1(_02567_),
    .S(_00308_),
    .X(_02515_));
 sky130_fd_sc_hd__mux2_1 _39510_ (.A0(_01623_),
    .A1(_01624_),
    .S(instr_jal),
    .X(_01625_));
 sky130_fd_sc_hd__mux2_1 _39511_ (.A0(_01626_),
    .A1(_02566_),
    .S(_00308_),
    .X(_02514_));
 sky130_fd_sc_hd__mux2_1 _39512_ (.A0(_01619_),
    .A1(_01620_),
    .S(instr_jal),
    .X(_01621_));
 sky130_fd_sc_hd__mux2_1 _39513_ (.A0(_01622_),
    .A1(_02565_),
    .S(_00308_),
    .X(_02513_));
 sky130_fd_sc_hd__mux2_1 _39514_ (.A0(_01615_),
    .A1(_01616_),
    .S(instr_jal),
    .X(_01617_));
 sky130_fd_sc_hd__mux2_1 _39515_ (.A0(_01618_),
    .A1(_02564_),
    .S(_00308_),
    .X(_02512_));
 sky130_fd_sc_hd__mux2_1 _39516_ (.A0(_01611_),
    .A1(_01612_),
    .S(instr_jal),
    .X(_01613_));
 sky130_fd_sc_hd__mux2_1 _39517_ (.A0(_01614_),
    .A1(_02563_),
    .S(_00308_),
    .X(_02511_));
 sky130_fd_sc_hd__mux2_1 _39518_ (.A0(_01607_),
    .A1(_01608_),
    .S(instr_jal),
    .X(_01609_));
 sky130_fd_sc_hd__mux2_1 _39519_ (.A0(_01610_),
    .A1(_02562_),
    .S(_00308_),
    .X(_02510_));
 sky130_fd_sc_hd__mux2_1 _39520_ (.A0(_01603_),
    .A1(_01604_),
    .S(instr_jal),
    .X(_01605_));
 sky130_fd_sc_hd__mux2_1 _39521_ (.A0(_01606_),
    .A1(_02561_),
    .S(_00308_),
    .X(_02509_));
 sky130_fd_sc_hd__mux2_1 _39522_ (.A0(_01599_),
    .A1(_01600_),
    .S(instr_jal),
    .X(_01601_));
 sky130_fd_sc_hd__mux2_1 _39523_ (.A0(_01602_),
    .A1(_02589_),
    .S(_00308_),
    .X(_02508_));
 sky130_fd_sc_hd__mux2_1 _39524_ (.A0(_01595_),
    .A1(_01596_),
    .S(instr_jal),
    .X(_01597_));
 sky130_fd_sc_hd__mux2_1 _39525_ (.A0(_01598_),
    .A1(_02588_),
    .S(_00308_),
    .X(_02507_));
 sky130_fd_sc_hd__mux2_1 _39526_ (.A0(_01591_),
    .A1(_01592_),
    .S(instr_jal),
    .X(_01593_));
 sky130_fd_sc_hd__mux2_1 _39527_ (.A0(_01594_),
    .A1(_02587_),
    .S(_00308_),
    .X(_02537_));
 sky130_fd_sc_hd__mux2_1 _39528_ (.A0(_01587_),
    .A1(_01588_),
    .S(instr_jal),
    .X(_01589_));
 sky130_fd_sc_hd__mux2_1 _39529_ (.A0(_01590_),
    .A1(_02586_),
    .S(_00308_),
    .X(_02536_));
 sky130_fd_sc_hd__mux2_1 _39530_ (.A0(_01583_),
    .A1(_01584_),
    .S(instr_jal),
    .X(_01585_));
 sky130_fd_sc_hd__mux2_1 _39531_ (.A0(_01586_),
    .A1(_02585_),
    .S(_00308_),
    .X(_02535_));
 sky130_fd_sc_hd__mux2_1 _39532_ (.A0(_01579_),
    .A1(_01580_),
    .S(instr_jal),
    .X(_01581_));
 sky130_fd_sc_hd__mux2_1 _39533_ (.A0(_01582_),
    .A1(_02584_),
    .S(_00308_),
    .X(_02534_));
 sky130_fd_sc_hd__mux2_1 _39534_ (.A0(_01575_),
    .A1(_01576_),
    .S(instr_jal),
    .X(_01577_));
 sky130_fd_sc_hd__mux2_1 _39535_ (.A0(_01578_),
    .A1(_02583_),
    .S(_00308_),
    .X(_02533_));
 sky130_fd_sc_hd__mux2_1 _39536_ (.A0(_01571_),
    .A1(_01572_),
    .S(instr_jal),
    .X(_01573_));
 sky130_fd_sc_hd__mux2_1 _39537_ (.A0(_01574_),
    .A1(_02582_),
    .S(_00308_),
    .X(_02532_));
 sky130_fd_sc_hd__mux2_1 _39538_ (.A0(_01567_),
    .A1(_01568_),
    .S(instr_jal),
    .X(_01569_));
 sky130_fd_sc_hd__mux2_1 _39539_ (.A0(_01570_),
    .A1(_02571_),
    .S(_00308_),
    .X(_02531_));
 sky130_fd_sc_hd__mux2_1 _39540_ (.A0(_01561_),
    .A1(_01562_),
    .S(instr_jal),
    .X(_01563_));
 sky130_fd_sc_hd__mux2_1 _39541_ (.A0(_02560_),
    .A1(_01563_),
    .S(decoder_trigger),
    .X(_01564_));
 sky130_fd_sc_hd__mux2_1 _39542_ (.A0(_01564_),
    .A1(_01565_),
    .S(_00309_),
    .X(_01566_));
 sky130_fd_sc_hd__mux2_1 _39543_ (.A0(_01566_),
    .A1(_02560_),
    .S(_00308_),
    .X(_02528_));
 sky130_fd_sc_hd__mux2_1 _39544_ (.A0(_02590_),
    .A1(_01557_),
    .S(instr_jal),
    .X(_01558_));
 sky130_fd_sc_hd__mux2_1 _39545_ (.A0(_02590_),
    .A1(_01558_),
    .S(decoder_trigger),
    .X(_01559_));
 sky130_fd_sc_hd__mux2_1 _39546_ (.A0(_01559_),
    .A1(_02590_),
    .S(_00309_),
    .X(_01560_));
 sky130_fd_sc_hd__mux2_1 _39547_ (.A0(_01560_),
    .A1(_02590_),
    .S(_00308_),
    .X(_02517_));
 sky130_fd_sc_hd__mux2_1 _39548_ (.A0(\cpuregs_rs1[31] ),
    .A1(_01462_),
    .S(is_lui_auipc_jal),
    .X(_01463_));
 sky130_fd_sc_hd__mux2_1 _39549_ (.A0(_01464_),
    .A1(_01463_),
    .S(_00297_),
    .X(_02499_));
 sky130_fd_sc_hd__mux2_1 _39550_ (.A0(\cpuregs_rs1[30] ),
    .A1(_01459_),
    .S(is_lui_auipc_jal),
    .X(_01460_));
 sky130_fd_sc_hd__mux2_1 _39551_ (.A0(_01461_),
    .A1(_01460_),
    .S(_00297_),
    .X(_02498_));
 sky130_fd_sc_hd__mux2_1 _39552_ (.A0(\cpuregs_rs1[29] ),
    .A1(_01456_),
    .S(is_lui_auipc_jal),
    .X(_01457_));
 sky130_fd_sc_hd__mux2_1 _39553_ (.A0(_01458_),
    .A1(_01457_),
    .S(_00297_),
    .X(_02496_));
 sky130_fd_sc_hd__mux2_1 _39554_ (.A0(\cpuregs_rs1[28] ),
    .A1(_01453_),
    .S(is_lui_auipc_jal),
    .X(_01454_));
 sky130_fd_sc_hd__mux2_1 _39555_ (.A0(_01455_),
    .A1(_01454_),
    .S(_00297_),
    .X(_02495_));
 sky130_fd_sc_hd__mux2_1 _39556_ (.A0(\cpuregs_rs1[27] ),
    .A1(_01450_),
    .S(is_lui_auipc_jal),
    .X(_01451_));
 sky130_fd_sc_hd__mux2_1 _39557_ (.A0(_01452_),
    .A1(_01451_),
    .S(_00297_),
    .X(_02494_));
 sky130_fd_sc_hd__mux2_1 _39558_ (.A0(\cpuregs_rs1[26] ),
    .A1(_01447_),
    .S(is_lui_auipc_jal),
    .X(_01448_));
 sky130_fd_sc_hd__mux2_1 _39559_ (.A0(_01449_),
    .A1(_01448_),
    .S(_00297_),
    .X(_02493_));
 sky130_fd_sc_hd__mux2_1 _39560_ (.A0(\cpuregs_rs1[25] ),
    .A1(_01444_),
    .S(is_lui_auipc_jal),
    .X(_01445_));
 sky130_fd_sc_hd__mux2_1 _39561_ (.A0(_01446_),
    .A1(_01445_),
    .S(_00297_),
    .X(_02492_));
 sky130_fd_sc_hd__mux2_1 _39562_ (.A0(\cpuregs_rs1[24] ),
    .A1(_01441_),
    .S(is_lui_auipc_jal),
    .X(_01442_));
 sky130_fd_sc_hd__mux2_1 _39563_ (.A0(_01443_),
    .A1(_01442_),
    .S(_00297_),
    .X(_02491_));
 sky130_fd_sc_hd__mux2_1 _39564_ (.A0(\cpuregs_rs1[23] ),
    .A1(_01438_),
    .S(is_lui_auipc_jal),
    .X(_01439_));
 sky130_fd_sc_hd__mux2_1 _39565_ (.A0(_01440_),
    .A1(_01439_),
    .S(_00297_),
    .X(_02490_));
 sky130_fd_sc_hd__mux2_1 _39566_ (.A0(\cpuregs_rs1[22] ),
    .A1(_01435_),
    .S(is_lui_auipc_jal),
    .X(_01436_));
 sky130_fd_sc_hd__mux2_1 _39567_ (.A0(_01437_),
    .A1(_01436_),
    .S(_00297_),
    .X(_02489_));
 sky130_fd_sc_hd__mux2_1 _39568_ (.A0(\cpuregs_rs1[21] ),
    .A1(_01432_),
    .S(is_lui_auipc_jal),
    .X(_01433_));
 sky130_fd_sc_hd__mux2_1 _39569_ (.A0(_01434_),
    .A1(_01433_),
    .S(_00297_),
    .X(_02488_));
 sky130_fd_sc_hd__mux2_1 _39570_ (.A0(\cpuregs_rs1[20] ),
    .A1(_01429_),
    .S(is_lui_auipc_jal),
    .X(_01430_));
 sky130_fd_sc_hd__mux2_1 _39571_ (.A0(_01431_),
    .A1(_01430_),
    .S(_00297_),
    .X(_02487_));
 sky130_fd_sc_hd__mux2_1 _39572_ (.A0(\cpuregs_rs1[19] ),
    .A1(_01426_),
    .S(is_lui_auipc_jal),
    .X(_01427_));
 sky130_fd_sc_hd__mux2_1 _39573_ (.A0(_01428_),
    .A1(_01427_),
    .S(_00297_),
    .X(_02485_));
 sky130_fd_sc_hd__mux2_1 _39574_ (.A0(\cpuregs_rs1[18] ),
    .A1(_01423_),
    .S(is_lui_auipc_jal),
    .X(_01424_));
 sky130_fd_sc_hd__mux2_1 _39575_ (.A0(_01425_),
    .A1(_01424_),
    .S(_00297_),
    .X(_02484_));
 sky130_fd_sc_hd__mux2_1 _39576_ (.A0(\cpuregs_rs1[17] ),
    .A1(_01420_),
    .S(is_lui_auipc_jal),
    .X(_01421_));
 sky130_fd_sc_hd__mux2_1 _39577_ (.A0(_01422_),
    .A1(_01421_),
    .S(_00297_),
    .X(_02483_));
 sky130_fd_sc_hd__mux2_1 _39578_ (.A0(\cpuregs_rs1[16] ),
    .A1(_01417_),
    .S(is_lui_auipc_jal),
    .X(_01418_));
 sky130_fd_sc_hd__mux2_1 _39579_ (.A0(_01419_),
    .A1(_01418_),
    .S(_00297_),
    .X(_02482_));
 sky130_fd_sc_hd__mux2_1 _39580_ (.A0(\cpuregs_rs1[15] ),
    .A1(_01414_),
    .S(is_lui_auipc_jal),
    .X(_01415_));
 sky130_fd_sc_hd__mux2_1 _39581_ (.A0(_01416_),
    .A1(_01415_),
    .S(_00297_),
    .X(_02481_));
 sky130_fd_sc_hd__mux2_1 _39582_ (.A0(\cpuregs_rs1[14] ),
    .A1(_01411_),
    .S(is_lui_auipc_jal),
    .X(_01412_));
 sky130_fd_sc_hd__mux2_1 _39583_ (.A0(_01413_),
    .A1(_01412_),
    .S(_00297_),
    .X(_02480_));
 sky130_fd_sc_hd__mux2_1 _39584_ (.A0(\cpuregs_rs1[13] ),
    .A1(_01408_),
    .S(is_lui_auipc_jal),
    .X(_01409_));
 sky130_fd_sc_hd__mux2_1 _39585_ (.A0(_01410_),
    .A1(_01409_),
    .S(_00297_),
    .X(_02479_));
 sky130_fd_sc_hd__mux2_1 _39586_ (.A0(\cpuregs_rs1[12] ),
    .A1(_01405_),
    .S(is_lui_auipc_jal),
    .X(_01406_));
 sky130_fd_sc_hd__mux2_1 _39587_ (.A0(_01407_),
    .A1(_01406_),
    .S(_00297_),
    .X(_02478_));
 sky130_fd_sc_hd__mux2_1 _39588_ (.A0(\cpuregs_rs1[11] ),
    .A1(_01402_),
    .S(is_lui_auipc_jal),
    .X(_01403_));
 sky130_fd_sc_hd__mux2_1 _39589_ (.A0(_01404_),
    .A1(_01403_),
    .S(_00297_),
    .X(_02477_));
 sky130_fd_sc_hd__mux2_1 _39590_ (.A0(\cpuregs_rs1[10] ),
    .A1(_01399_),
    .S(is_lui_auipc_jal),
    .X(_01400_));
 sky130_fd_sc_hd__mux2_1 _39591_ (.A0(_01401_),
    .A1(_01400_),
    .S(_00297_),
    .X(_02476_));
 sky130_fd_sc_hd__mux2_1 _39592_ (.A0(\cpuregs_rs1[9] ),
    .A1(_01396_),
    .S(is_lui_auipc_jal),
    .X(_01397_));
 sky130_fd_sc_hd__mux2_1 _39593_ (.A0(_01398_),
    .A1(_01397_),
    .S(_00297_),
    .X(_02506_));
 sky130_fd_sc_hd__mux2_1 _39594_ (.A0(\cpuregs_rs1[8] ),
    .A1(_01393_),
    .S(is_lui_auipc_jal),
    .X(_01394_));
 sky130_fd_sc_hd__mux2_1 _39595_ (.A0(_01395_),
    .A1(_01394_),
    .S(_00297_),
    .X(_02505_));
 sky130_fd_sc_hd__mux2_1 _39596_ (.A0(\cpuregs_rs1[7] ),
    .A1(_01390_),
    .S(is_lui_auipc_jal),
    .X(_01391_));
 sky130_fd_sc_hd__mux2_1 _39597_ (.A0(_01392_),
    .A1(_01391_),
    .S(_00297_),
    .X(_02504_));
 sky130_fd_sc_hd__mux2_1 _39598_ (.A0(\cpuregs_rs1[6] ),
    .A1(_01387_),
    .S(is_lui_auipc_jal),
    .X(_01388_));
 sky130_fd_sc_hd__mux2_1 _39599_ (.A0(_01389_),
    .A1(_01388_),
    .S(_00297_),
    .X(_02503_));
 sky130_fd_sc_hd__mux2_1 _39600_ (.A0(\cpuregs_rs1[5] ),
    .A1(_01384_),
    .S(is_lui_auipc_jal),
    .X(_01385_));
 sky130_fd_sc_hd__mux2_1 _39601_ (.A0(_01386_),
    .A1(_01385_),
    .S(_00297_),
    .X(_02502_));
 sky130_fd_sc_hd__mux2_1 _39602_ (.A0(\cpuregs_rs1[4] ),
    .A1(_01381_),
    .S(is_lui_auipc_jal),
    .X(_01382_));
 sky130_fd_sc_hd__mux2_1 _39603_ (.A0(_01383_),
    .A1(_01382_),
    .S(_00297_),
    .X(_02501_));
 sky130_fd_sc_hd__mux2_1 _39604_ (.A0(\cpuregs_rs1[3] ),
    .A1(_01378_),
    .S(is_lui_auipc_jal),
    .X(_01379_));
 sky130_fd_sc_hd__mux2_1 _39605_ (.A0(_01380_),
    .A1(_01379_),
    .S(_00297_),
    .X(_02500_));
 sky130_fd_sc_hd__mux2_1 _39606_ (.A0(\cpuregs_rs1[2] ),
    .A1(_01375_),
    .S(is_lui_auipc_jal),
    .X(_01376_));
 sky130_fd_sc_hd__mux2_1 _39607_ (.A0(_01377_),
    .A1(_01376_),
    .S(_00297_),
    .X(_02497_));
 sky130_fd_sc_hd__mux2_1 _39608_ (.A0(\cpuregs_rs1[1] ),
    .A1(_01372_),
    .S(is_lui_auipc_jal),
    .X(_01373_));
 sky130_fd_sc_hd__mux2_1 _39609_ (.A0(_01374_),
    .A1(_01373_),
    .S(_00297_),
    .X(_02486_));
 sky130_fd_sc_hd__mux2_1 _39610_ (.A0(\cpuregs_rs1[0] ),
    .A1(_01369_),
    .S(is_lui_auipc_jal),
    .X(_01370_));
 sky130_fd_sc_hd__mux2_1 _39611_ (.A0(_01371_),
    .A1(_01370_),
    .S(_00297_),
    .X(_02475_));
 sky130_fd_sc_hd__mux2_1 _39612_ (.A0(_01367_),
    .A1(\decoded_imm[31] ),
    .S(_01304_),
    .X(_01368_));
 sky130_fd_sc_hd__mux2_1 _39613_ (.A0(_01368_),
    .A1(\cpuregs_rs1[31] ),
    .S(\cpu_state[3] ),
    .X(_02467_));
 sky130_fd_sc_hd__mux2_1 _39614_ (.A0(_01365_),
    .A1(\decoded_imm[30] ),
    .S(_01304_),
    .X(_01366_));
 sky130_fd_sc_hd__mux2_1 _39615_ (.A0(_01366_),
    .A1(\cpuregs_rs1[30] ),
    .S(\cpu_state[3] ),
    .X(_02466_));
 sky130_fd_sc_hd__mux2_1 _39616_ (.A0(_01363_),
    .A1(\decoded_imm[29] ),
    .S(_01304_),
    .X(_01364_));
 sky130_fd_sc_hd__mux2_1 _39617_ (.A0(_01364_),
    .A1(\cpuregs_rs1[29] ),
    .S(\cpu_state[3] ),
    .X(_02464_));
 sky130_fd_sc_hd__mux2_1 _39618_ (.A0(_01361_),
    .A1(\decoded_imm[28] ),
    .S(_01304_),
    .X(_01362_));
 sky130_fd_sc_hd__mux2_1 _39619_ (.A0(_01362_),
    .A1(\cpuregs_rs1[28] ),
    .S(\cpu_state[3] ),
    .X(_02463_));
 sky130_fd_sc_hd__mux2_1 _39620_ (.A0(_01359_),
    .A1(\decoded_imm[27] ),
    .S(_01304_),
    .X(_01360_));
 sky130_fd_sc_hd__mux2_1 _39621_ (.A0(_01360_),
    .A1(\cpuregs_rs1[27] ),
    .S(\cpu_state[3] ),
    .X(_02462_));
 sky130_fd_sc_hd__mux2_1 _39622_ (.A0(_01357_),
    .A1(\decoded_imm[26] ),
    .S(_01304_),
    .X(_01358_));
 sky130_fd_sc_hd__mux2_1 _39623_ (.A0(_01358_),
    .A1(\cpuregs_rs1[26] ),
    .S(\cpu_state[3] ),
    .X(_02461_));
 sky130_fd_sc_hd__mux2_1 _39624_ (.A0(_01355_),
    .A1(\decoded_imm[25] ),
    .S(_01304_),
    .X(_01356_));
 sky130_fd_sc_hd__mux2_1 _39625_ (.A0(_01356_),
    .A1(\cpuregs_rs1[25] ),
    .S(\cpu_state[3] ),
    .X(_02460_));
 sky130_fd_sc_hd__mux2_1 _39626_ (.A0(_01353_),
    .A1(\decoded_imm[24] ),
    .S(_01304_),
    .X(_01354_));
 sky130_fd_sc_hd__mux2_1 _39627_ (.A0(_01354_),
    .A1(\cpuregs_rs1[24] ),
    .S(\cpu_state[3] ),
    .X(_02459_));
 sky130_fd_sc_hd__mux2_1 _39628_ (.A0(_01351_),
    .A1(\decoded_imm[23] ),
    .S(_01304_),
    .X(_01352_));
 sky130_fd_sc_hd__mux2_1 _39629_ (.A0(_01352_),
    .A1(\cpuregs_rs1[23] ),
    .S(\cpu_state[3] ),
    .X(_02458_));
 sky130_fd_sc_hd__mux2_1 _39630_ (.A0(_01349_),
    .A1(\decoded_imm[22] ),
    .S(_01304_),
    .X(_01350_));
 sky130_fd_sc_hd__mux2_1 _39631_ (.A0(_01350_),
    .A1(\cpuregs_rs1[22] ),
    .S(\cpu_state[3] ),
    .X(_02457_));
 sky130_fd_sc_hd__mux2_1 _39632_ (.A0(_01347_),
    .A1(\decoded_imm[21] ),
    .S(_01304_),
    .X(_01348_));
 sky130_fd_sc_hd__mux2_1 _39633_ (.A0(_01348_),
    .A1(\cpuregs_rs1[21] ),
    .S(\cpu_state[3] ),
    .X(_02456_));
 sky130_fd_sc_hd__mux2_1 _39634_ (.A0(_01345_),
    .A1(\decoded_imm[20] ),
    .S(_01304_),
    .X(_01346_));
 sky130_fd_sc_hd__mux2_1 _39635_ (.A0(_01346_),
    .A1(\cpuregs_rs1[20] ),
    .S(\cpu_state[3] ),
    .X(_02455_));
 sky130_fd_sc_hd__mux2_1 _39636_ (.A0(_01343_),
    .A1(\decoded_imm[19] ),
    .S(_01304_),
    .X(_01344_));
 sky130_fd_sc_hd__mux2_1 _39637_ (.A0(_01344_),
    .A1(\cpuregs_rs1[19] ),
    .S(\cpu_state[3] ),
    .X(_02453_));
 sky130_fd_sc_hd__mux2_1 _39638_ (.A0(_01341_),
    .A1(\decoded_imm[18] ),
    .S(_01304_),
    .X(_01342_));
 sky130_fd_sc_hd__mux2_1 _39639_ (.A0(_01342_),
    .A1(\cpuregs_rs1[18] ),
    .S(\cpu_state[3] ),
    .X(_02452_));
 sky130_fd_sc_hd__mux2_1 _39640_ (.A0(_01339_),
    .A1(\decoded_imm[17] ),
    .S(_01304_),
    .X(_01340_));
 sky130_fd_sc_hd__mux2_1 _39641_ (.A0(_01340_),
    .A1(\cpuregs_rs1[17] ),
    .S(\cpu_state[3] ),
    .X(_02451_));
 sky130_fd_sc_hd__mux2_1 _39642_ (.A0(_01337_),
    .A1(\decoded_imm[16] ),
    .S(_01304_),
    .X(_01338_));
 sky130_fd_sc_hd__mux2_1 _39643_ (.A0(_01338_),
    .A1(\cpuregs_rs1[16] ),
    .S(\cpu_state[3] ),
    .X(_02450_));
 sky130_fd_sc_hd__mux2_1 _39644_ (.A0(_01335_),
    .A1(\decoded_imm[15] ),
    .S(_01304_),
    .X(_01336_));
 sky130_fd_sc_hd__mux2_1 _39645_ (.A0(_01336_),
    .A1(\cpuregs_rs1[15] ),
    .S(\cpu_state[3] ),
    .X(_02449_));
 sky130_fd_sc_hd__mux2_1 _39646_ (.A0(_01333_),
    .A1(\decoded_imm[14] ),
    .S(_01304_),
    .X(_01334_));
 sky130_fd_sc_hd__mux2_1 _39647_ (.A0(_01334_),
    .A1(\cpuregs_rs1[14] ),
    .S(\cpu_state[3] ),
    .X(_02448_));
 sky130_fd_sc_hd__mux2_1 _39648_ (.A0(_01331_),
    .A1(\decoded_imm[13] ),
    .S(_01304_),
    .X(_01332_));
 sky130_fd_sc_hd__mux2_1 _39649_ (.A0(_01332_),
    .A1(\cpuregs_rs1[13] ),
    .S(\cpu_state[3] ),
    .X(_02447_));
 sky130_fd_sc_hd__mux2_1 _39650_ (.A0(_01329_),
    .A1(\decoded_imm[12] ),
    .S(_01304_),
    .X(_01330_));
 sky130_fd_sc_hd__mux2_1 _39651_ (.A0(_01330_),
    .A1(\cpuregs_rs1[12] ),
    .S(\cpu_state[3] ),
    .X(_02446_));
 sky130_fd_sc_hd__mux2_1 _39652_ (.A0(_01327_),
    .A1(\decoded_imm[11] ),
    .S(_01304_),
    .X(_01328_));
 sky130_fd_sc_hd__mux2_1 _39653_ (.A0(_01328_),
    .A1(\cpuregs_rs1[11] ),
    .S(\cpu_state[3] ),
    .X(_02445_));
 sky130_fd_sc_hd__mux2_1 _39654_ (.A0(_01325_),
    .A1(\decoded_imm[10] ),
    .S(_01304_),
    .X(_01326_));
 sky130_fd_sc_hd__mux2_1 _39655_ (.A0(_01326_),
    .A1(\cpuregs_rs1[10] ),
    .S(\cpu_state[3] ),
    .X(_02444_));
 sky130_fd_sc_hd__mux2_1 _39656_ (.A0(_01323_),
    .A1(\decoded_imm[9] ),
    .S(_01304_),
    .X(_01324_));
 sky130_fd_sc_hd__mux2_1 _39657_ (.A0(_01324_),
    .A1(\cpuregs_rs1[9] ),
    .S(\cpu_state[3] ),
    .X(_02474_));
 sky130_fd_sc_hd__mux2_1 _39658_ (.A0(_01321_),
    .A1(\decoded_imm[8] ),
    .S(_01304_),
    .X(_01322_));
 sky130_fd_sc_hd__mux2_1 _39659_ (.A0(_01322_),
    .A1(\cpuregs_rs1[8] ),
    .S(\cpu_state[3] ),
    .X(_02473_));
 sky130_fd_sc_hd__mux2_1 _39660_ (.A0(_01319_),
    .A1(\decoded_imm[7] ),
    .S(_01304_),
    .X(_01320_));
 sky130_fd_sc_hd__mux2_1 _39661_ (.A0(_01320_),
    .A1(\cpuregs_rs1[7] ),
    .S(\cpu_state[3] ),
    .X(_02472_));
 sky130_fd_sc_hd__mux2_1 _39662_ (.A0(_01317_),
    .A1(\decoded_imm[6] ),
    .S(_01304_),
    .X(_01318_));
 sky130_fd_sc_hd__mux2_1 _39663_ (.A0(_01318_),
    .A1(\cpuregs_rs1[6] ),
    .S(\cpu_state[3] ),
    .X(_02471_));
 sky130_fd_sc_hd__mux2_1 _39664_ (.A0(_01315_),
    .A1(\decoded_imm[5] ),
    .S(_01304_),
    .X(_01316_));
 sky130_fd_sc_hd__mux2_1 _39665_ (.A0(_01316_),
    .A1(\cpuregs_rs1[5] ),
    .S(\cpu_state[3] ),
    .X(_02470_));
 sky130_fd_sc_hd__mux2_1 _39666_ (.A0(\decoded_imm[4] ),
    .A1(\decoded_imm_uj[4] ),
    .S(is_slli_srli_srai),
    .X(_01313_));
 sky130_fd_sc_hd__mux2_1 _39667_ (.A0(_01313_),
    .A1(\decoded_imm[4] ),
    .S(_01304_),
    .X(_01314_));
 sky130_fd_sc_hd__mux2_1 _39668_ (.A0(_01314_),
    .A1(\cpuregs_rs1[4] ),
    .S(\cpu_state[3] ),
    .X(_02469_));
 sky130_fd_sc_hd__mux2_1 _39669_ (.A0(\decoded_imm[3] ),
    .A1(\decoded_imm_uj[3] ),
    .S(is_slli_srli_srai),
    .X(_01311_));
 sky130_fd_sc_hd__mux2_1 _39670_ (.A0(_01311_),
    .A1(\decoded_imm[3] ),
    .S(_01304_),
    .X(_01312_));
 sky130_fd_sc_hd__mux2_1 _39671_ (.A0(_01312_),
    .A1(\cpuregs_rs1[3] ),
    .S(\cpu_state[3] ),
    .X(_02468_));
 sky130_fd_sc_hd__mux2_1 _39672_ (.A0(\decoded_imm[2] ),
    .A1(\decoded_imm_uj[2] ),
    .S(is_slli_srli_srai),
    .X(_01309_));
 sky130_fd_sc_hd__mux2_1 _39673_ (.A0(_01309_),
    .A1(\decoded_imm[2] ),
    .S(_01304_),
    .X(_01310_));
 sky130_fd_sc_hd__mux2_1 _39674_ (.A0(_01310_),
    .A1(\cpuregs_rs1[2] ),
    .S(\cpu_state[3] ),
    .X(_02465_));
 sky130_fd_sc_hd__mux2_1 _39675_ (.A0(\decoded_imm[1] ),
    .A1(\decoded_imm_uj[1] ),
    .S(is_slli_srli_srai),
    .X(_01307_));
 sky130_fd_sc_hd__mux2_1 _39676_ (.A0(_01307_),
    .A1(\decoded_imm[1] ),
    .S(_01304_),
    .X(_01308_));
 sky130_fd_sc_hd__mux2_1 _39677_ (.A0(_01308_),
    .A1(\cpuregs_rs1[1] ),
    .S(\cpu_state[3] ),
    .X(_02454_));
 sky130_fd_sc_hd__mux2_1 _39678_ (.A0(\decoded_imm[0] ),
    .A1(\decoded_imm_uj[11] ),
    .S(is_slli_srli_srai),
    .X(_01305_));
 sky130_fd_sc_hd__mux2_1 _39679_ (.A0(_01305_),
    .A1(\decoded_imm[0] ),
    .S(_01304_),
    .X(_01306_));
 sky130_fd_sc_hd__mux2_1 _39680_ (.A0(_01306_),
    .A1(\cpuregs_rs1[0] ),
    .S(\cpu_state[3] ),
    .X(_02443_));
 sky130_fd_sc_hd__mux2_1 _39681_ (.A0(_01302_),
    .A1(\cpuregs_rs1[31] ),
    .S(instr_timer),
    .X(_01303_));
 sky130_fd_sc_hd__mux2_1 _39682_ (.A0(_01302_),
    .A1(_01303_),
    .S(\cpu_state[2] ),
    .X(_02435_));
 sky130_fd_sc_hd__mux2_1 _39683_ (.A0(_01299_),
    .A1(\cpuregs_rs1[30] ),
    .S(instr_timer),
    .X(_01300_));
 sky130_fd_sc_hd__mux2_1 _39684_ (.A0(_01299_),
    .A1(_01300_),
    .S(\cpu_state[2] ),
    .X(_02434_));
 sky130_fd_sc_hd__mux2_1 _39685_ (.A0(_01296_),
    .A1(\cpuregs_rs1[29] ),
    .S(instr_timer),
    .X(_01297_));
 sky130_fd_sc_hd__mux2_1 _39686_ (.A0(_01296_),
    .A1(_01297_),
    .S(\cpu_state[2] ),
    .X(_02432_));
 sky130_fd_sc_hd__mux2_1 _39687_ (.A0(_01293_),
    .A1(\cpuregs_rs1[28] ),
    .S(instr_timer),
    .X(_01294_));
 sky130_fd_sc_hd__mux2_1 _39688_ (.A0(_01293_),
    .A1(_01294_),
    .S(\cpu_state[2] ),
    .X(_02431_));
 sky130_fd_sc_hd__mux2_1 _39689_ (.A0(_01290_),
    .A1(\cpuregs_rs1[27] ),
    .S(instr_timer),
    .X(_01291_));
 sky130_fd_sc_hd__mux2_1 _39690_ (.A0(_01290_),
    .A1(_01291_),
    .S(\cpu_state[2] ),
    .X(_02430_));
 sky130_fd_sc_hd__mux2_1 _39691_ (.A0(_01287_),
    .A1(\cpuregs_rs1[26] ),
    .S(instr_timer),
    .X(_01288_));
 sky130_fd_sc_hd__mux2_1 _39692_ (.A0(_01287_),
    .A1(_01288_),
    .S(\cpu_state[2] ),
    .X(_02429_));
 sky130_fd_sc_hd__mux2_1 _39693_ (.A0(_01284_),
    .A1(\cpuregs_rs1[25] ),
    .S(instr_timer),
    .X(_01285_));
 sky130_fd_sc_hd__mux2_1 _39694_ (.A0(_01284_),
    .A1(_01285_),
    .S(\cpu_state[2] ),
    .X(_02428_));
 sky130_fd_sc_hd__mux2_1 _39695_ (.A0(_01281_),
    .A1(\cpuregs_rs1[24] ),
    .S(instr_timer),
    .X(_01282_));
 sky130_fd_sc_hd__mux2_1 _39696_ (.A0(_01281_),
    .A1(_01282_),
    .S(\cpu_state[2] ),
    .X(_02427_));
 sky130_fd_sc_hd__mux2_1 _39697_ (.A0(_01278_),
    .A1(\cpuregs_rs1[23] ),
    .S(instr_timer),
    .X(_01279_));
 sky130_fd_sc_hd__mux2_1 _39698_ (.A0(_01278_),
    .A1(_01279_),
    .S(\cpu_state[2] ),
    .X(_02426_));
 sky130_fd_sc_hd__mux2_1 _39699_ (.A0(_01275_),
    .A1(\cpuregs_rs1[22] ),
    .S(instr_timer),
    .X(_01276_));
 sky130_fd_sc_hd__mux2_1 _39700_ (.A0(_01275_),
    .A1(_01276_),
    .S(\cpu_state[2] ),
    .X(_02425_));
 sky130_fd_sc_hd__mux2_1 _39701_ (.A0(_01272_),
    .A1(\cpuregs_rs1[21] ),
    .S(instr_timer),
    .X(_01273_));
 sky130_fd_sc_hd__mux2_1 _39702_ (.A0(_01272_),
    .A1(_01273_),
    .S(\cpu_state[2] ),
    .X(_02424_));
 sky130_fd_sc_hd__mux2_1 _39703_ (.A0(_01269_),
    .A1(\cpuregs_rs1[20] ),
    .S(instr_timer),
    .X(_01270_));
 sky130_fd_sc_hd__mux2_1 _39704_ (.A0(_01269_),
    .A1(_01270_),
    .S(\cpu_state[2] ),
    .X(_02423_));
 sky130_fd_sc_hd__mux2_1 _39705_ (.A0(_01266_),
    .A1(\cpuregs_rs1[19] ),
    .S(instr_timer),
    .X(_01267_));
 sky130_fd_sc_hd__mux2_1 _39706_ (.A0(_01266_),
    .A1(_01267_),
    .S(\cpu_state[2] ),
    .X(_02421_));
 sky130_fd_sc_hd__mux2_1 _39707_ (.A0(_01263_),
    .A1(\cpuregs_rs1[18] ),
    .S(instr_timer),
    .X(_01264_));
 sky130_fd_sc_hd__mux2_1 _39708_ (.A0(_01263_),
    .A1(_01264_),
    .S(\cpu_state[2] ),
    .X(_02420_));
 sky130_fd_sc_hd__mux2_1 _39709_ (.A0(_01260_),
    .A1(\cpuregs_rs1[17] ),
    .S(instr_timer),
    .X(_01261_));
 sky130_fd_sc_hd__mux2_1 _39710_ (.A0(_01260_),
    .A1(_01261_),
    .S(\cpu_state[2] ),
    .X(_02419_));
 sky130_fd_sc_hd__mux2_1 _39711_ (.A0(_01257_),
    .A1(\cpuregs_rs1[16] ),
    .S(instr_timer),
    .X(_01258_));
 sky130_fd_sc_hd__mux2_1 _39712_ (.A0(_01257_),
    .A1(_01258_),
    .S(\cpu_state[2] ),
    .X(_02418_));
 sky130_fd_sc_hd__mux2_1 _39713_ (.A0(_01254_),
    .A1(\cpuregs_rs1[15] ),
    .S(instr_timer),
    .X(_01255_));
 sky130_fd_sc_hd__mux2_1 _39714_ (.A0(_01254_),
    .A1(_01255_),
    .S(\cpu_state[2] ),
    .X(_02417_));
 sky130_fd_sc_hd__mux2_1 _39715_ (.A0(_01251_),
    .A1(\cpuregs_rs1[14] ),
    .S(instr_timer),
    .X(_01252_));
 sky130_fd_sc_hd__mux2_1 _39716_ (.A0(_01251_),
    .A1(_01252_),
    .S(\cpu_state[2] ),
    .X(_02416_));
 sky130_fd_sc_hd__mux2_1 _39717_ (.A0(_01248_),
    .A1(\cpuregs_rs1[13] ),
    .S(instr_timer),
    .X(_01249_));
 sky130_fd_sc_hd__mux2_1 _39718_ (.A0(_01248_),
    .A1(_01249_),
    .S(\cpu_state[2] ),
    .X(_02415_));
 sky130_fd_sc_hd__mux2_1 _39719_ (.A0(_01245_),
    .A1(\cpuregs_rs1[12] ),
    .S(instr_timer),
    .X(_01246_));
 sky130_fd_sc_hd__mux2_1 _39720_ (.A0(_01245_),
    .A1(_01246_),
    .S(\cpu_state[2] ),
    .X(_02414_));
 sky130_fd_sc_hd__mux2_1 _39721_ (.A0(_01242_),
    .A1(\cpuregs_rs1[11] ),
    .S(instr_timer),
    .X(_01243_));
 sky130_fd_sc_hd__mux2_1 _39722_ (.A0(_01242_),
    .A1(_01243_),
    .S(\cpu_state[2] ),
    .X(_02413_));
 sky130_fd_sc_hd__mux2_1 _39723_ (.A0(_01239_),
    .A1(\cpuregs_rs1[10] ),
    .S(instr_timer),
    .X(_01240_));
 sky130_fd_sc_hd__mux2_1 _39724_ (.A0(_01239_),
    .A1(_01240_),
    .S(\cpu_state[2] ),
    .X(_02412_));
 sky130_fd_sc_hd__mux2_1 _39725_ (.A0(_01236_),
    .A1(\cpuregs_rs1[9] ),
    .S(instr_timer),
    .X(_01237_));
 sky130_fd_sc_hd__mux2_1 _39726_ (.A0(_01236_),
    .A1(_01237_),
    .S(\cpu_state[2] ),
    .X(_02442_));
 sky130_fd_sc_hd__mux2_1 _39727_ (.A0(_01233_),
    .A1(\cpuregs_rs1[8] ),
    .S(instr_timer),
    .X(_01234_));
 sky130_fd_sc_hd__mux2_1 _39728_ (.A0(_01233_),
    .A1(_01234_),
    .S(\cpu_state[2] ),
    .X(_02441_));
 sky130_fd_sc_hd__mux2_1 _39729_ (.A0(_01230_),
    .A1(\cpuregs_rs1[7] ),
    .S(instr_timer),
    .X(_01231_));
 sky130_fd_sc_hd__mux2_1 _39730_ (.A0(_01230_),
    .A1(_01231_),
    .S(\cpu_state[2] ),
    .X(_02440_));
 sky130_fd_sc_hd__mux2_1 _39731_ (.A0(_01227_),
    .A1(\cpuregs_rs1[6] ),
    .S(instr_timer),
    .X(_01228_));
 sky130_fd_sc_hd__mux2_1 _39732_ (.A0(_01227_),
    .A1(_01228_),
    .S(\cpu_state[2] ),
    .X(_02439_));
 sky130_fd_sc_hd__mux2_1 _39733_ (.A0(_01224_),
    .A1(\cpuregs_rs1[5] ),
    .S(instr_timer),
    .X(_01225_));
 sky130_fd_sc_hd__mux2_1 _39734_ (.A0(_01224_),
    .A1(_01225_),
    .S(\cpu_state[2] ),
    .X(_02438_));
 sky130_fd_sc_hd__mux2_1 _39735_ (.A0(_01221_),
    .A1(\cpuregs_rs1[4] ),
    .S(instr_timer),
    .X(_01222_));
 sky130_fd_sc_hd__mux2_1 _39736_ (.A0(_01221_),
    .A1(_01222_),
    .S(\cpu_state[2] ),
    .X(_02437_));
 sky130_fd_sc_hd__mux2_1 _39737_ (.A0(_01218_),
    .A1(\cpuregs_rs1[3] ),
    .S(instr_timer),
    .X(_01219_));
 sky130_fd_sc_hd__mux2_1 _39738_ (.A0(_01218_),
    .A1(_01219_),
    .S(\cpu_state[2] ),
    .X(_02436_));
 sky130_fd_sc_hd__mux2_1 _39739_ (.A0(_01215_),
    .A1(\cpuregs_rs1[2] ),
    .S(instr_timer),
    .X(_01216_));
 sky130_fd_sc_hd__mux2_1 _39740_ (.A0(_01215_),
    .A1(_01216_),
    .S(\cpu_state[2] ),
    .X(_02433_));
 sky130_fd_sc_hd__mux2_1 _39741_ (.A0(_01212_),
    .A1(\cpuregs_rs1[1] ),
    .S(instr_timer),
    .X(_01213_));
 sky130_fd_sc_hd__mux2_1 _39742_ (.A0(_01212_),
    .A1(_01213_),
    .S(\cpu_state[2] ),
    .X(_02422_));
 sky130_fd_sc_hd__mux2_1 _39743_ (.A0(_01209_),
    .A1(\cpuregs_rs1[0] ),
    .S(instr_timer),
    .X(_01210_));
 sky130_fd_sc_hd__mux2_1 _39744_ (.A0(_01209_),
    .A1(_01210_),
    .S(\cpu_state[2] ),
    .X(_02411_));
 sky130_fd_sc_hd__mux4_1 _39745_ (.A0(_01202_),
    .A1(_01203_),
    .A2(_01204_),
    .A3(_01205_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_01206_));
 sky130_fd_sc_hd__mux4_1 _39746_ (.A0(_01181_),
    .A1(_01182_),
    .A2(_01183_),
    .A3(_01184_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_01185_));
 sky130_fd_sc_hd__mux4_1 _39747_ (.A0(_01186_),
    .A1(_01187_),
    .A2(_01188_),
    .A3(_01189_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_01190_));
 sky130_fd_sc_hd__mux4_1 _39748_ (.A0(_01191_),
    .A1(_01192_),
    .A2(_01193_),
    .A3(_01194_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_01195_));
 sky130_fd_sc_hd__mux4_1 _39749_ (.A0(_01196_),
    .A1(_01197_),
    .A2(_01198_),
    .A3(_01199_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_01200_));
 sky130_fd_sc_hd__mux4_1 _39750_ (.A0(_01185_),
    .A1(_01190_),
    .A2(_01195_),
    .A3(_01200_),
    .S0(_00360_),
    .S1(_00362_),
    .X(_01201_));
 sky130_fd_sc_hd__mux4_1 _39751_ (.A0(_01175_),
    .A1(_01176_),
    .A2(_01177_),
    .A3(_01178_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_01179_));
 sky130_fd_sc_hd__mux4_1 _39752_ (.A0(_01154_),
    .A1(_01155_),
    .A2(_01156_),
    .A3(_01157_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_01158_));
 sky130_fd_sc_hd__mux4_1 _39753_ (.A0(_01159_),
    .A1(_01160_),
    .A2(_01161_),
    .A3(_01162_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_01163_));
 sky130_fd_sc_hd__mux4_1 _39754_ (.A0(_01164_),
    .A1(_01165_),
    .A2(_01166_),
    .A3(_01167_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_01168_));
 sky130_fd_sc_hd__mux4_1 _39755_ (.A0(_01169_),
    .A1(_01170_),
    .A2(_01171_),
    .A3(_01172_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_01173_));
 sky130_fd_sc_hd__mux4_1 _39756_ (.A0(_01158_),
    .A1(_01163_),
    .A2(_01168_),
    .A3(_01173_),
    .S0(_00360_),
    .S1(_00362_),
    .X(_01174_));
 sky130_fd_sc_hd__mux4_1 _39757_ (.A0(_01148_),
    .A1(_01149_),
    .A2(_01150_),
    .A3(_01151_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_01152_));
 sky130_fd_sc_hd__mux4_1 _39758_ (.A0(_01127_),
    .A1(_01128_),
    .A2(_01129_),
    .A3(_01130_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_01131_));
 sky130_fd_sc_hd__mux4_1 _39759_ (.A0(_01132_),
    .A1(_01133_),
    .A2(_01134_),
    .A3(_01135_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_01136_));
 sky130_fd_sc_hd__mux4_1 _39760_ (.A0(_01137_),
    .A1(_01138_),
    .A2(_01139_),
    .A3(_01140_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_01141_));
 sky130_fd_sc_hd__mux4_1 _39761_ (.A0(_01142_),
    .A1(_01143_),
    .A2(_01144_),
    .A3(_01145_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_01146_));
 sky130_fd_sc_hd__mux4_1 _39762_ (.A0(_01131_),
    .A1(_01136_),
    .A2(_01141_),
    .A3(_01146_),
    .S0(_00360_),
    .S1(_00362_),
    .X(_01147_));
 sky130_fd_sc_hd__mux4_1 _39763_ (.A0(_01121_),
    .A1(_01122_),
    .A2(_01123_),
    .A3(_01124_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_01125_));
 sky130_fd_sc_hd__mux4_1 _39764_ (.A0(_01100_),
    .A1(_01101_),
    .A2(_01102_),
    .A3(_01103_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_01104_));
 sky130_fd_sc_hd__mux4_1 _39765_ (.A0(_01105_),
    .A1(_01106_),
    .A2(_01107_),
    .A3(_01108_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_01109_));
 sky130_fd_sc_hd__mux4_1 _39766_ (.A0(_01110_),
    .A1(_01111_),
    .A2(_01112_),
    .A3(_01113_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_01114_));
 sky130_fd_sc_hd__mux4_1 _39767_ (.A0(_01115_),
    .A1(_01116_),
    .A2(_01117_),
    .A3(_01118_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_01119_));
 sky130_fd_sc_hd__mux4_1 _39768_ (.A0(_01104_),
    .A1(_01109_),
    .A2(_01114_),
    .A3(_01119_),
    .S0(_00360_),
    .S1(_00362_),
    .X(_01120_));
 sky130_fd_sc_hd__mux4_1 _39769_ (.A0(_01094_),
    .A1(_01095_),
    .A2(_01096_),
    .A3(_01097_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_01098_));
 sky130_fd_sc_hd__mux4_1 _39770_ (.A0(_01073_),
    .A1(_01074_),
    .A2(_01075_),
    .A3(_01076_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_01077_));
 sky130_fd_sc_hd__mux4_1 _39771_ (.A0(_01078_),
    .A1(_01079_),
    .A2(_01080_),
    .A3(_01081_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_01082_));
 sky130_fd_sc_hd__mux4_1 _39772_ (.A0(_01083_),
    .A1(_01084_),
    .A2(_01085_),
    .A3(_01086_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_01087_));
 sky130_fd_sc_hd__mux4_1 _39773_ (.A0(_01088_),
    .A1(_01089_),
    .A2(_01090_),
    .A3(_01091_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_01092_));
 sky130_fd_sc_hd__mux4_1 _39774_ (.A0(_01077_),
    .A1(_01082_),
    .A2(_01087_),
    .A3(_01092_),
    .S0(_00360_),
    .S1(_00362_),
    .X(_01093_));
 sky130_fd_sc_hd__mux4_1 _39775_ (.A0(_01067_),
    .A1(_01068_),
    .A2(_01069_),
    .A3(_01070_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_01071_));
 sky130_fd_sc_hd__mux4_1 _39776_ (.A0(_01046_),
    .A1(_01047_),
    .A2(_01048_),
    .A3(_01049_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_01050_));
 sky130_fd_sc_hd__mux4_1 _39777_ (.A0(_01051_),
    .A1(_01052_),
    .A2(_01053_),
    .A3(_01054_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_01055_));
 sky130_fd_sc_hd__mux4_1 _39778_ (.A0(_01056_),
    .A1(_01057_),
    .A2(_01058_),
    .A3(_01059_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_01060_));
 sky130_fd_sc_hd__mux4_1 _39779_ (.A0(_01061_),
    .A1(_01062_),
    .A2(_01063_),
    .A3(_01064_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_01065_));
 sky130_fd_sc_hd__mux4_1 _39780_ (.A0(_01050_),
    .A1(_01055_),
    .A2(_01060_),
    .A3(_01065_),
    .S0(_00360_),
    .S1(_00362_),
    .X(_01066_));
 sky130_fd_sc_hd__mux4_1 _39781_ (.A0(_01040_),
    .A1(_01041_),
    .A2(_01042_),
    .A3(_01043_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_01044_));
 sky130_fd_sc_hd__mux4_1 _39782_ (.A0(_01019_),
    .A1(_01020_),
    .A2(_01021_),
    .A3(_01022_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_01023_));
 sky130_fd_sc_hd__mux4_1 _39783_ (.A0(_01024_),
    .A1(_01025_),
    .A2(_01026_),
    .A3(_01027_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_01028_));
 sky130_fd_sc_hd__mux4_1 _39784_ (.A0(_01029_),
    .A1(_01030_),
    .A2(_01031_),
    .A3(_01032_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_01033_));
 sky130_fd_sc_hd__mux4_1 _39785_ (.A0(_01034_),
    .A1(_01035_),
    .A2(_01036_),
    .A3(_01037_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_01038_));
 sky130_fd_sc_hd__mux4_1 _39786_ (.A0(_01023_),
    .A1(_01028_),
    .A2(_01033_),
    .A3(_01038_),
    .S0(_00360_),
    .S1(_00362_),
    .X(_01039_));
 sky130_fd_sc_hd__mux4_1 _39787_ (.A0(_01013_),
    .A1(_01014_),
    .A2(_01015_),
    .A3(_01016_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_01017_));
 sky130_fd_sc_hd__mux4_1 _39788_ (.A0(_00992_),
    .A1(_00993_),
    .A2(_00994_),
    .A3(_00995_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00996_));
 sky130_fd_sc_hd__mux4_1 _39789_ (.A0(_00997_),
    .A1(_00998_),
    .A2(_00999_),
    .A3(_01000_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_01001_));
 sky130_fd_sc_hd__mux4_1 _39790_ (.A0(_01002_),
    .A1(_01003_),
    .A2(_01004_),
    .A3(_01005_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_01006_));
 sky130_fd_sc_hd__mux4_1 _39791_ (.A0(_01007_),
    .A1(_01008_),
    .A2(_01009_),
    .A3(_01010_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_01011_));
 sky130_fd_sc_hd__mux4_1 _39792_ (.A0(_00996_),
    .A1(_01001_),
    .A2(_01006_),
    .A3(_01011_),
    .S0(_00360_),
    .S1(_00362_),
    .X(_01012_));
 sky130_fd_sc_hd__mux4_1 _39793_ (.A0(_00986_),
    .A1(_00987_),
    .A2(_00988_),
    .A3(_00989_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00990_));
 sky130_fd_sc_hd__mux4_1 _39794_ (.A0(_00965_),
    .A1(_00966_),
    .A2(_00967_),
    .A3(_00968_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00969_));
 sky130_fd_sc_hd__mux4_1 _39795_ (.A0(_00970_),
    .A1(_00971_),
    .A2(_00972_),
    .A3(_00973_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00974_));
 sky130_fd_sc_hd__mux4_1 _39796_ (.A0(_00975_),
    .A1(_00976_),
    .A2(_00977_),
    .A3(_00978_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00979_));
 sky130_fd_sc_hd__mux4_1 _39797_ (.A0(_00980_),
    .A1(_00981_),
    .A2(_00982_),
    .A3(_00983_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00984_));
 sky130_fd_sc_hd__mux4_1 _39798_ (.A0(_00969_),
    .A1(_00974_),
    .A2(_00979_),
    .A3(_00984_),
    .S0(_00360_),
    .S1(_00362_),
    .X(_00985_));
 sky130_fd_sc_hd__mux4_1 _39799_ (.A0(_00959_),
    .A1(_00960_),
    .A2(_00961_),
    .A3(_00962_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00963_));
 sky130_fd_sc_hd__mux4_1 _39800_ (.A0(_00938_),
    .A1(_00939_),
    .A2(_00940_),
    .A3(_00941_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00942_));
 sky130_fd_sc_hd__mux4_1 _39801_ (.A0(_00943_),
    .A1(_00944_),
    .A2(_00945_),
    .A3(_00946_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00947_));
 sky130_fd_sc_hd__mux4_1 _39802_ (.A0(_00948_),
    .A1(_00949_),
    .A2(_00950_),
    .A3(_00951_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00952_));
 sky130_fd_sc_hd__mux4_1 _39803_ (.A0(_00953_),
    .A1(_00954_),
    .A2(_00955_),
    .A3(_00956_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00957_));
 sky130_fd_sc_hd__mux4_1 _39804_ (.A0(_00942_),
    .A1(_00947_),
    .A2(_00952_),
    .A3(_00957_),
    .S0(_00360_),
    .S1(_00362_),
    .X(_00958_));
 sky130_fd_sc_hd__mux4_1 _39805_ (.A0(_00932_),
    .A1(_00933_),
    .A2(_00934_),
    .A3(_00935_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00936_));
 sky130_fd_sc_hd__mux4_1 _39806_ (.A0(_00911_),
    .A1(_00912_),
    .A2(_00913_),
    .A3(_00914_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00915_));
 sky130_fd_sc_hd__mux4_1 _39807_ (.A0(_00916_),
    .A1(_00917_),
    .A2(_00918_),
    .A3(_00919_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00920_));
 sky130_fd_sc_hd__mux4_1 _39808_ (.A0(_00921_),
    .A1(_00922_),
    .A2(_00923_),
    .A3(_00924_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00925_));
 sky130_fd_sc_hd__mux4_1 _39809_ (.A0(_00926_),
    .A1(_00927_),
    .A2(_00928_),
    .A3(_00929_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00930_));
 sky130_fd_sc_hd__mux4_1 _39810_ (.A0(_00915_),
    .A1(_00920_),
    .A2(_00925_),
    .A3(_00930_),
    .S0(_00360_),
    .S1(_00362_),
    .X(_00931_));
 sky130_fd_sc_hd__mux4_1 _39811_ (.A0(_00905_),
    .A1(_00906_),
    .A2(_00907_),
    .A3(_00908_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00909_));
 sky130_fd_sc_hd__mux4_1 _39812_ (.A0(_00884_),
    .A1(_00885_),
    .A2(_00886_),
    .A3(_00887_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00888_));
 sky130_fd_sc_hd__mux4_1 _39813_ (.A0(_00889_),
    .A1(_00890_),
    .A2(_00891_),
    .A3(_00892_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00893_));
 sky130_fd_sc_hd__mux4_1 _39814_ (.A0(_00894_),
    .A1(_00895_),
    .A2(_00896_),
    .A3(_00897_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00898_));
 sky130_fd_sc_hd__mux4_1 _39815_ (.A0(_00899_),
    .A1(_00900_),
    .A2(_00901_),
    .A3(_00902_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00903_));
 sky130_fd_sc_hd__mux4_1 _39816_ (.A0(_00888_),
    .A1(_00893_),
    .A2(_00898_),
    .A3(_00903_),
    .S0(_00360_),
    .S1(_00362_),
    .X(_00904_));
 sky130_fd_sc_hd__mux4_1 _39817_ (.A0(_00878_),
    .A1(_00879_),
    .A2(_00880_),
    .A3(_00881_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00882_));
 sky130_fd_sc_hd__mux4_1 _39818_ (.A0(_00857_),
    .A1(_00858_),
    .A2(_00859_),
    .A3(_00860_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00861_));
 sky130_fd_sc_hd__mux4_1 _39819_ (.A0(_00862_),
    .A1(_00863_),
    .A2(_00864_),
    .A3(_00865_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00866_));
 sky130_fd_sc_hd__mux4_1 _39820_ (.A0(_00867_),
    .A1(_00868_),
    .A2(_00869_),
    .A3(_00870_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00871_));
 sky130_fd_sc_hd__mux4_1 _39821_ (.A0(_00872_),
    .A1(_00873_),
    .A2(_00874_),
    .A3(_00875_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00876_));
 sky130_fd_sc_hd__mux4_1 _39822_ (.A0(_00861_),
    .A1(_00866_),
    .A2(_00871_),
    .A3(_00876_),
    .S0(_00360_),
    .S1(_00362_),
    .X(_00877_));
 sky130_fd_sc_hd__mux4_1 _39823_ (.A0(_00851_),
    .A1(_00852_),
    .A2(_00853_),
    .A3(_00854_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00855_));
 sky130_fd_sc_hd__mux4_1 _39824_ (.A0(_00830_),
    .A1(_00831_),
    .A2(_00832_),
    .A3(_00833_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00834_));
 sky130_fd_sc_hd__mux4_1 _39825_ (.A0(_00835_),
    .A1(_00836_),
    .A2(_00837_),
    .A3(_00838_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00839_));
 sky130_fd_sc_hd__mux4_1 _39826_ (.A0(_00840_),
    .A1(_00841_),
    .A2(_00842_),
    .A3(_00843_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00844_));
 sky130_fd_sc_hd__mux4_1 _39827_ (.A0(_00845_),
    .A1(_00846_),
    .A2(_00847_),
    .A3(_00848_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00849_));
 sky130_fd_sc_hd__mux4_1 _39828_ (.A0(_00834_),
    .A1(_00839_),
    .A2(_00844_),
    .A3(_00849_),
    .S0(_00360_),
    .S1(_00362_),
    .X(_00850_));
 sky130_fd_sc_hd__mux4_1 _39829_ (.A0(_00824_),
    .A1(_00825_),
    .A2(_00826_),
    .A3(_00827_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00828_));
 sky130_fd_sc_hd__mux4_1 _39830_ (.A0(_00803_),
    .A1(_00804_),
    .A2(_00805_),
    .A3(_00806_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00807_));
 sky130_fd_sc_hd__mux4_1 _39831_ (.A0(_00808_),
    .A1(_00809_),
    .A2(_00810_),
    .A3(_00811_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00812_));
 sky130_fd_sc_hd__mux4_1 _39832_ (.A0(_00813_),
    .A1(_00814_),
    .A2(_00815_),
    .A3(_00816_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00817_));
 sky130_fd_sc_hd__mux4_1 _39833_ (.A0(_00818_),
    .A1(_00819_),
    .A2(_00820_),
    .A3(_00821_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00822_));
 sky130_fd_sc_hd__mux4_1 _39834_ (.A0(_00807_),
    .A1(_00812_),
    .A2(_00817_),
    .A3(_00822_),
    .S0(_00360_),
    .S1(_00362_),
    .X(_00823_));
 sky130_fd_sc_hd__mux4_1 _39835_ (.A0(_00797_),
    .A1(_00798_),
    .A2(_00799_),
    .A3(_00800_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00801_));
 sky130_fd_sc_hd__mux4_1 _39836_ (.A0(_00776_),
    .A1(_00777_),
    .A2(_00778_),
    .A3(_00779_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00780_));
 sky130_fd_sc_hd__mux4_1 _39837_ (.A0(_00781_),
    .A1(_00782_),
    .A2(_00783_),
    .A3(_00784_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00785_));
 sky130_fd_sc_hd__mux4_1 _39838_ (.A0(_00786_),
    .A1(_00787_),
    .A2(_00788_),
    .A3(_00789_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00790_));
 sky130_fd_sc_hd__mux4_1 _39839_ (.A0(_00791_),
    .A1(_00792_),
    .A2(_00793_),
    .A3(_00794_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00795_));
 sky130_fd_sc_hd__mux4_1 _39840_ (.A0(_00780_),
    .A1(_00785_),
    .A2(_00790_),
    .A3(_00795_),
    .S0(_00360_),
    .S1(_00362_),
    .X(_00796_));
 sky130_fd_sc_hd__mux4_1 _39841_ (.A0(_00770_),
    .A1(_00771_),
    .A2(_00772_),
    .A3(_00773_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00774_));
 sky130_fd_sc_hd__mux4_1 _39842_ (.A0(_00749_),
    .A1(_00750_),
    .A2(_00751_),
    .A3(_00752_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00753_));
 sky130_fd_sc_hd__mux4_1 _39843_ (.A0(_00754_),
    .A1(_00755_),
    .A2(_00756_),
    .A3(_00757_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00758_));
 sky130_fd_sc_hd__mux4_1 _39844_ (.A0(_00759_),
    .A1(_00760_),
    .A2(_00761_),
    .A3(_00762_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00763_));
 sky130_fd_sc_hd__mux4_1 _39845_ (.A0(_00764_),
    .A1(_00765_),
    .A2(_00766_),
    .A3(_00767_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00768_));
 sky130_fd_sc_hd__mux4_1 _39846_ (.A0(_00753_),
    .A1(_00758_),
    .A2(_00763_),
    .A3(_00768_),
    .S0(_00360_),
    .S1(_00362_),
    .X(_00769_));
 sky130_fd_sc_hd__mux4_1 _39847_ (.A0(_00743_),
    .A1(_00744_),
    .A2(_00745_),
    .A3(_00746_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00747_));
 sky130_fd_sc_hd__mux4_1 _39848_ (.A0(_00722_),
    .A1(_00723_),
    .A2(_00724_),
    .A3(_00725_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00726_));
 sky130_fd_sc_hd__mux4_1 _39849_ (.A0(_00727_),
    .A1(_00728_),
    .A2(_00729_),
    .A3(_00730_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00731_));
 sky130_fd_sc_hd__mux4_1 _39850_ (.A0(_00732_),
    .A1(_00733_),
    .A2(_00734_),
    .A3(_00735_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00736_));
 sky130_fd_sc_hd__mux4_1 _39851_ (.A0(_00737_),
    .A1(_00738_),
    .A2(_00739_),
    .A3(_00740_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00741_));
 sky130_fd_sc_hd__mux4_1 _39852_ (.A0(_00726_),
    .A1(_00731_),
    .A2(_00736_),
    .A3(_00741_),
    .S0(_00360_),
    .S1(_00362_),
    .X(_00742_));
 sky130_fd_sc_hd__mux4_1 _39853_ (.A0(_00716_),
    .A1(_00717_),
    .A2(_00718_),
    .A3(_00719_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00720_));
 sky130_fd_sc_hd__mux4_1 _39854_ (.A0(_00695_),
    .A1(_00696_),
    .A2(_00697_),
    .A3(_00698_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00699_));
 sky130_fd_sc_hd__mux4_1 _39855_ (.A0(_00700_),
    .A1(_00701_),
    .A2(_00702_),
    .A3(_00703_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00704_));
 sky130_fd_sc_hd__mux4_1 _39856_ (.A0(_00705_),
    .A1(_00706_),
    .A2(_00707_),
    .A3(_00708_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00709_));
 sky130_fd_sc_hd__mux4_1 _39857_ (.A0(_00710_),
    .A1(_00711_),
    .A2(_00712_),
    .A3(_00713_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00714_));
 sky130_fd_sc_hd__mux4_1 _39858_ (.A0(_00699_),
    .A1(_00704_),
    .A2(_00709_),
    .A3(_00714_),
    .S0(_00360_),
    .S1(_00362_),
    .X(_00715_));
 sky130_fd_sc_hd__mux4_1 _39859_ (.A0(_00689_),
    .A1(_00690_),
    .A2(_00691_),
    .A3(_00692_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00693_));
 sky130_fd_sc_hd__mux4_1 _39860_ (.A0(_00668_),
    .A1(_00669_),
    .A2(_00670_),
    .A3(_00671_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00672_));
 sky130_fd_sc_hd__mux4_1 _39861_ (.A0(_00673_),
    .A1(_00674_),
    .A2(_00675_),
    .A3(_00676_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00677_));
 sky130_fd_sc_hd__mux4_1 _39862_ (.A0(_00678_),
    .A1(_00679_),
    .A2(_00680_),
    .A3(_00681_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00682_));
 sky130_fd_sc_hd__mux4_1 _39863_ (.A0(_00683_),
    .A1(_00684_),
    .A2(_00685_),
    .A3(_00686_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00687_));
 sky130_fd_sc_hd__mux4_1 _39864_ (.A0(_00672_),
    .A1(_00677_),
    .A2(_00682_),
    .A3(_00687_),
    .S0(_00360_),
    .S1(_00362_),
    .X(_00688_));
 sky130_fd_sc_hd__mux4_1 _39865_ (.A0(_00662_),
    .A1(_00663_),
    .A2(_00664_),
    .A3(_00665_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00666_));
 sky130_fd_sc_hd__mux4_1 _39866_ (.A0(_00641_),
    .A1(_00642_),
    .A2(_00643_),
    .A3(_00644_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00645_));
 sky130_fd_sc_hd__mux4_1 _39867_ (.A0(_00646_),
    .A1(_00647_),
    .A2(_00648_),
    .A3(_00649_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00650_));
 sky130_fd_sc_hd__mux4_1 _39868_ (.A0(_00651_),
    .A1(_00652_),
    .A2(_00653_),
    .A3(_00654_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00655_));
 sky130_fd_sc_hd__mux4_1 _39869_ (.A0(_00656_),
    .A1(_00657_),
    .A2(_00658_),
    .A3(_00659_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00660_));
 sky130_fd_sc_hd__mux4_1 _39870_ (.A0(_00645_),
    .A1(_00650_),
    .A2(_00655_),
    .A3(_00660_),
    .S0(_00360_),
    .S1(_00362_),
    .X(_00661_));
 sky130_fd_sc_hd__mux4_1 _39871_ (.A0(_00635_),
    .A1(_00636_),
    .A2(_00637_),
    .A3(_00638_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00639_));
 sky130_fd_sc_hd__mux4_1 _39872_ (.A0(_00614_),
    .A1(_00615_),
    .A2(_00616_),
    .A3(_00617_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00618_));
 sky130_fd_sc_hd__mux4_1 _39873_ (.A0(_00619_),
    .A1(_00620_),
    .A2(_00621_),
    .A3(_00622_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00623_));
 sky130_fd_sc_hd__mux4_1 _39874_ (.A0(_00624_),
    .A1(_00625_),
    .A2(_00626_),
    .A3(_00627_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00628_));
 sky130_fd_sc_hd__mux4_1 _39875_ (.A0(_00629_),
    .A1(_00630_),
    .A2(_00631_),
    .A3(_00632_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00633_));
 sky130_fd_sc_hd__mux4_1 _39876_ (.A0(_00618_),
    .A1(_00623_),
    .A2(_00628_),
    .A3(_00633_),
    .S0(_00360_),
    .S1(_00362_),
    .X(_00634_));
 sky130_fd_sc_hd__mux4_1 _39877_ (.A0(_00608_),
    .A1(_00609_),
    .A2(_00610_),
    .A3(_00611_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00612_));
 sky130_fd_sc_hd__mux4_1 _39878_ (.A0(_00587_),
    .A1(_00588_),
    .A2(_00589_),
    .A3(_00590_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00591_));
 sky130_fd_sc_hd__mux4_1 _39879_ (.A0(_00592_),
    .A1(_00593_),
    .A2(_00594_),
    .A3(_00595_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00596_));
 sky130_fd_sc_hd__mux4_1 _39880_ (.A0(_00597_),
    .A1(_00598_),
    .A2(_00599_),
    .A3(_00600_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00601_));
 sky130_fd_sc_hd__mux4_1 _39881_ (.A0(_00602_),
    .A1(_00603_),
    .A2(_00604_),
    .A3(_00605_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00606_));
 sky130_fd_sc_hd__mux4_1 _39882_ (.A0(_00591_),
    .A1(_00596_),
    .A2(_00601_),
    .A3(_00606_),
    .S0(_00360_),
    .S1(_00362_),
    .X(_00607_));
 sky130_fd_sc_hd__mux4_1 _39883_ (.A0(_00581_),
    .A1(_00582_),
    .A2(_00583_),
    .A3(_00584_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00585_));
 sky130_fd_sc_hd__mux4_1 _39884_ (.A0(_00560_),
    .A1(_00561_),
    .A2(_00562_),
    .A3(_00563_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00564_));
 sky130_fd_sc_hd__mux4_1 _39885_ (.A0(_00565_),
    .A1(_00566_),
    .A2(_00567_),
    .A3(_00568_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00569_));
 sky130_fd_sc_hd__mux4_1 _39886_ (.A0(_00570_),
    .A1(_00571_),
    .A2(_00572_),
    .A3(_00573_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00574_));
 sky130_fd_sc_hd__mux4_1 _39887_ (.A0(_00575_),
    .A1(_00576_),
    .A2(_00577_),
    .A3(_00578_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00579_));
 sky130_fd_sc_hd__mux4_1 _39888_ (.A0(_00564_),
    .A1(_00569_),
    .A2(_00574_),
    .A3(_00579_),
    .S0(_00360_),
    .S1(_00362_),
    .X(_00580_));
 sky130_fd_sc_hd__mux4_1 _39889_ (.A0(_00554_),
    .A1(_00555_),
    .A2(_00556_),
    .A3(_00557_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00558_));
 sky130_fd_sc_hd__mux4_1 _39890_ (.A0(_00533_),
    .A1(_00534_),
    .A2(_00535_),
    .A3(_00536_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00537_));
 sky130_fd_sc_hd__mux4_1 _39891_ (.A0(_00538_),
    .A1(_00539_),
    .A2(_00540_),
    .A3(_00541_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00542_));
 sky130_fd_sc_hd__mux4_1 _39892_ (.A0(_00543_),
    .A1(_00544_),
    .A2(_00545_),
    .A3(_00546_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00547_));
 sky130_fd_sc_hd__mux4_1 _39893_ (.A0(_00548_),
    .A1(_00549_),
    .A2(_00550_),
    .A3(_00551_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00552_));
 sky130_fd_sc_hd__mux4_1 _39894_ (.A0(_00537_),
    .A1(_00542_),
    .A2(_00547_),
    .A3(_00552_),
    .S0(_00360_),
    .S1(_00362_),
    .X(_00553_));
 sky130_fd_sc_hd__mux4_1 _39895_ (.A0(_00527_),
    .A1(_00528_),
    .A2(_00529_),
    .A3(_00530_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00531_));
 sky130_fd_sc_hd__mux4_1 _39896_ (.A0(_00506_),
    .A1(_00507_),
    .A2(_00508_),
    .A3(_00509_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00510_));
 sky130_fd_sc_hd__mux4_1 _39897_ (.A0(_00511_),
    .A1(_00512_),
    .A2(_00513_),
    .A3(_00514_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00515_));
 sky130_fd_sc_hd__mux4_1 _39898_ (.A0(_00516_),
    .A1(_00517_),
    .A2(_00518_),
    .A3(_00519_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00520_));
 sky130_fd_sc_hd__mux4_1 _39899_ (.A0(_00521_),
    .A1(_00522_),
    .A2(_00523_),
    .A3(_00524_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00525_));
 sky130_fd_sc_hd__mux4_1 _39900_ (.A0(_00510_),
    .A1(_00515_),
    .A2(_00520_),
    .A3(_00525_),
    .S0(_00360_),
    .S1(_00362_),
    .X(_00526_));
 sky130_fd_sc_hd__mux4_1 _39901_ (.A0(_00500_),
    .A1(_00501_),
    .A2(_00502_),
    .A3(_00503_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00504_));
 sky130_fd_sc_hd__mux4_1 _39902_ (.A0(_00479_),
    .A1(_00480_),
    .A2(_00481_),
    .A3(_00482_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00483_));
 sky130_fd_sc_hd__mux4_1 _39903_ (.A0(_00484_),
    .A1(_00485_),
    .A2(_00486_),
    .A3(_00487_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00488_));
 sky130_fd_sc_hd__mux4_1 _39904_ (.A0(_00489_),
    .A1(_00490_),
    .A2(_00491_),
    .A3(_00492_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00493_));
 sky130_fd_sc_hd__mux4_1 _39905_ (.A0(_00494_),
    .A1(_00495_),
    .A2(_00496_),
    .A3(_00497_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00498_));
 sky130_fd_sc_hd__mux4_1 _39906_ (.A0(_00483_),
    .A1(_00488_),
    .A2(_00493_),
    .A3(_00498_),
    .S0(_00360_),
    .S1(_00362_),
    .X(_00499_));
 sky130_fd_sc_hd__mux4_1 _39907_ (.A0(_00473_),
    .A1(_00474_),
    .A2(_00475_),
    .A3(_00476_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00477_));
 sky130_fd_sc_hd__mux4_1 _39908_ (.A0(_00452_),
    .A1(_00453_),
    .A2(_00454_),
    .A3(_00455_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00456_));
 sky130_fd_sc_hd__mux4_1 _39909_ (.A0(_00457_),
    .A1(_00458_),
    .A2(_00459_),
    .A3(_00460_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00461_));
 sky130_fd_sc_hd__mux4_1 _39910_ (.A0(_00462_),
    .A1(_00463_),
    .A2(_00464_),
    .A3(_00465_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00466_));
 sky130_fd_sc_hd__mux4_1 _39911_ (.A0(_00467_),
    .A1(_00468_),
    .A2(_00469_),
    .A3(_00470_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00471_));
 sky130_fd_sc_hd__mux4_1 _39912_ (.A0(_00456_),
    .A1(_00461_),
    .A2(_00466_),
    .A3(_00471_),
    .S0(_00360_),
    .S1(_00362_),
    .X(_00472_));
 sky130_fd_sc_hd__mux4_1 _39913_ (.A0(_00446_),
    .A1(_00447_),
    .A2(_00448_),
    .A3(_00449_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00450_));
 sky130_fd_sc_hd__mux4_1 _39914_ (.A0(_00425_),
    .A1(_00426_),
    .A2(_00427_),
    .A3(_00428_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00429_));
 sky130_fd_sc_hd__mux4_1 _39915_ (.A0(_00430_),
    .A1(_00431_),
    .A2(_00432_),
    .A3(_00433_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00434_));
 sky130_fd_sc_hd__mux4_1 _39916_ (.A0(_00435_),
    .A1(_00436_),
    .A2(_00437_),
    .A3(_00438_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00439_));
 sky130_fd_sc_hd__mux4_1 _39917_ (.A0(_00440_),
    .A1(_00441_),
    .A2(_00442_),
    .A3(_00443_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00444_));
 sky130_fd_sc_hd__mux4_1 _39918_ (.A0(_00429_),
    .A1(_00434_),
    .A2(_00439_),
    .A3(_00444_),
    .S0(_00360_),
    .S1(_00362_),
    .X(_00445_));
 sky130_fd_sc_hd__mux4_1 _39919_ (.A0(_00419_),
    .A1(_00420_),
    .A2(_00421_),
    .A3(_00422_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00423_));
 sky130_fd_sc_hd__mux4_1 _39920_ (.A0(_00398_),
    .A1(_00399_),
    .A2(_00400_),
    .A3(_00401_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00402_));
 sky130_fd_sc_hd__mux4_1 _39921_ (.A0(_00403_),
    .A1(_00404_),
    .A2(_00405_),
    .A3(_00406_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00407_));
 sky130_fd_sc_hd__mux4_1 _39922_ (.A0(_00408_),
    .A1(_00409_),
    .A2(_00410_),
    .A3(_00411_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00412_));
 sky130_fd_sc_hd__mux4_1 _39923_ (.A0(_00413_),
    .A1(_00414_),
    .A2(_00415_),
    .A3(_00416_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00417_));
 sky130_fd_sc_hd__mux4_1 _39924_ (.A0(_00402_),
    .A1(_00407_),
    .A2(_00412_),
    .A3(_00417_),
    .S0(_00360_),
    .S1(_00362_),
    .X(_00418_));
 sky130_fd_sc_hd__mux4_1 _39925_ (.A0(_00392_),
    .A1(_00393_),
    .A2(_00394_),
    .A3(_00395_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00396_));
 sky130_fd_sc_hd__mux4_1 _39926_ (.A0(_00371_),
    .A1(_00372_),
    .A2(_00373_),
    .A3(_00374_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00375_));
 sky130_fd_sc_hd__mux4_1 _39927_ (.A0(_00376_),
    .A1(_00377_),
    .A2(_00378_),
    .A3(_00379_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00380_));
 sky130_fd_sc_hd__mux4_1 _39928_ (.A0(_00381_),
    .A1(_00382_),
    .A2(_00383_),
    .A3(_00384_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00385_));
 sky130_fd_sc_hd__mux4_1 _39929_ (.A0(_00386_),
    .A1(_00387_),
    .A2(_00388_),
    .A3(_00389_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00390_));
 sky130_fd_sc_hd__mux4_1 _39930_ (.A0(_00375_),
    .A1(_00380_),
    .A2(_00385_),
    .A3(_00390_),
    .S0(_00360_),
    .S1(_00362_),
    .X(_00391_));
 sky130_fd_sc_hd__mux4_1 _39931_ (.A0(\cpuregs[16][0] ),
    .A1(\cpuregs[17][0] ),
    .A2(\cpuregs[18][0] ),
    .A3(\cpuregs[19][0] ),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00369_));
 sky130_fd_sc_hd__mux4_1 _39932_ (.A0(\cpuregs[0][0] ),
    .A1(\cpuregs[1][0] ),
    .A2(\cpuregs[2][0] ),
    .A3(\cpuregs[3][0] ),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00359_));
 sky130_fd_sc_hd__mux4_1 _39933_ (.A0(\cpuregs[4][0] ),
    .A1(\cpuregs[5][0] ),
    .A2(\cpuregs[6][0] ),
    .A3(\cpuregs[7][0] ),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00361_));
 sky130_fd_sc_hd__mux4_1 _39934_ (.A0(\cpuregs[8][0] ),
    .A1(\cpuregs[9][0] ),
    .A2(\cpuregs[10][0] ),
    .A3(\cpuregs[11][0] ),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00363_));
 sky130_fd_sc_hd__mux4_1 _39935_ (.A0(\cpuregs[12][0] ),
    .A1(\cpuregs[13][0] ),
    .A2(\cpuregs[14][0] ),
    .A3(\cpuregs[15][0] ),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00364_));
 sky130_fd_sc_hd__mux4_1 _39936_ (.A0(_00359_),
    .A1(_00361_),
    .A2(_00363_),
    .A3(_00364_),
    .S0(_00360_),
    .S1(_00362_),
    .X(_00365_));
 sky130_fd_sc_hd__mux4_1 _39937_ (.A0(_02581_),
    .A1(_01681_),
    .A2(_01679_),
    .A3(_02581_),
    .S0(_19782_),
    .S1(_00309_),
    .X(_01682_));
 sky130_fd_sc_hd__mux4_1 _39938_ (.A0(_02580_),
    .A1(_01677_),
    .A2(_01675_),
    .A3(_02580_),
    .S0(_19782_),
    .S1(_00309_),
    .X(_01678_));
 sky130_fd_sc_hd__mux4_1 _39939_ (.A0(_02579_),
    .A1(_01673_),
    .A2(_01671_),
    .A3(_02579_),
    .S0(_19782_),
    .S1(_00309_),
    .X(_01674_));
 sky130_fd_sc_hd__mux4_1 _39940_ (.A0(_02578_),
    .A1(_01669_),
    .A2(_01667_),
    .A3(_02578_),
    .S0(_19782_),
    .S1(_00309_),
    .X(_01670_));
 sky130_fd_sc_hd__mux4_1 _39941_ (.A0(_02577_),
    .A1(_01665_),
    .A2(_01663_),
    .A3(_02577_),
    .S0(_19782_),
    .S1(_00309_),
    .X(_01666_));
 sky130_fd_sc_hd__mux4_1 _39942_ (.A0(_02576_),
    .A1(_01661_),
    .A2(_01659_),
    .A3(_02576_),
    .S0(_19782_),
    .S1(_00309_),
    .X(_01662_));
 sky130_fd_sc_hd__mux4_1 _39943_ (.A0(_02575_),
    .A1(_01657_),
    .A2(_01655_),
    .A3(_02575_),
    .S0(_19782_),
    .S1(_00309_),
    .X(_01658_));
 sky130_fd_sc_hd__mux4_1 _39944_ (.A0(_02574_),
    .A1(_01653_),
    .A2(_01651_),
    .A3(_02574_),
    .S0(_19782_),
    .S1(_00309_),
    .X(_01654_));
 sky130_fd_sc_hd__mux4_1 _39945_ (.A0(_02573_),
    .A1(_01649_),
    .A2(_01647_),
    .A3(_02573_),
    .S0(_19782_),
    .S1(_00309_),
    .X(_01650_));
 sky130_fd_sc_hd__mux4_1 _39946_ (.A0(_02572_),
    .A1(_01645_),
    .A2(_01643_),
    .A3(_02572_),
    .S0(_19782_),
    .S1(_00309_),
    .X(_01646_));
 sky130_fd_sc_hd__mux4_1 _39947_ (.A0(_02570_),
    .A1(_01641_),
    .A2(_01639_),
    .A3(_02570_),
    .S0(_19782_),
    .S1(_00309_),
    .X(_01642_));
 sky130_fd_sc_hd__mux4_1 _39948_ (.A0(_02569_),
    .A1(_01637_),
    .A2(_01635_),
    .A3(_02569_),
    .S0(_19782_),
    .S1(_00309_),
    .X(_01638_));
 sky130_fd_sc_hd__mux4_1 _39949_ (.A0(_02568_),
    .A1(_01633_),
    .A2(_01631_),
    .A3(_02568_),
    .S0(_19782_),
    .S1(_00309_),
    .X(_01634_));
 sky130_fd_sc_hd__mux4_1 _39950_ (.A0(_02567_),
    .A1(_01629_),
    .A2(_01627_),
    .A3(_02567_),
    .S0(_19782_),
    .S1(_00309_),
    .X(_01630_));
 sky130_fd_sc_hd__mux4_1 _39951_ (.A0(_02566_),
    .A1(_01625_),
    .A2(_01623_),
    .A3(_02566_),
    .S0(_19782_),
    .S1(_00309_),
    .X(_01626_));
 sky130_fd_sc_hd__mux4_1 _39952_ (.A0(_02565_),
    .A1(_01621_),
    .A2(_01619_),
    .A3(_02565_),
    .S0(_19782_),
    .S1(_00309_),
    .X(_01622_));
 sky130_fd_sc_hd__mux4_1 _39953_ (.A0(_02564_),
    .A1(_01617_),
    .A2(_01615_),
    .A3(_02564_),
    .S0(_19782_),
    .S1(_00309_),
    .X(_01618_));
 sky130_fd_sc_hd__mux4_1 _39954_ (.A0(_02563_),
    .A1(_01613_),
    .A2(_01611_),
    .A3(_02563_),
    .S0(_19782_),
    .S1(_00309_),
    .X(_01614_));
 sky130_fd_sc_hd__mux4_1 _39955_ (.A0(_02562_),
    .A1(_01609_),
    .A2(_01607_),
    .A3(_02562_),
    .S0(_19782_),
    .S1(_00309_),
    .X(_01610_));
 sky130_fd_sc_hd__mux4_1 _39956_ (.A0(_02561_),
    .A1(_01605_),
    .A2(_01603_),
    .A3(_02561_),
    .S0(_19782_),
    .S1(_00309_),
    .X(_01606_));
 sky130_fd_sc_hd__mux4_1 _39957_ (.A0(_02589_),
    .A1(_01601_),
    .A2(_01599_),
    .A3(_02589_),
    .S0(_19782_),
    .S1(_00309_),
    .X(_01602_));
 sky130_fd_sc_hd__mux4_1 _39958_ (.A0(_02588_),
    .A1(_01597_),
    .A2(_01595_),
    .A3(_02588_),
    .S0(_19782_),
    .S1(_00309_),
    .X(_01598_));
 sky130_fd_sc_hd__mux4_1 _39959_ (.A0(_02587_),
    .A1(_01593_),
    .A2(_01591_),
    .A3(_02587_),
    .S0(_19782_),
    .S1(_00309_),
    .X(_01594_));
 sky130_fd_sc_hd__mux4_1 _39960_ (.A0(_02586_),
    .A1(_01589_),
    .A2(_01587_),
    .A3(_02586_),
    .S0(_19782_),
    .S1(_00309_),
    .X(_01590_));
 sky130_fd_sc_hd__mux4_1 _39961_ (.A0(_02585_),
    .A1(_01585_),
    .A2(_01583_),
    .A3(_02585_),
    .S0(_19782_),
    .S1(_00309_),
    .X(_01586_));
 sky130_fd_sc_hd__mux4_1 _39962_ (.A0(_02584_),
    .A1(_01581_),
    .A2(_01579_),
    .A3(_02584_),
    .S0(_19782_),
    .S1(_00309_),
    .X(_01582_));
 sky130_fd_sc_hd__mux4_1 _39963_ (.A0(_02583_),
    .A1(_01577_),
    .A2(_01575_),
    .A3(_02583_),
    .S0(_19782_),
    .S1(_00309_),
    .X(_01578_));
 sky130_fd_sc_hd__mux4_1 _39964_ (.A0(_02582_),
    .A1(_01573_),
    .A2(_01571_),
    .A3(_02582_),
    .S0(_19782_),
    .S1(_00309_),
    .X(_01574_));
 sky130_fd_sc_hd__mux4_1 _39965_ (.A0(_02571_),
    .A1(_01569_),
    .A2(_01567_),
    .A3(_02571_),
    .S0(_19782_),
    .S1(_00309_),
    .X(_01570_));
 sky130_fd_sc_hd__dfxtp_2 _39966_ (.CLK(clk),
    .D(_02687_),
    .Q(\alu_shl[0] ));
 sky130_fd_sc_hd__dfxtp_2 _39967_ (.CLK(clk),
    .D(_02688_),
    .Q(\alu_shl[1] ));
 sky130_fd_sc_hd__dfxtp_2 _39968_ (.CLK(clk),
    .D(_02689_),
    .Q(\alu_shl[2] ));
 sky130_fd_sc_hd__dfxtp_2 _39969_ (.CLK(clk),
    .D(_02690_),
    .Q(\alu_shl[3] ));
 sky130_fd_sc_hd__dfxtp_2 _39970_ (.CLK(clk),
    .D(_02691_),
    .Q(\alu_shl[4] ));
 sky130_fd_sc_hd__dfxtp_2 _39971_ (.CLK(clk),
    .D(_02692_),
    .Q(\alu_shl[5] ));
 sky130_fd_sc_hd__dfxtp_2 _39972_ (.CLK(clk),
    .D(_02693_),
    .Q(\alu_shl[6] ));
 sky130_fd_sc_hd__dfxtp_2 _39973_ (.CLK(clk),
    .D(_02694_),
    .Q(\alu_shl[7] ));
 sky130_fd_sc_hd__dfxtp_2 _39974_ (.CLK(clk),
    .D(_02695_),
    .Q(\alu_shl[8] ));
 sky130_fd_sc_hd__dfxtp_2 _39975_ (.CLK(clk),
    .D(_02696_),
    .Q(\alu_shl[9] ));
 sky130_fd_sc_hd__dfxtp_2 _39976_ (.CLK(clk),
    .D(_02697_),
    .Q(\alu_shl[10] ));
 sky130_fd_sc_hd__dfxtp_2 _39977_ (.CLK(clk),
    .D(_02698_),
    .Q(\alu_shl[11] ));
 sky130_fd_sc_hd__dfxtp_2 _39978_ (.CLK(clk),
    .D(_02699_),
    .Q(\alu_shl[12] ));
 sky130_fd_sc_hd__dfxtp_2 _39979_ (.CLK(clk),
    .D(_02700_),
    .Q(\alu_shl[13] ));
 sky130_fd_sc_hd__dfxtp_2 _39980_ (.CLK(clk),
    .D(_02701_),
    .Q(\alu_shl[14] ));
 sky130_fd_sc_hd__dfxtp_2 _39981_ (.CLK(clk),
    .D(_02702_),
    .Q(\alu_shl[15] ));
 sky130_fd_sc_hd__dfxtp_2 _39982_ (.CLK(clk),
    .D(_02703_),
    .Q(alu_wait));
 sky130_fd_sc_hd__dfxtp_2 _39983_ (.CLK(clk),
    .D(_02704_),
    .Q(\latched_rd[3] ));
 sky130_fd_sc_hd__dfxtp_2 _39984_ (.CLK(clk),
    .D(_02705_),
    .Q(\latched_rd[2] ));
 sky130_fd_sc_hd__dfxtp_2 _39985_ (.CLK(clk),
    .D(_02706_),
    .Q(\latched_rd[1] ));
 sky130_fd_sc_hd__dfxtp_2 _39986_ (.CLK(clk),
    .D(_02707_),
    .Q(\latched_rd[0] ));
 sky130_fd_sc_hd__dfxtp_2 _39987_ (.CLK(clk),
    .D(_02708_),
    .Q(\decoded_imm[31] ));
 sky130_fd_sc_hd__dfxtp_2 _39988_ (.CLK(clk),
    .D(_02709_),
    .Q(\decoded_imm[30] ));
 sky130_fd_sc_hd__dfxtp_2 _39989_ (.CLK(clk),
    .D(_02710_),
    .Q(\decoded_imm[29] ));
 sky130_fd_sc_hd__dfxtp_2 _39990_ (.CLK(clk),
    .D(_02711_),
    .Q(\decoded_imm[28] ));
 sky130_fd_sc_hd__dfxtp_2 _39991_ (.CLK(clk),
    .D(_02712_),
    .Q(\decoded_imm[27] ));
 sky130_fd_sc_hd__dfxtp_2 _39992_ (.CLK(clk),
    .D(_02713_),
    .Q(\decoded_imm[26] ));
 sky130_fd_sc_hd__dfxtp_2 _39993_ (.CLK(clk),
    .D(_02714_),
    .Q(\decoded_imm[25] ));
 sky130_fd_sc_hd__dfxtp_2 _39994_ (.CLK(clk),
    .D(_02715_),
    .Q(\decoded_imm[24] ));
 sky130_fd_sc_hd__dfxtp_2 _39995_ (.CLK(clk),
    .D(_02716_),
    .Q(\decoded_imm[23] ));
 sky130_fd_sc_hd__dfxtp_2 _39996_ (.CLK(clk),
    .D(_02717_),
    .Q(\decoded_imm[22] ));
 sky130_fd_sc_hd__dfxtp_2 _39997_ (.CLK(clk),
    .D(_02718_),
    .Q(\decoded_imm[21] ));
 sky130_fd_sc_hd__dfxtp_2 _39998_ (.CLK(clk),
    .D(_02719_),
    .Q(\decoded_imm[20] ));
 sky130_fd_sc_hd__dfxtp_2 _39999_ (.CLK(clk),
    .D(_02720_),
    .Q(\decoded_imm[19] ));
 sky130_fd_sc_hd__dfxtp_2 _40000_ (.CLK(clk),
    .D(_02721_),
    .Q(\decoded_imm[18] ));
 sky130_fd_sc_hd__dfxtp_2 _40001_ (.CLK(clk),
    .D(_02722_),
    .Q(\decoded_imm[17] ));
 sky130_fd_sc_hd__dfxtp_2 _40002_ (.CLK(clk),
    .D(_02723_),
    .Q(\decoded_imm[16] ));
 sky130_fd_sc_hd__dfxtp_2 _40003_ (.CLK(clk),
    .D(_02724_),
    .Q(\decoded_imm[15] ));
 sky130_fd_sc_hd__dfxtp_2 _40004_ (.CLK(clk),
    .D(_02725_),
    .Q(\decoded_imm[14] ));
 sky130_fd_sc_hd__dfxtp_2 _40005_ (.CLK(clk),
    .D(_02726_),
    .Q(\decoded_imm[13] ));
 sky130_fd_sc_hd__dfxtp_2 _40006_ (.CLK(clk),
    .D(_02727_),
    .Q(\decoded_imm[12] ));
 sky130_fd_sc_hd__dfxtp_2 _40007_ (.CLK(clk),
    .D(_02728_),
    .Q(\decoded_imm[11] ));
 sky130_fd_sc_hd__dfxtp_2 _40008_ (.CLK(clk),
    .D(_02729_),
    .Q(\decoded_imm[10] ));
 sky130_fd_sc_hd__dfxtp_2 _40009_ (.CLK(clk),
    .D(_02730_),
    .Q(\decoded_imm[9] ));
 sky130_fd_sc_hd__dfxtp_2 _40010_ (.CLK(clk),
    .D(_02731_),
    .Q(\decoded_imm[8] ));
 sky130_fd_sc_hd__dfxtp_2 _40011_ (.CLK(clk),
    .D(_02732_),
    .Q(\decoded_imm[7] ));
 sky130_fd_sc_hd__dfxtp_2 _40012_ (.CLK(clk),
    .D(_02733_),
    .Q(\decoded_imm[6] ));
 sky130_fd_sc_hd__dfxtp_2 _40013_ (.CLK(clk),
    .D(_02734_),
    .Q(\decoded_imm[5] ));
 sky130_fd_sc_hd__dfxtp_2 _40014_ (.CLK(clk),
    .D(_02735_),
    .Q(\decoded_imm[4] ));
 sky130_fd_sc_hd__dfxtp_2 _40015_ (.CLK(clk),
    .D(_02736_),
    .Q(\decoded_imm[3] ));
 sky130_fd_sc_hd__dfxtp_2 _40016_ (.CLK(clk),
    .D(_02737_),
    .Q(\decoded_imm[2] ));
 sky130_fd_sc_hd__dfxtp_2 _40017_ (.CLK(clk),
    .D(_02738_),
    .Q(\decoded_imm[1] ));
 sky130_fd_sc_hd__dfxtp_2 _40018_ (.CLK(clk),
    .D(_02739_),
    .Q(\irq_pending[31] ));
 sky130_fd_sc_hd__dfxtp_2 _40019_ (.CLK(clk),
    .D(_02740_),
    .Q(\irq_pending[30] ));
 sky130_fd_sc_hd__dfxtp_2 _40020_ (.CLK(clk),
    .D(_02741_),
    .Q(\irq_pending[29] ));
 sky130_fd_sc_hd__dfxtp_2 _40021_ (.CLK(clk),
    .D(_02742_),
    .Q(\irq_pending[28] ));
 sky130_fd_sc_hd__dfxtp_2 _40022_ (.CLK(clk),
    .D(_02743_),
    .Q(\irq_pending[27] ));
 sky130_fd_sc_hd__dfxtp_2 _40023_ (.CLK(clk),
    .D(_02744_),
    .Q(\irq_pending[26] ));
 sky130_fd_sc_hd__dfxtp_2 _40024_ (.CLK(clk),
    .D(_02745_),
    .Q(\irq_pending[25] ));
 sky130_fd_sc_hd__dfxtp_2 _40025_ (.CLK(clk),
    .D(_02746_),
    .Q(\irq_pending[24] ));
 sky130_fd_sc_hd__dfxtp_2 _40026_ (.CLK(clk),
    .D(_02747_),
    .Q(\irq_pending[23] ));
 sky130_fd_sc_hd__dfxtp_2 _40027_ (.CLK(clk),
    .D(_02748_),
    .Q(\irq_pending[22] ));
 sky130_fd_sc_hd__dfxtp_2 _40028_ (.CLK(clk),
    .D(_02749_),
    .Q(\irq_pending[21] ));
 sky130_fd_sc_hd__dfxtp_2 _40029_ (.CLK(clk),
    .D(_02750_),
    .Q(\irq_pending[20] ));
 sky130_fd_sc_hd__dfxtp_2 _40030_ (.CLK(clk),
    .D(_02751_),
    .Q(\irq_pending[19] ));
 sky130_fd_sc_hd__dfxtp_2 _40031_ (.CLK(clk),
    .D(_02752_),
    .Q(\irq_pending[18] ));
 sky130_fd_sc_hd__dfxtp_2 _40032_ (.CLK(clk),
    .D(_02753_),
    .Q(\irq_pending[17] ));
 sky130_fd_sc_hd__dfxtp_2 _40033_ (.CLK(clk),
    .D(_02754_),
    .Q(\irq_pending[16] ));
 sky130_fd_sc_hd__dfxtp_2 _40034_ (.CLK(clk),
    .D(_02755_),
    .Q(\irq_pending[15] ));
 sky130_fd_sc_hd__dfxtp_2 _40035_ (.CLK(clk),
    .D(_02756_),
    .Q(\irq_pending[14] ));
 sky130_fd_sc_hd__dfxtp_2 _40036_ (.CLK(clk),
    .D(_02757_),
    .Q(\irq_pending[13] ));
 sky130_fd_sc_hd__dfxtp_2 _40037_ (.CLK(clk),
    .D(_02758_),
    .Q(\irq_pending[12] ));
 sky130_fd_sc_hd__dfxtp_2 _40038_ (.CLK(clk),
    .D(_02759_),
    .Q(\irq_pending[11] ));
 sky130_fd_sc_hd__dfxtp_2 _40039_ (.CLK(clk),
    .D(_02760_),
    .Q(\irq_pending[10] ));
 sky130_fd_sc_hd__dfxtp_2 _40040_ (.CLK(clk),
    .D(_02761_),
    .Q(\irq_pending[9] ));
 sky130_fd_sc_hd__dfxtp_2 _40041_ (.CLK(clk),
    .D(_02762_),
    .Q(\irq_pending[8] ));
 sky130_fd_sc_hd__dfxtp_2 _40042_ (.CLK(clk),
    .D(_02763_),
    .Q(\irq_pending[7] ));
 sky130_fd_sc_hd__dfxtp_2 _40043_ (.CLK(clk),
    .D(_02764_),
    .Q(\irq_pending[6] ));
 sky130_fd_sc_hd__dfxtp_2 _40044_ (.CLK(clk),
    .D(_02765_),
    .Q(\irq_pending[5] ));
 sky130_fd_sc_hd__dfxtp_2 _40045_ (.CLK(clk),
    .D(_02766_),
    .Q(\irq_pending[4] ));
 sky130_fd_sc_hd__dfxtp_2 _40046_ (.CLK(clk),
    .D(_02767_),
    .Q(\irq_pending[3] ));
 sky130_fd_sc_hd__dfxtp_2 _40047_ (.CLK(clk),
    .D(_02768_),
    .Q(\irq_pending[1] ));
 sky130_fd_sc_hd__dfxtp_2 _40048_ (.CLK(clk),
    .D(_02769_),
    .Q(\irq_pending[0] ));
 sky130_fd_sc_hd__dfxtp_2 _40049_ (.CLK(clk),
    .D(_02770_),
    .Q(\reg_next_pc[0] ));
 sky130_fd_sc_hd__dfxtp_2 _40050_ (.CLK(clk),
    .D(_00045_),
    .Q(\mem_wordsize[0] ));
 sky130_fd_sc_hd__dfxtp_2 _40051_ (.CLK(clk),
    .D(_00046_),
    .Q(\mem_wordsize[1] ));
 sky130_fd_sc_hd__dfxtp_2 _40052_ (.CLK(clk),
    .D(_00047_),
    .Q(\mem_wordsize[2] ));
 sky130_fd_sc_hd__dfxtp_2 _40053_ (.CLK(clk),
    .D(_19784_),
    .Q(\reg_out[0] ));
 sky130_fd_sc_hd__dfxtp_2 _40054_ (.CLK(clk),
    .D(_19795_),
    .Q(\reg_out[1] ));
 sky130_fd_sc_hd__dfxtp_2 _40055_ (.CLK(clk),
    .D(_19806_),
    .Q(\reg_out[2] ));
 sky130_fd_sc_hd__dfxtp_2 _40056_ (.CLK(clk),
    .D(_19809_),
    .Q(\reg_out[3] ));
 sky130_fd_sc_hd__dfxtp_2 _40057_ (.CLK(clk),
    .D(_19810_),
    .Q(\reg_out[4] ));
 sky130_fd_sc_hd__dfxtp_2 _40058_ (.CLK(clk),
    .D(_19811_),
    .Q(\reg_out[5] ));
 sky130_fd_sc_hd__dfxtp_2 _40059_ (.CLK(clk),
    .D(_19812_),
    .Q(\reg_out[6] ));
 sky130_fd_sc_hd__dfxtp_2 _40060_ (.CLK(clk),
    .D(_19813_),
    .Q(\reg_out[7] ));
 sky130_fd_sc_hd__dfxtp_2 _40061_ (.CLK(clk),
    .D(_19814_),
    .Q(\reg_out[8] ));
 sky130_fd_sc_hd__dfxtp_2 _40062_ (.CLK(clk),
    .D(_19815_),
    .Q(\reg_out[9] ));
 sky130_fd_sc_hd__dfxtp_2 _40063_ (.CLK(clk),
    .D(_19785_),
    .Q(\reg_out[10] ));
 sky130_fd_sc_hd__dfxtp_2 _40064_ (.CLK(clk),
    .D(_19786_),
    .Q(\reg_out[11] ));
 sky130_fd_sc_hd__dfxtp_2 _40065_ (.CLK(clk),
    .D(_19787_),
    .Q(\reg_out[12] ));
 sky130_fd_sc_hd__dfxtp_2 _40066_ (.CLK(clk),
    .D(_19788_),
    .Q(\reg_out[13] ));
 sky130_fd_sc_hd__dfxtp_2 _40067_ (.CLK(clk),
    .D(_19789_),
    .Q(\reg_out[14] ));
 sky130_fd_sc_hd__dfxtp_2 _40068_ (.CLK(clk),
    .D(_19790_),
    .Q(\reg_out[15] ));
 sky130_fd_sc_hd__dfxtp_2 _40069_ (.CLK(clk),
    .D(_19791_),
    .Q(\reg_out[16] ));
 sky130_fd_sc_hd__dfxtp_2 _40070_ (.CLK(clk),
    .D(_19792_),
    .Q(\reg_out[17] ));
 sky130_fd_sc_hd__dfxtp_2 _40071_ (.CLK(clk),
    .D(_19793_),
    .Q(\reg_out[18] ));
 sky130_fd_sc_hd__dfxtp_2 _40072_ (.CLK(clk),
    .D(_19794_),
    .Q(\reg_out[19] ));
 sky130_fd_sc_hd__dfxtp_2 _40073_ (.CLK(clk),
    .D(_19796_),
    .Q(\reg_out[20] ));
 sky130_fd_sc_hd__dfxtp_2 _40074_ (.CLK(clk),
    .D(_19797_),
    .Q(\reg_out[21] ));
 sky130_fd_sc_hd__dfxtp_2 _40075_ (.CLK(clk),
    .D(_19798_),
    .Q(\reg_out[22] ));
 sky130_fd_sc_hd__dfxtp_2 _40076_ (.CLK(clk),
    .D(_19799_),
    .Q(\reg_out[23] ));
 sky130_fd_sc_hd__dfxtp_2 _40077_ (.CLK(clk),
    .D(_19800_),
    .Q(\reg_out[24] ));
 sky130_fd_sc_hd__dfxtp_2 _40078_ (.CLK(clk),
    .D(_19801_),
    .Q(\reg_out[25] ));
 sky130_fd_sc_hd__dfxtp_2 _40079_ (.CLK(clk),
    .D(_19802_),
    .Q(\reg_out[26] ));
 sky130_fd_sc_hd__dfxtp_2 _40080_ (.CLK(clk),
    .D(_19803_),
    .Q(\reg_out[27] ));
 sky130_fd_sc_hd__dfxtp_2 _40081_ (.CLK(clk),
    .D(_19804_),
    .Q(\reg_out[28] ));
 sky130_fd_sc_hd__dfxtp_2 _40082_ (.CLK(clk),
    .D(_19805_),
    .Q(\reg_out[29] ));
 sky130_fd_sc_hd__dfxtp_2 _40083_ (.CLK(clk),
    .D(_19807_),
    .Q(\reg_out[30] ));
 sky130_fd_sc_hd__dfxtp_2 _40084_ (.CLK(clk),
    .D(_19808_),
    .Q(\reg_out[31] ));
 sky130_fd_sc_hd__dfxtp_2 _40085_ (.CLK(clk),
    .D(_00004_),
    .Q(\irq_pending[2] ));
 sky130_fd_sc_hd__dfxtp_2 _40086_ (.CLK(clk),
    .D(_00003_),
    .Q(decoder_trigger));
 sky130_fd_sc_hd__dfxtp_2 _40087_ (.CLK(clk),
    .D(\alu_out[0] ),
    .Q(\alu_out_q[0] ));
 sky130_fd_sc_hd__dfxtp_2 _40088_ (.CLK(clk),
    .D(\alu_out[1] ),
    .Q(\alu_out_q[1] ));
 sky130_fd_sc_hd__dfxtp_2 _40089_ (.CLK(clk),
    .D(\alu_out[2] ),
    .Q(\alu_out_q[2] ));
 sky130_fd_sc_hd__dfxtp_2 _40090_ (.CLK(clk),
    .D(\alu_out[3] ),
    .Q(\alu_out_q[3] ));
 sky130_fd_sc_hd__dfxtp_2 _40091_ (.CLK(clk),
    .D(\alu_out[4] ),
    .Q(\alu_out_q[4] ));
 sky130_fd_sc_hd__dfxtp_2 _40092_ (.CLK(clk),
    .D(\alu_out[5] ),
    .Q(\alu_out_q[5] ));
 sky130_fd_sc_hd__dfxtp_2 _40093_ (.CLK(clk),
    .D(\alu_out[6] ),
    .Q(\alu_out_q[6] ));
 sky130_fd_sc_hd__dfxtp_2 _40094_ (.CLK(clk),
    .D(\alu_out[7] ),
    .Q(\alu_out_q[7] ));
 sky130_fd_sc_hd__dfxtp_2 _40095_ (.CLK(clk),
    .D(\alu_out[8] ),
    .Q(\alu_out_q[8] ));
 sky130_fd_sc_hd__dfxtp_2 _40096_ (.CLK(clk),
    .D(\alu_out[9] ),
    .Q(\alu_out_q[9] ));
 sky130_fd_sc_hd__dfxtp_2 _40097_ (.CLK(clk),
    .D(\alu_out[10] ),
    .Q(\alu_out_q[10] ));
 sky130_fd_sc_hd__dfxtp_2 _40098_ (.CLK(clk),
    .D(\alu_out[11] ),
    .Q(\alu_out_q[11] ));
 sky130_fd_sc_hd__dfxtp_2 _40099_ (.CLK(clk),
    .D(\alu_out[12] ),
    .Q(\alu_out_q[12] ));
 sky130_fd_sc_hd__dfxtp_2 _40100_ (.CLK(clk),
    .D(\alu_out[13] ),
    .Q(\alu_out_q[13] ));
 sky130_fd_sc_hd__dfxtp_2 _40101_ (.CLK(clk),
    .D(\alu_out[14] ),
    .Q(\alu_out_q[14] ));
 sky130_fd_sc_hd__dfxtp_2 _40102_ (.CLK(clk),
    .D(\alu_out[15] ),
    .Q(\alu_out_q[15] ));
 sky130_fd_sc_hd__dfxtp_2 _40103_ (.CLK(clk),
    .D(\alu_out[16] ),
    .Q(\alu_out_q[16] ));
 sky130_fd_sc_hd__dfxtp_2 _40104_ (.CLK(clk),
    .D(\alu_out[17] ),
    .Q(\alu_out_q[17] ));
 sky130_fd_sc_hd__dfxtp_2 _40105_ (.CLK(clk),
    .D(\alu_out[18] ),
    .Q(\alu_out_q[18] ));
 sky130_fd_sc_hd__dfxtp_2 _40106_ (.CLK(clk),
    .D(\alu_out[19] ),
    .Q(\alu_out_q[19] ));
 sky130_fd_sc_hd__dfxtp_2 _40107_ (.CLK(clk),
    .D(\alu_out[20] ),
    .Q(\alu_out_q[20] ));
 sky130_fd_sc_hd__dfxtp_2 _40108_ (.CLK(clk),
    .D(\alu_out[21] ),
    .Q(\alu_out_q[21] ));
 sky130_fd_sc_hd__dfxtp_2 _40109_ (.CLK(clk),
    .D(\alu_out[22] ),
    .Q(\alu_out_q[22] ));
 sky130_fd_sc_hd__dfxtp_2 _40110_ (.CLK(clk),
    .D(\alu_out[23] ),
    .Q(\alu_out_q[23] ));
 sky130_fd_sc_hd__dfxtp_2 _40111_ (.CLK(clk),
    .D(\alu_out[24] ),
    .Q(\alu_out_q[24] ));
 sky130_fd_sc_hd__dfxtp_2 _40112_ (.CLK(clk),
    .D(\alu_out[25] ),
    .Q(\alu_out_q[25] ));
 sky130_fd_sc_hd__dfxtp_2 _40113_ (.CLK(clk),
    .D(\alu_out[26] ),
    .Q(\alu_out_q[26] ));
 sky130_fd_sc_hd__dfxtp_2 _40114_ (.CLK(clk),
    .D(\alu_out[27] ),
    .Q(\alu_out_q[27] ));
 sky130_fd_sc_hd__dfxtp_2 _40115_ (.CLK(clk),
    .D(\alu_out[28] ),
    .Q(\alu_out_q[28] ));
 sky130_fd_sc_hd__dfxtp_2 _40116_ (.CLK(clk),
    .D(\alu_out[29] ),
    .Q(\alu_out_q[29] ));
 sky130_fd_sc_hd__dfxtp_2 _40117_ (.CLK(clk),
    .D(\alu_out[30] ),
    .Q(\alu_out_q[30] ));
 sky130_fd_sc_hd__dfxtp_2 _40118_ (.CLK(clk),
    .D(\alu_out[31] ),
    .Q(\alu_out_q[31] ));
 sky130_fd_sc_hd__dfxtp_2 _40119_ (.CLK(clk),
    .D(_00005_),
    .Q(is_lui_auipc_jal));
 sky130_fd_sc_hd__dfxtp_2 _40120_ (.CLK(clk),
    .D(_00006_),
    .Q(is_slti_blt_slt));
 sky130_fd_sc_hd__dfxtp_2 _40121_ (.CLK(clk),
    .D(_00007_),
    .Q(is_sltiu_bltu_sltu));
 sky130_fd_sc_hd__dfxtp_2 _40122_ (.CLK(clk),
    .D(_02591_),
    .Q(\alu_add_sub[0] ));
 sky130_fd_sc_hd__dfxtp_2 _40123_ (.CLK(clk),
    .D(_02602_),
    .Q(\alu_add_sub[1] ));
 sky130_fd_sc_hd__dfxtp_2 _40124_ (.CLK(clk),
    .D(_02613_),
    .Q(\alu_add_sub[2] ));
 sky130_fd_sc_hd__dfxtp_2 _40125_ (.CLK(clk),
    .D(_02616_),
    .Q(\alu_add_sub[3] ));
 sky130_fd_sc_hd__dfxtp_2 _40126_ (.CLK(clk),
    .D(_02617_),
    .Q(\alu_add_sub[4] ));
 sky130_fd_sc_hd__dfxtp_2 _40127_ (.CLK(clk),
    .D(_02618_),
    .Q(\alu_add_sub[5] ));
 sky130_fd_sc_hd__dfxtp_2 _40128_ (.CLK(clk),
    .D(_02619_),
    .Q(\alu_add_sub[6] ));
 sky130_fd_sc_hd__dfxtp_2 _40129_ (.CLK(clk),
    .D(_02620_),
    .Q(\alu_add_sub[7] ));
 sky130_fd_sc_hd__dfxtp_2 _40130_ (.CLK(clk),
    .D(_02621_),
    .Q(\alu_add_sub[8] ));
 sky130_fd_sc_hd__dfxtp_2 _40131_ (.CLK(clk),
    .D(_02622_),
    .Q(\alu_add_sub[9] ));
 sky130_fd_sc_hd__dfxtp_2 _40132_ (.CLK(clk),
    .D(_02592_),
    .Q(\alu_add_sub[10] ));
 sky130_fd_sc_hd__dfxtp_2 _40133_ (.CLK(clk),
    .D(_02593_),
    .Q(\alu_add_sub[11] ));
 sky130_fd_sc_hd__dfxtp_2 _40134_ (.CLK(clk),
    .D(_02594_),
    .Q(\alu_add_sub[12] ));
 sky130_fd_sc_hd__dfxtp_2 _40135_ (.CLK(clk),
    .D(_02595_),
    .Q(\alu_add_sub[13] ));
 sky130_fd_sc_hd__dfxtp_2 _40136_ (.CLK(clk),
    .D(_02596_),
    .Q(\alu_add_sub[14] ));
 sky130_fd_sc_hd__dfxtp_2 _40137_ (.CLK(clk),
    .D(_02597_),
    .Q(\alu_add_sub[15] ));
 sky130_fd_sc_hd__dfxtp_2 _40138_ (.CLK(clk),
    .D(_02598_),
    .Q(\alu_add_sub[16] ));
 sky130_fd_sc_hd__dfxtp_2 _40139_ (.CLK(clk),
    .D(_02599_),
    .Q(\alu_add_sub[17] ));
 sky130_fd_sc_hd__dfxtp_2 _40140_ (.CLK(clk),
    .D(_02600_),
    .Q(\alu_add_sub[18] ));
 sky130_fd_sc_hd__dfxtp_2 _40141_ (.CLK(clk),
    .D(_02601_),
    .Q(\alu_add_sub[19] ));
 sky130_fd_sc_hd__dfxtp_2 _40142_ (.CLK(clk),
    .D(_02603_),
    .Q(\alu_add_sub[20] ));
 sky130_fd_sc_hd__dfxtp_2 _40143_ (.CLK(clk),
    .D(_02604_),
    .Q(\alu_add_sub[21] ));
 sky130_fd_sc_hd__dfxtp_2 _40144_ (.CLK(clk),
    .D(_02605_),
    .Q(\alu_add_sub[22] ));
 sky130_fd_sc_hd__dfxtp_2 _40145_ (.CLK(clk),
    .D(_02606_),
    .Q(\alu_add_sub[23] ));
 sky130_fd_sc_hd__dfxtp_2 _40146_ (.CLK(clk),
    .D(_02607_),
    .Q(\alu_add_sub[24] ));
 sky130_fd_sc_hd__dfxtp_2 _40147_ (.CLK(clk),
    .D(_02608_),
    .Q(\alu_add_sub[25] ));
 sky130_fd_sc_hd__dfxtp_2 _40148_ (.CLK(clk),
    .D(_02609_),
    .Q(\alu_add_sub[26] ));
 sky130_fd_sc_hd__dfxtp_2 _40149_ (.CLK(clk),
    .D(_02610_),
    .Q(\alu_add_sub[27] ));
 sky130_fd_sc_hd__dfxtp_2 _40150_ (.CLK(clk),
    .D(_02611_),
    .Q(\alu_add_sub[28] ));
 sky130_fd_sc_hd__dfxtp_2 _40151_ (.CLK(clk),
    .D(_02612_),
    .Q(\alu_add_sub[29] ));
 sky130_fd_sc_hd__dfxtp_2 _40152_ (.CLK(clk),
    .D(_02614_),
    .Q(\alu_add_sub[30] ));
 sky130_fd_sc_hd__dfxtp_2 _40153_ (.CLK(clk),
    .D(_02615_),
    .Q(\alu_add_sub[31] ));
 sky130_fd_sc_hd__dfxtp_2 _40154_ (.CLK(clk),
    .D(_19819_),
    .Q(\alu_shl[16] ));
 sky130_fd_sc_hd__dfxtp_2 _40155_ (.CLK(clk),
    .D(_19820_),
    .Q(\alu_shl[17] ));
 sky130_fd_sc_hd__dfxtp_2 _40156_ (.CLK(clk),
    .D(_19821_),
    .Q(\alu_shl[18] ));
 sky130_fd_sc_hd__dfxtp_2 _40157_ (.CLK(clk),
    .D(_19822_),
    .Q(\alu_shl[19] ));
 sky130_fd_sc_hd__dfxtp_2 _40158_ (.CLK(clk),
    .D(_19823_),
    .Q(\alu_shl[20] ));
 sky130_fd_sc_hd__dfxtp_2 _40159_ (.CLK(clk),
    .D(_19824_),
    .Q(\alu_shl[21] ));
 sky130_fd_sc_hd__dfxtp_2 _40160_ (.CLK(clk),
    .D(_19825_),
    .Q(\alu_shl[22] ));
 sky130_fd_sc_hd__dfxtp_2 _40161_ (.CLK(clk),
    .D(_19826_),
    .Q(\alu_shl[23] ));
 sky130_fd_sc_hd__dfxtp_2 _40162_ (.CLK(clk),
    .D(_19827_),
    .Q(\alu_shl[24] ));
 sky130_fd_sc_hd__dfxtp_2 _40163_ (.CLK(clk),
    .D(_19828_),
    .Q(\alu_shl[25] ));
 sky130_fd_sc_hd__dfxtp_2 _40164_ (.CLK(clk),
    .D(_19829_),
    .Q(\alu_shl[26] ));
 sky130_fd_sc_hd__dfxtp_2 _40165_ (.CLK(clk),
    .D(_19830_),
    .Q(\alu_shl[27] ));
 sky130_fd_sc_hd__dfxtp_2 _40166_ (.CLK(clk),
    .D(_19831_),
    .Q(\alu_shl[28] ));
 sky130_fd_sc_hd__dfxtp_2 _40167_ (.CLK(clk),
    .D(_19832_),
    .Q(\alu_shl[29] ));
 sky130_fd_sc_hd__dfxtp_2 _40168_ (.CLK(clk),
    .D(_19833_),
    .Q(\alu_shl[30] ));
 sky130_fd_sc_hd__dfxtp_2 _40169_ (.CLK(clk),
    .D(_19834_),
    .Q(\alu_shl[31] ));
 sky130_fd_sc_hd__dfxtp_2 _40170_ (.CLK(clk),
    .D(_19835_),
    .Q(\alu_shr[0] ));
 sky130_fd_sc_hd__dfxtp_2 _40171_ (.CLK(clk),
    .D(_19846_),
    .Q(\alu_shr[1] ));
 sky130_fd_sc_hd__dfxtp_2 _40172_ (.CLK(clk),
    .D(_19857_),
    .Q(\alu_shr[2] ));
 sky130_fd_sc_hd__dfxtp_2 _40173_ (.CLK(clk),
    .D(_19860_),
    .Q(\alu_shr[3] ));
 sky130_fd_sc_hd__dfxtp_2 _40174_ (.CLK(clk),
    .D(_19861_),
    .Q(\alu_shr[4] ));
 sky130_fd_sc_hd__dfxtp_2 _40175_ (.CLK(clk),
    .D(_19862_),
    .Q(\alu_shr[5] ));
 sky130_fd_sc_hd__dfxtp_2 _40176_ (.CLK(clk),
    .D(_19863_),
    .Q(\alu_shr[6] ));
 sky130_fd_sc_hd__dfxtp_2 _40177_ (.CLK(clk),
    .D(_19864_),
    .Q(\alu_shr[7] ));
 sky130_fd_sc_hd__dfxtp_2 _40178_ (.CLK(clk),
    .D(_19865_),
    .Q(\alu_shr[8] ));
 sky130_fd_sc_hd__dfxtp_2 _40179_ (.CLK(clk),
    .D(_19866_),
    .Q(\alu_shr[9] ));
 sky130_fd_sc_hd__dfxtp_2 _40180_ (.CLK(clk),
    .D(_19836_),
    .Q(\alu_shr[10] ));
 sky130_fd_sc_hd__dfxtp_2 _40181_ (.CLK(clk),
    .D(_19837_),
    .Q(\alu_shr[11] ));
 sky130_fd_sc_hd__dfxtp_2 _40182_ (.CLK(clk),
    .D(_19838_),
    .Q(\alu_shr[12] ));
 sky130_fd_sc_hd__dfxtp_2 _40183_ (.CLK(clk),
    .D(_19839_),
    .Q(\alu_shr[13] ));
 sky130_fd_sc_hd__dfxtp_2 _40184_ (.CLK(clk),
    .D(_19840_),
    .Q(\alu_shr[14] ));
 sky130_fd_sc_hd__dfxtp_2 _40185_ (.CLK(clk),
    .D(_19841_),
    .Q(\alu_shr[15] ));
 sky130_fd_sc_hd__dfxtp_2 _40186_ (.CLK(clk),
    .D(_19842_),
    .Q(\alu_shr[16] ));
 sky130_fd_sc_hd__dfxtp_2 _40187_ (.CLK(clk),
    .D(_19843_),
    .Q(\alu_shr[17] ));
 sky130_fd_sc_hd__dfxtp_2 _40188_ (.CLK(clk),
    .D(_19844_),
    .Q(\alu_shr[18] ));
 sky130_fd_sc_hd__dfxtp_2 _40189_ (.CLK(clk),
    .D(_19845_),
    .Q(\alu_shr[19] ));
 sky130_fd_sc_hd__dfxtp_2 _40190_ (.CLK(clk),
    .D(_19847_),
    .Q(\alu_shr[20] ));
 sky130_fd_sc_hd__dfxtp_2 _40191_ (.CLK(clk),
    .D(_19848_),
    .Q(\alu_shr[21] ));
 sky130_fd_sc_hd__dfxtp_2 _40192_ (.CLK(clk),
    .D(_19849_),
    .Q(\alu_shr[22] ));
 sky130_fd_sc_hd__dfxtp_2 _40193_ (.CLK(clk),
    .D(_19850_),
    .Q(\alu_shr[23] ));
 sky130_fd_sc_hd__dfxtp_2 _40194_ (.CLK(clk),
    .D(_19851_),
    .Q(\alu_shr[24] ));
 sky130_fd_sc_hd__dfxtp_2 _40195_ (.CLK(clk),
    .D(_19852_),
    .Q(\alu_shr[25] ));
 sky130_fd_sc_hd__dfxtp_2 _40196_ (.CLK(clk),
    .D(_19853_),
    .Q(\alu_shr[26] ));
 sky130_fd_sc_hd__dfxtp_2 _40197_ (.CLK(clk),
    .D(_19854_),
    .Q(\alu_shr[27] ));
 sky130_fd_sc_hd__dfxtp_2 _40198_ (.CLK(clk),
    .D(_19855_),
    .Q(\alu_shr[28] ));
 sky130_fd_sc_hd__dfxtp_2 _40199_ (.CLK(clk),
    .D(_19856_),
    .Q(\alu_shr[29] ));
 sky130_fd_sc_hd__dfxtp_2 _40200_ (.CLK(clk),
    .D(_19858_),
    .Q(\alu_shr[30] ));
 sky130_fd_sc_hd__dfxtp_2 _40201_ (.CLK(clk),
    .D(_19859_),
    .Q(\alu_shr[31] ));
 sky130_fd_sc_hd__dfxtp_2 _40202_ (.CLK(clk),
    .D(_00000_),
    .Q(alu_eq));
 sky130_fd_sc_hd__dfxtp_2 _40203_ (.CLK(clk),
    .D(_00002_),
    .Q(alu_ltu));
 sky130_fd_sc_hd__dfxtp_2 _40204_ (.CLK(clk),
    .D(_00001_),
    .Q(alu_lts));
 sky130_fd_sc_hd__dfxtp_2 _40205_ (.CLK(clk),
    .D(_02623_),
    .Q(\pcpi_mul.rd[0] ));
 sky130_fd_sc_hd__dfxtp_2 _40206_ (.CLK(clk),
    .D(_02624_),
    .Q(\pcpi_mul.rd[1] ));
 sky130_fd_sc_hd__dfxtp_2 _40207_ (.CLK(clk),
    .D(_02625_),
    .Q(\pcpi_mul.rd[2] ));
 sky130_fd_sc_hd__dfxtp_2 _40208_ (.CLK(clk),
    .D(_02626_),
    .Q(\pcpi_mul.rd[3] ));
 sky130_fd_sc_hd__dfxtp_2 _40209_ (.CLK(clk),
    .D(_02627_),
    .Q(\pcpi_mul.rd[4] ));
 sky130_fd_sc_hd__dfxtp_2 _40210_ (.CLK(clk),
    .D(_02628_),
    .Q(\pcpi_mul.rd[5] ));
 sky130_fd_sc_hd__dfxtp_2 _40211_ (.CLK(clk),
    .D(_02683_),
    .Q(\pcpi_mul.rd[6] ));
 sky130_fd_sc_hd__dfxtp_2 _40212_ (.CLK(clk),
    .D(_02684_),
    .Q(\pcpi_mul.rd[7] ));
 sky130_fd_sc_hd__dfxtp_2 _40213_ (.CLK(clk),
    .D(_02685_),
    .Q(\pcpi_mul.rd[8] ));
 sky130_fd_sc_hd__dfxtp_2 _40214_ (.CLK(clk),
    .D(_02686_),
    .Q(\pcpi_mul.rd[9] ));
 sky130_fd_sc_hd__dfxtp_2 _40215_ (.CLK(clk),
    .D(_02629_),
    .Q(\pcpi_mul.rd[10] ));
 sky130_fd_sc_hd__dfxtp_2 _40216_ (.CLK(clk),
    .D(_02630_),
    .Q(\pcpi_mul.rd[11] ));
 sky130_fd_sc_hd__dfxtp_2 _40217_ (.CLK(clk),
    .D(_02631_),
    .Q(\pcpi_mul.rd[12] ));
 sky130_fd_sc_hd__dfxtp_2 _40218_ (.CLK(clk),
    .D(_02632_),
    .Q(\pcpi_mul.rd[13] ));
 sky130_fd_sc_hd__dfxtp_2 _40219_ (.CLK(clk),
    .D(_02633_),
    .Q(\pcpi_mul.rd[14] ));
 sky130_fd_sc_hd__dfxtp_2 _40220_ (.CLK(clk),
    .D(_02634_),
    .Q(\pcpi_mul.rd[15] ));
 sky130_fd_sc_hd__dfxtp_2 _40221_ (.CLK(clk),
    .D(_02635_),
    .Q(\pcpi_mul.rd[16] ));
 sky130_fd_sc_hd__dfxtp_2 _40222_ (.CLK(clk),
    .D(_02636_),
    .Q(\pcpi_mul.rd[17] ));
 sky130_fd_sc_hd__dfxtp_2 _40223_ (.CLK(clk),
    .D(_02637_),
    .Q(\pcpi_mul.rd[18] ));
 sky130_fd_sc_hd__dfxtp_2 _40224_ (.CLK(clk),
    .D(_02638_),
    .Q(\pcpi_mul.rd[19] ));
 sky130_fd_sc_hd__dfxtp_2 _40225_ (.CLK(clk),
    .D(_02639_),
    .Q(\pcpi_mul.rd[20] ));
 sky130_fd_sc_hd__dfxtp_2 _40226_ (.CLK(clk),
    .D(_02640_),
    .Q(\pcpi_mul.rd[21] ));
 sky130_fd_sc_hd__dfxtp_2 _40227_ (.CLK(clk),
    .D(_02641_),
    .Q(\pcpi_mul.rd[22] ));
 sky130_fd_sc_hd__dfxtp_2 _40228_ (.CLK(clk),
    .D(_02642_),
    .Q(\pcpi_mul.rd[23] ));
 sky130_fd_sc_hd__dfxtp_2 _40229_ (.CLK(clk),
    .D(_02643_),
    .Q(\pcpi_mul.rd[24] ));
 sky130_fd_sc_hd__dfxtp_2 _40230_ (.CLK(clk),
    .D(_02644_),
    .Q(\pcpi_mul.rd[25] ));
 sky130_fd_sc_hd__dfxtp_2 _40231_ (.CLK(clk),
    .D(_02645_),
    .Q(\pcpi_mul.rd[26] ));
 sky130_fd_sc_hd__dfxtp_2 _40232_ (.CLK(clk),
    .D(_02646_),
    .Q(\pcpi_mul.rd[27] ));
 sky130_fd_sc_hd__dfxtp_2 _40233_ (.CLK(clk),
    .D(_02647_),
    .Q(\pcpi_mul.rd[28] ));
 sky130_fd_sc_hd__dfxtp_2 _40234_ (.CLK(clk),
    .D(_02648_),
    .Q(\pcpi_mul.rd[29] ));
 sky130_fd_sc_hd__dfxtp_2 _40235_ (.CLK(clk),
    .D(_02649_),
    .Q(\pcpi_mul.rd[30] ));
 sky130_fd_sc_hd__dfxtp_2 _40236_ (.CLK(clk),
    .D(_02650_),
    .Q(\pcpi_mul.rd[31] ));
 sky130_fd_sc_hd__dfxtp_2 _40237_ (.CLK(clk),
    .D(_02651_),
    .Q(\pcpi_mul.rd[32] ));
 sky130_fd_sc_hd__dfxtp_2 _40238_ (.CLK(clk),
    .D(_02652_),
    .Q(\pcpi_mul.rd[33] ));
 sky130_fd_sc_hd__dfxtp_2 _40239_ (.CLK(clk),
    .D(_02653_),
    .Q(\pcpi_mul.rd[34] ));
 sky130_fd_sc_hd__dfxtp_2 _40240_ (.CLK(clk),
    .D(_02654_),
    .Q(\pcpi_mul.rd[35] ));
 sky130_fd_sc_hd__dfxtp_2 _40241_ (.CLK(clk),
    .D(_02655_),
    .Q(\pcpi_mul.rd[36] ));
 sky130_fd_sc_hd__dfxtp_2 _40242_ (.CLK(clk),
    .D(_02656_),
    .Q(\pcpi_mul.rd[37] ));
 sky130_fd_sc_hd__dfxtp_2 _40243_ (.CLK(clk),
    .D(_02657_),
    .Q(\pcpi_mul.rd[38] ));
 sky130_fd_sc_hd__dfxtp_2 _40244_ (.CLK(clk),
    .D(_02658_),
    .Q(\pcpi_mul.rd[39] ));
 sky130_fd_sc_hd__dfxtp_2 _40245_ (.CLK(clk),
    .D(_02659_),
    .Q(\pcpi_mul.rd[40] ));
 sky130_fd_sc_hd__dfxtp_2 _40246_ (.CLK(clk),
    .D(_02660_),
    .Q(\pcpi_mul.rd[41] ));
 sky130_fd_sc_hd__dfxtp_2 _40247_ (.CLK(clk),
    .D(_02661_),
    .Q(\pcpi_mul.rd[42] ));
 sky130_fd_sc_hd__dfxtp_2 _40248_ (.CLK(clk),
    .D(_02662_),
    .Q(\pcpi_mul.rd[43] ));
 sky130_fd_sc_hd__dfxtp_2 _40249_ (.CLK(clk),
    .D(_02663_),
    .Q(\pcpi_mul.rd[44] ));
 sky130_fd_sc_hd__dfxtp_2 _40250_ (.CLK(clk),
    .D(_02664_),
    .Q(\pcpi_mul.rd[45] ));
 sky130_fd_sc_hd__dfxtp_2 _40251_ (.CLK(clk),
    .D(_02665_),
    .Q(\pcpi_mul.rd[46] ));
 sky130_fd_sc_hd__dfxtp_2 _40252_ (.CLK(clk),
    .D(_02666_),
    .Q(\pcpi_mul.rd[47] ));
 sky130_fd_sc_hd__dfxtp_2 _40253_ (.CLK(clk),
    .D(_02667_),
    .Q(\pcpi_mul.rd[48] ));
 sky130_fd_sc_hd__dfxtp_2 _40254_ (.CLK(clk),
    .D(_02668_),
    .Q(\pcpi_mul.rd[49] ));
 sky130_fd_sc_hd__dfxtp_2 _40255_ (.CLK(clk),
    .D(_02669_),
    .Q(\pcpi_mul.rd[50] ));
 sky130_fd_sc_hd__dfxtp_2 _40256_ (.CLK(clk),
    .D(_02670_),
    .Q(\pcpi_mul.rd[51] ));
 sky130_fd_sc_hd__dfxtp_2 _40257_ (.CLK(clk),
    .D(_02671_),
    .Q(\pcpi_mul.rd[52] ));
 sky130_fd_sc_hd__dfxtp_2 _40258_ (.CLK(clk),
    .D(_02672_),
    .Q(\pcpi_mul.rd[53] ));
 sky130_fd_sc_hd__dfxtp_2 _40259_ (.CLK(clk),
    .D(_02673_),
    .Q(\pcpi_mul.rd[54] ));
 sky130_fd_sc_hd__dfxtp_2 _40260_ (.CLK(clk),
    .D(_02674_),
    .Q(\pcpi_mul.rd[55] ));
 sky130_fd_sc_hd__dfxtp_2 _40261_ (.CLK(clk),
    .D(_02675_),
    .Q(\pcpi_mul.rd[56] ));
 sky130_fd_sc_hd__dfxtp_2 _40262_ (.CLK(clk),
    .D(_02676_),
    .Q(\pcpi_mul.rd[57] ));
 sky130_fd_sc_hd__dfxtp_2 _40263_ (.CLK(clk),
    .D(_02677_),
    .Q(\pcpi_mul.rd[58] ));
 sky130_fd_sc_hd__dfxtp_2 _40264_ (.CLK(clk),
    .D(_02678_),
    .Q(\pcpi_mul.rd[59] ));
 sky130_fd_sc_hd__dfxtp_2 _40265_ (.CLK(clk),
    .D(_02679_),
    .Q(\pcpi_mul.rd[60] ));
 sky130_fd_sc_hd__dfxtp_2 _40266_ (.CLK(clk),
    .D(_02680_),
    .Q(\pcpi_mul.rd[61] ));
 sky130_fd_sc_hd__dfxtp_2 _40267_ (.CLK(clk),
    .D(_02681_),
    .Q(\pcpi_mul.rd[62] ));
 sky130_fd_sc_hd__dfxtp_2 _40268_ (.CLK(clk),
    .D(_02682_),
    .Q(\pcpi_mul.rd[63] ));
 sky130_fd_sc_hd__dfxtp_2 _40269_ (.CLK(clk),
    .D(\pcpi_mul.instr_any_mulh ),
    .Q(\pcpi_mul.shift_out ));
 sky130_fd_sc_hd__dfxtp_2 _40270_ (.CLK(clk),
    .D(_00038_),
    .Q(\cpu_state[0] ));
 sky130_fd_sc_hd__dfxtp_2 _40271_ (.CLK(clk),
    .D(_00039_),
    .Q(\cpu_state[1] ));
 sky130_fd_sc_hd__dfxtp_2 _40272_ (.CLK(clk),
    .D(_00040_),
    .Q(\cpu_state[2] ));
 sky130_fd_sc_hd__dfxtp_2 _40273_ (.CLK(clk),
    .D(_00041_),
    .Q(\cpu_state[3] ));
 sky130_fd_sc_hd__dfxtp_2 _40274_ (.CLK(clk),
    .D(_00042_),
    .Q(\cpu_state[4] ));
 sky130_fd_sc_hd__dfxtp_2 _40275_ (.CLK(clk),
    .D(_00043_),
    .Q(\cpu_state[5] ));
 sky130_fd_sc_hd__dfxtp_2 _40276_ (.CLK(clk),
    .D(_00044_),
    .Q(\cpu_state[6] ));
 sky130_fd_sc_hd__dfxtp_2 _40277_ (.CLK(clk),
    .D(_02771_),
    .Q(\cpuregs[8][0] ));
 sky130_fd_sc_hd__dfxtp_2 _40278_ (.CLK(clk),
    .D(_02772_),
    .Q(\cpuregs[8][1] ));
 sky130_fd_sc_hd__dfxtp_2 _40279_ (.CLK(clk),
    .D(_02773_),
    .Q(\cpuregs[8][2] ));
 sky130_fd_sc_hd__dfxtp_2 _40280_ (.CLK(clk),
    .D(_02774_),
    .Q(\cpuregs[8][3] ));
 sky130_fd_sc_hd__dfxtp_2 _40281_ (.CLK(clk),
    .D(_02775_),
    .Q(\cpuregs[8][4] ));
 sky130_fd_sc_hd__dfxtp_2 _40282_ (.CLK(clk),
    .D(_02776_),
    .Q(\cpuregs[8][5] ));
 sky130_fd_sc_hd__dfxtp_2 _40283_ (.CLK(clk),
    .D(_02777_),
    .Q(\cpuregs[8][6] ));
 sky130_fd_sc_hd__dfxtp_2 _40284_ (.CLK(clk),
    .D(_02778_),
    .Q(\cpuregs[8][7] ));
 sky130_fd_sc_hd__dfxtp_2 _40285_ (.CLK(clk),
    .D(_02779_),
    .Q(\cpuregs[8][8] ));
 sky130_fd_sc_hd__dfxtp_2 _40286_ (.CLK(clk),
    .D(_02780_),
    .Q(\cpuregs[8][9] ));
 sky130_fd_sc_hd__dfxtp_2 _40287_ (.CLK(clk),
    .D(_02781_),
    .Q(\cpuregs[8][10] ));
 sky130_fd_sc_hd__dfxtp_2 _40288_ (.CLK(clk),
    .D(_02782_),
    .Q(\cpuregs[8][11] ));
 sky130_fd_sc_hd__dfxtp_2 _40289_ (.CLK(clk),
    .D(_02783_),
    .Q(\cpuregs[8][12] ));
 sky130_fd_sc_hd__dfxtp_2 _40290_ (.CLK(clk),
    .D(_02784_),
    .Q(\cpuregs[8][13] ));
 sky130_fd_sc_hd__dfxtp_2 _40291_ (.CLK(clk),
    .D(_02785_),
    .Q(\cpuregs[8][14] ));
 sky130_fd_sc_hd__dfxtp_2 _40292_ (.CLK(clk),
    .D(_02786_),
    .Q(\cpuregs[8][15] ));
 sky130_fd_sc_hd__dfxtp_2 _40293_ (.CLK(clk),
    .D(_02787_),
    .Q(\cpuregs[8][16] ));
 sky130_fd_sc_hd__dfxtp_2 _40294_ (.CLK(clk),
    .D(_02788_),
    .Q(\cpuregs[8][17] ));
 sky130_fd_sc_hd__dfxtp_2 _40295_ (.CLK(clk),
    .D(_02789_),
    .Q(\cpuregs[8][18] ));
 sky130_fd_sc_hd__dfxtp_2 _40296_ (.CLK(clk),
    .D(_02790_),
    .Q(\cpuregs[8][19] ));
 sky130_fd_sc_hd__dfxtp_2 _40297_ (.CLK(clk),
    .D(_02791_),
    .Q(\cpuregs[8][20] ));
 sky130_fd_sc_hd__dfxtp_2 _40298_ (.CLK(clk),
    .D(_02792_),
    .Q(\cpuregs[8][21] ));
 sky130_fd_sc_hd__dfxtp_2 _40299_ (.CLK(clk),
    .D(_02793_),
    .Q(\cpuregs[8][22] ));
 sky130_fd_sc_hd__dfxtp_2 _40300_ (.CLK(clk),
    .D(_02794_),
    .Q(\cpuregs[8][23] ));
 sky130_fd_sc_hd__dfxtp_2 _40301_ (.CLK(clk),
    .D(_02795_),
    .Q(\cpuregs[8][24] ));
 sky130_fd_sc_hd__dfxtp_2 _40302_ (.CLK(clk),
    .D(_02796_),
    .Q(\cpuregs[8][25] ));
 sky130_fd_sc_hd__dfxtp_2 _40303_ (.CLK(clk),
    .D(_02797_),
    .Q(\cpuregs[8][26] ));
 sky130_fd_sc_hd__dfxtp_2 _40304_ (.CLK(clk),
    .D(_02798_),
    .Q(\cpuregs[8][27] ));
 sky130_fd_sc_hd__dfxtp_2 _40305_ (.CLK(clk),
    .D(_02799_),
    .Q(\cpuregs[8][28] ));
 sky130_fd_sc_hd__dfxtp_2 _40306_ (.CLK(clk),
    .D(_02800_),
    .Q(\cpuregs[8][29] ));
 sky130_fd_sc_hd__dfxtp_2 _40307_ (.CLK(clk),
    .D(_02801_),
    .Q(\cpuregs[8][30] ));
 sky130_fd_sc_hd__dfxtp_2 _40308_ (.CLK(clk),
    .D(_02802_),
    .Q(\cpuregs[8][31] ));
 sky130_fd_sc_hd__dfxtp_2 _40309_ (.CLK(clk),
    .D(_02803_),
    .Q(\cpuregs[14][0] ));
 sky130_fd_sc_hd__dfxtp_2 _40310_ (.CLK(clk),
    .D(_02804_),
    .Q(\cpuregs[14][1] ));
 sky130_fd_sc_hd__dfxtp_2 _40311_ (.CLK(clk),
    .D(_02805_),
    .Q(\cpuregs[14][2] ));
 sky130_fd_sc_hd__dfxtp_2 _40312_ (.CLK(clk),
    .D(_02806_),
    .Q(\cpuregs[14][3] ));
 sky130_fd_sc_hd__dfxtp_2 _40313_ (.CLK(clk),
    .D(_02807_),
    .Q(\cpuregs[14][4] ));
 sky130_fd_sc_hd__dfxtp_2 _40314_ (.CLK(clk),
    .D(_02808_),
    .Q(\cpuregs[14][5] ));
 sky130_fd_sc_hd__dfxtp_2 _40315_ (.CLK(clk),
    .D(_02809_),
    .Q(\cpuregs[14][6] ));
 sky130_fd_sc_hd__dfxtp_2 _40316_ (.CLK(clk),
    .D(_02810_),
    .Q(\cpuregs[14][7] ));
 sky130_fd_sc_hd__dfxtp_2 _40317_ (.CLK(clk),
    .D(_02811_),
    .Q(\cpuregs[14][8] ));
 sky130_fd_sc_hd__dfxtp_2 _40318_ (.CLK(clk),
    .D(_02812_),
    .Q(\cpuregs[14][9] ));
 sky130_fd_sc_hd__dfxtp_2 _40319_ (.CLK(clk),
    .D(_02813_),
    .Q(\cpuregs[14][10] ));
 sky130_fd_sc_hd__dfxtp_2 _40320_ (.CLK(clk),
    .D(_02814_),
    .Q(\cpuregs[14][11] ));
 sky130_fd_sc_hd__dfxtp_2 _40321_ (.CLK(clk),
    .D(_02815_),
    .Q(\cpuregs[14][12] ));
 sky130_fd_sc_hd__dfxtp_2 _40322_ (.CLK(clk),
    .D(_02816_),
    .Q(\cpuregs[14][13] ));
 sky130_fd_sc_hd__dfxtp_2 _40323_ (.CLK(clk),
    .D(_02817_),
    .Q(\cpuregs[14][14] ));
 sky130_fd_sc_hd__dfxtp_2 _40324_ (.CLK(clk),
    .D(_02818_),
    .Q(\cpuregs[14][15] ));
 sky130_fd_sc_hd__dfxtp_2 _40325_ (.CLK(clk),
    .D(_02819_),
    .Q(\cpuregs[14][16] ));
 sky130_fd_sc_hd__dfxtp_2 _40326_ (.CLK(clk),
    .D(_02820_),
    .Q(\cpuregs[14][17] ));
 sky130_fd_sc_hd__dfxtp_2 _40327_ (.CLK(clk),
    .D(_02821_),
    .Q(\cpuregs[14][18] ));
 sky130_fd_sc_hd__dfxtp_2 _40328_ (.CLK(clk),
    .D(_02822_),
    .Q(\cpuregs[14][19] ));
 sky130_fd_sc_hd__dfxtp_2 _40329_ (.CLK(clk),
    .D(_02823_),
    .Q(\cpuregs[14][20] ));
 sky130_fd_sc_hd__dfxtp_2 _40330_ (.CLK(clk),
    .D(_02824_),
    .Q(\cpuregs[14][21] ));
 sky130_fd_sc_hd__dfxtp_2 _40331_ (.CLK(clk),
    .D(_02825_),
    .Q(\cpuregs[14][22] ));
 sky130_fd_sc_hd__dfxtp_2 _40332_ (.CLK(clk),
    .D(_02826_),
    .Q(\cpuregs[14][23] ));
 sky130_fd_sc_hd__dfxtp_2 _40333_ (.CLK(clk),
    .D(_02827_),
    .Q(\cpuregs[14][24] ));
 sky130_fd_sc_hd__dfxtp_2 _40334_ (.CLK(clk),
    .D(_02828_),
    .Q(\cpuregs[14][25] ));
 sky130_fd_sc_hd__dfxtp_2 _40335_ (.CLK(clk),
    .D(_02829_),
    .Q(\cpuregs[14][26] ));
 sky130_fd_sc_hd__dfxtp_2 _40336_ (.CLK(clk),
    .D(_02830_),
    .Q(\cpuregs[14][27] ));
 sky130_fd_sc_hd__dfxtp_2 _40337_ (.CLK(clk),
    .D(_02831_),
    .Q(\cpuregs[14][28] ));
 sky130_fd_sc_hd__dfxtp_2 _40338_ (.CLK(clk),
    .D(_02832_),
    .Q(\cpuregs[14][29] ));
 sky130_fd_sc_hd__dfxtp_2 _40339_ (.CLK(clk),
    .D(_02833_),
    .Q(\cpuregs[14][30] ));
 sky130_fd_sc_hd__dfxtp_2 _40340_ (.CLK(clk),
    .D(_02834_),
    .Q(\cpuregs[14][31] ));
 sky130_fd_sc_hd__dfxtp_2 _40341_ (.CLK(clk),
    .D(_02835_),
    .Q(\cpuregs[0][0] ));
 sky130_fd_sc_hd__dfxtp_2 _40342_ (.CLK(clk),
    .D(_02836_),
    .Q(\cpuregs[0][1] ));
 sky130_fd_sc_hd__dfxtp_2 _40343_ (.CLK(clk),
    .D(_02837_),
    .Q(\cpuregs[0][2] ));
 sky130_fd_sc_hd__dfxtp_2 _40344_ (.CLK(clk),
    .D(_02838_),
    .Q(\cpuregs[0][3] ));
 sky130_fd_sc_hd__dfxtp_2 _40345_ (.CLK(clk),
    .D(_02839_),
    .Q(\cpuregs[0][4] ));
 sky130_fd_sc_hd__dfxtp_2 _40346_ (.CLK(clk),
    .D(_02840_),
    .Q(\cpuregs[0][5] ));
 sky130_fd_sc_hd__dfxtp_2 _40347_ (.CLK(clk),
    .D(_02841_),
    .Q(\cpuregs[0][6] ));
 sky130_fd_sc_hd__dfxtp_2 _40348_ (.CLK(clk),
    .D(_02842_),
    .Q(\cpuregs[0][7] ));
 sky130_fd_sc_hd__dfxtp_2 _40349_ (.CLK(clk),
    .D(_02843_),
    .Q(\cpuregs[0][8] ));
 sky130_fd_sc_hd__dfxtp_2 _40350_ (.CLK(clk),
    .D(_02844_),
    .Q(\cpuregs[0][9] ));
 sky130_fd_sc_hd__dfxtp_2 _40351_ (.CLK(clk),
    .D(_02845_),
    .Q(\cpuregs[0][10] ));
 sky130_fd_sc_hd__dfxtp_2 _40352_ (.CLK(clk),
    .D(_02846_),
    .Q(\cpuregs[0][11] ));
 sky130_fd_sc_hd__dfxtp_2 _40353_ (.CLK(clk),
    .D(_02847_),
    .Q(\cpuregs[0][12] ));
 sky130_fd_sc_hd__dfxtp_2 _40354_ (.CLK(clk),
    .D(_02848_),
    .Q(\cpuregs[0][13] ));
 sky130_fd_sc_hd__dfxtp_2 _40355_ (.CLK(clk),
    .D(_02849_),
    .Q(\cpuregs[0][14] ));
 sky130_fd_sc_hd__dfxtp_2 _40356_ (.CLK(clk),
    .D(_02850_),
    .Q(\cpuregs[0][15] ));
 sky130_fd_sc_hd__dfxtp_2 _40357_ (.CLK(clk),
    .D(_02851_),
    .Q(\cpuregs[0][16] ));
 sky130_fd_sc_hd__dfxtp_2 _40358_ (.CLK(clk),
    .D(_02852_),
    .Q(\cpuregs[0][17] ));
 sky130_fd_sc_hd__dfxtp_2 _40359_ (.CLK(clk),
    .D(_02853_),
    .Q(\cpuregs[0][18] ));
 sky130_fd_sc_hd__dfxtp_2 _40360_ (.CLK(clk),
    .D(_02854_),
    .Q(\cpuregs[0][19] ));
 sky130_fd_sc_hd__dfxtp_2 _40361_ (.CLK(clk),
    .D(_02855_),
    .Q(\cpuregs[0][20] ));
 sky130_fd_sc_hd__dfxtp_2 _40362_ (.CLK(clk),
    .D(_02856_),
    .Q(\cpuregs[0][21] ));
 sky130_fd_sc_hd__dfxtp_2 _40363_ (.CLK(clk),
    .D(_02857_),
    .Q(\cpuregs[0][22] ));
 sky130_fd_sc_hd__dfxtp_2 _40364_ (.CLK(clk),
    .D(_02858_),
    .Q(\cpuregs[0][23] ));
 sky130_fd_sc_hd__dfxtp_2 _40365_ (.CLK(clk),
    .D(_02859_),
    .Q(\cpuregs[0][24] ));
 sky130_fd_sc_hd__dfxtp_2 _40366_ (.CLK(clk),
    .D(_02860_),
    .Q(\cpuregs[0][25] ));
 sky130_fd_sc_hd__dfxtp_2 _40367_ (.CLK(clk),
    .D(_02861_),
    .Q(\cpuregs[0][26] ));
 sky130_fd_sc_hd__dfxtp_2 _40368_ (.CLK(clk),
    .D(_02862_),
    .Q(\cpuregs[0][27] ));
 sky130_fd_sc_hd__dfxtp_2 _40369_ (.CLK(clk),
    .D(_02863_),
    .Q(\cpuregs[0][28] ));
 sky130_fd_sc_hd__dfxtp_2 _40370_ (.CLK(clk),
    .D(_02864_),
    .Q(\cpuregs[0][29] ));
 sky130_fd_sc_hd__dfxtp_2 _40371_ (.CLK(clk),
    .D(_02865_),
    .Q(\cpuregs[0][30] ));
 sky130_fd_sc_hd__dfxtp_2 _40372_ (.CLK(clk),
    .D(_02866_),
    .Q(\cpuregs[0][31] ));
 sky130_fd_sc_hd__dfxtp_2 _40373_ (.CLK(clk),
    .D(_02867_),
    .Q(\cpuregs[10][0] ));
 sky130_fd_sc_hd__dfxtp_2 _40374_ (.CLK(clk),
    .D(_02868_),
    .Q(\cpuregs[10][1] ));
 sky130_fd_sc_hd__dfxtp_2 _40375_ (.CLK(clk),
    .D(_02869_),
    .Q(\cpuregs[10][2] ));
 sky130_fd_sc_hd__dfxtp_2 _40376_ (.CLK(clk),
    .D(_02870_),
    .Q(\cpuregs[10][3] ));
 sky130_fd_sc_hd__dfxtp_2 _40377_ (.CLK(clk),
    .D(_02871_),
    .Q(\cpuregs[10][4] ));
 sky130_fd_sc_hd__dfxtp_2 _40378_ (.CLK(clk),
    .D(_02872_),
    .Q(\cpuregs[10][5] ));
 sky130_fd_sc_hd__dfxtp_2 _40379_ (.CLK(clk),
    .D(_02873_),
    .Q(\cpuregs[10][6] ));
 sky130_fd_sc_hd__dfxtp_2 _40380_ (.CLK(clk),
    .D(_02874_),
    .Q(\cpuregs[10][7] ));
 sky130_fd_sc_hd__dfxtp_2 _40381_ (.CLK(clk),
    .D(_02875_),
    .Q(\cpuregs[10][8] ));
 sky130_fd_sc_hd__dfxtp_2 _40382_ (.CLK(clk),
    .D(_02876_),
    .Q(\cpuregs[10][9] ));
 sky130_fd_sc_hd__dfxtp_2 _40383_ (.CLK(clk),
    .D(_02877_),
    .Q(\cpuregs[10][10] ));
 sky130_fd_sc_hd__dfxtp_2 _40384_ (.CLK(clk),
    .D(_02878_),
    .Q(\cpuregs[10][11] ));
 sky130_fd_sc_hd__dfxtp_2 _40385_ (.CLK(clk),
    .D(_02879_),
    .Q(\cpuregs[10][12] ));
 sky130_fd_sc_hd__dfxtp_2 _40386_ (.CLK(clk),
    .D(_02880_),
    .Q(\cpuregs[10][13] ));
 sky130_fd_sc_hd__dfxtp_2 _40387_ (.CLK(clk),
    .D(_02881_),
    .Q(\cpuregs[10][14] ));
 sky130_fd_sc_hd__dfxtp_2 _40388_ (.CLK(clk),
    .D(_02882_),
    .Q(\cpuregs[10][15] ));
 sky130_fd_sc_hd__dfxtp_2 _40389_ (.CLK(clk),
    .D(_02883_),
    .Q(\cpuregs[10][16] ));
 sky130_fd_sc_hd__dfxtp_2 _40390_ (.CLK(clk),
    .D(_02884_),
    .Q(\cpuregs[10][17] ));
 sky130_fd_sc_hd__dfxtp_2 _40391_ (.CLK(clk),
    .D(_02885_),
    .Q(\cpuregs[10][18] ));
 sky130_fd_sc_hd__dfxtp_2 _40392_ (.CLK(clk),
    .D(_02886_),
    .Q(\cpuregs[10][19] ));
 sky130_fd_sc_hd__dfxtp_2 _40393_ (.CLK(clk),
    .D(_02887_),
    .Q(\cpuregs[10][20] ));
 sky130_fd_sc_hd__dfxtp_2 _40394_ (.CLK(clk),
    .D(_02888_),
    .Q(\cpuregs[10][21] ));
 sky130_fd_sc_hd__dfxtp_2 _40395_ (.CLK(clk),
    .D(_02889_),
    .Q(\cpuregs[10][22] ));
 sky130_fd_sc_hd__dfxtp_2 _40396_ (.CLK(clk),
    .D(_02890_),
    .Q(\cpuregs[10][23] ));
 sky130_fd_sc_hd__dfxtp_2 _40397_ (.CLK(clk),
    .D(_02891_),
    .Q(\cpuregs[10][24] ));
 sky130_fd_sc_hd__dfxtp_2 _40398_ (.CLK(clk),
    .D(_02892_),
    .Q(\cpuregs[10][25] ));
 sky130_fd_sc_hd__dfxtp_2 _40399_ (.CLK(clk),
    .D(_02893_),
    .Q(\cpuregs[10][26] ));
 sky130_fd_sc_hd__dfxtp_2 _40400_ (.CLK(clk),
    .D(_02894_),
    .Q(\cpuregs[10][27] ));
 sky130_fd_sc_hd__dfxtp_2 _40401_ (.CLK(clk),
    .D(_02895_),
    .Q(\cpuregs[10][28] ));
 sky130_fd_sc_hd__dfxtp_2 _40402_ (.CLK(clk),
    .D(_02896_),
    .Q(\cpuregs[10][29] ));
 sky130_fd_sc_hd__dfxtp_2 _40403_ (.CLK(clk),
    .D(_02897_),
    .Q(\cpuregs[10][30] ));
 sky130_fd_sc_hd__dfxtp_2 _40404_ (.CLK(clk),
    .D(_02898_),
    .Q(\cpuregs[10][31] ));
 sky130_fd_sc_hd__dfxtp_2 _40405_ (.CLK(clk),
    .D(_02899_),
    .Q(\cpuregs[18][0] ));
 sky130_fd_sc_hd__dfxtp_2 _40406_ (.CLK(clk),
    .D(_02900_),
    .Q(\cpuregs[18][1] ));
 sky130_fd_sc_hd__dfxtp_2 _40407_ (.CLK(clk),
    .D(_02901_),
    .Q(\cpuregs[18][2] ));
 sky130_fd_sc_hd__dfxtp_2 _40408_ (.CLK(clk),
    .D(_02902_),
    .Q(\cpuregs[18][3] ));
 sky130_fd_sc_hd__dfxtp_2 _40409_ (.CLK(clk),
    .D(_02903_),
    .Q(\cpuregs[18][4] ));
 sky130_fd_sc_hd__dfxtp_2 _40410_ (.CLK(clk),
    .D(_02904_),
    .Q(\cpuregs[18][5] ));
 sky130_fd_sc_hd__dfxtp_2 _40411_ (.CLK(clk),
    .D(_02905_),
    .Q(\cpuregs[18][6] ));
 sky130_fd_sc_hd__dfxtp_2 _40412_ (.CLK(clk),
    .D(_02906_),
    .Q(\cpuregs[18][7] ));
 sky130_fd_sc_hd__dfxtp_2 _40413_ (.CLK(clk),
    .D(_02907_),
    .Q(\cpuregs[18][8] ));
 sky130_fd_sc_hd__dfxtp_2 _40414_ (.CLK(clk),
    .D(_02908_),
    .Q(\cpuregs[18][9] ));
 sky130_fd_sc_hd__dfxtp_2 _40415_ (.CLK(clk),
    .D(_02909_),
    .Q(\cpuregs[18][10] ));
 sky130_fd_sc_hd__dfxtp_2 _40416_ (.CLK(clk),
    .D(_02910_),
    .Q(\cpuregs[18][11] ));
 sky130_fd_sc_hd__dfxtp_2 _40417_ (.CLK(clk),
    .D(_02911_),
    .Q(\cpuregs[18][12] ));
 sky130_fd_sc_hd__dfxtp_2 _40418_ (.CLK(clk),
    .D(_02912_),
    .Q(\cpuregs[18][13] ));
 sky130_fd_sc_hd__dfxtp_2 _40419_ (.CLK(clk),
    .D(_02913_),
    .Q(\cpuregs[18][14] ));
 sky130_fd_sc_hd__dfxtp_2 _40420_ (.CLK(clk),
    .D(_02914_),
    .Q(\cpuregs[18][15] ));
 sky130_fd_sc_hd__dfxtp_2 _40421_ (.CLK(clk),
    .D(_02915_),
    .Q(\cpuregs[18][16] ));
 sky130_fd_sc_hd__dfxtp_2 _40422_ (.CLK(clk),
    .D(_02916_),
    .Q(\cpuregs[18][17] ));
 sky130_fd_sc_hd__dfxtp_2 _40423_ (.CLK(clk),
    .D(_02917_),
    .Q(\cpuregs[18][18] ));
 sky130_fd_sc_hd__dfxtp_2 _40424_ (.CLK(clk),
    .D(_02918_),
    .Q(\cpuregs[18][19] ));
 sky130_fd_sc_hd__dfxtp_2 _40425_ (.CLK(clk),
    .D(_02919_),
    .Q(\cpuregs[18][20] ));
 sky130_fd_sc_hd__dfxtp_2 _40426_ (.CLK(clk),
    .D(_02920_),
    .Q(\cpuregs[18][21] ));
 sky130_fd_sc_hd__dfxtp_2 _40427_ (.CLK(clk),
    .D(_02921_),
    .Q(\cpuregs[18][22] ));
 sky130_fd_sc_hd__dfxtp_2 _40428_ (.CLK(clk),
    .D(_02922_),
    .Q(\cpuregs[18][23] ));
 sky130_fd_sc_hd__dfxtp_2 _40429_ (.CLK(clk),
    .D(_02923_),
    .Q(\cpuregs[18][24] ));
 sky130_fd_sc_hd__dfxtp_2 _40430_ (.CLK(clk),
    .D(_02924_),
    .Q(\cpuregs[18][25] ));
 sky130_fd_sc_hd__dfxtp_2 _40431_ (.CLK(clk),
    .D(_02925_),
    .Q(\cpuregs[18][26] ));
 sky130_fd_sc_hd__dfxtp_2 _40432_ (.CLK(clk),
    .D(_02926_),
    .Q(\cpuregs[18][27] ));
 sky130_fd_sc_hd__dfxtp_2 _40433_ (.CLK(clk),
    .D(_02927_),
    .Q(\cpuregs[18][28] ));
 sky130_fd_sc_hd__dfxtp_2 _40434_ (.CLK(clk),
    .D(_02928_),
    .Q(\cpuregs[18][29] ));
 sky130_fd_sc_hd__dfxtp_2 _40435_ (.CLK(clk),
    .D(_02929_),
    .Q(\cpuregs[18][30] ));
 sky130_fd_sc_hd__dfxtp_2 _40436_ (.CLK(clk),
    .D(_02930_),
    .Q(\cpuregs[18][31] ));
 sky130_fd_sc_hd__dfxtp_2 _40437_ (.CLK(clk),
    .D(_02931_),
    .Q(\mem_rdata_q[0] ));
 sky130_fd_sc_hd__dfxtp_2 _40438_ (.CLK(clk),
    .D(_02932_),
    .Q(\mem_rdata_q[1] ));
 sky130_fd_sc_hd__dfxtp_2 _40439_ (.CLK(clk),
    .D(_02933_),
    .Q(\mem_rdata_q[2] ));
 sky130_fd_sc_hd__dfxtp_2 _40440_ (.CLK(clk),
    .D(_02934_),
    .Q(\mem_rdata_q[3] ));
 sky130_fd_sc_hd__dfxtp_2 _40441_ (.CLK(clk),
    .D(_02935_),
    .Q(\mem_rdata_q[4] ));
 sky130_fd_sc_hd__dfxtp_2 _40442_ (.CLK(clk),
    .D(_02936_),
    .Q(\mem_rdata_q[5] ));
 sky130_fd_sc_hd__dfxtp_2 _40443_ (.CLK(clk),
    .D(_02937_),
    .Q(\mem_rdata_q[6] ));
 sky130_fd_sc_hd__dfxtp_2 _40444_ (.CLK(clk),
    .D(_02938_),
    .Q(\mem_rdata_q[7] ));
 sky130_fd_sc_hd__dfxtp_2 _40445_ (.CLK(clk),
    .D(_02939_),
    .Q(\mem_rdata_q[8] ));
 sky130_fd_sc_hd__dfxtp_2 _40446_ (.CLK(clk),
    .D(_02940_),
    .Q(\mem_rdata_q[9] ));
 sky130_fd_sc_hd__dfxtp_2 _40447_ (.CLK(clk),
    .D(_02941_),
    .Q(\mem_rdata_q[10] ));
 sky130_fd_sc_hd__dfxtp_2 _40448_ (.CLK(clk),
    .D(_02942_),
    .Q(\mem_rdata_q[11] ));
 sky130_fd_sc_hd__dfxtp_2 _40449_ (.CLK(clk),
    .D(_02943_),
    .Q(\mem_rdata_q[12] ));
 sky130_fd_sc_hd__dfxtp_2 _40450_ (.CLK(clk),
    .D(_02944_),
    .Q(\mem_rdata_q[13] ));
 sky130_fd_sc_hd__dfxtp_2 _40451_ (.CLK(clk),
    .D(_02945_),
    .Q(\mem_rdata_q[14] ));
 sky130_fd_sc_hd__dfxtp_2 _40452_ (.CLK(clk),
    .D(_02946_),
    .Q(\mem_rdata_q[15] ));
 sky130_fd_sc_hd__dfxtp_2 _40453_ (.CLK(clk),
    .D(_02947_),
    .Q(\mem_rdata_q[16] ));
 sky130_fd_sc_hd__dfxtp_2 _40454_ (.CLK(clk),
    .D(_02948_),
    .Q(\mem_rdata_q[17] ));
 sky130_fd_sc_hd__dfxtp_2 _40455_ (.CLK(clk),
    .D(_02949_),
    .Q(\mem_rdata_q[18] ));
 sky130_fd_sc_hd__dfxtp_2 _40456_ (.CLK(clk),
    .D(_02950_),
    .Q(\mem_rdata_q[19] ));
 sky130_fd_sc_hd__dfxtp_2 _40457_ (.CLK(clk),
    .D(_02951_),
    .Q(\mem_rdata_q[20] ));
 sky130_fd_sc_hd__dfxtp_2 _40458_ (.CLK(clk),
    .D(_02952_),
    .Q(\mem_rdata_q[21] ));
 sky130_fd_sc_hd__dfxtp_2 _40459_ (.CLK(clk),
    .D(_02953_),
    .Q(\mem_rdata_q[22] ));
 sky130_fd_sc_hd__dfxtp_2 _40460_ (.CLK(clk),
    .D(_02954_),
    .Q(\mem_rdata_q[23] ));
 sky130_fd_sc_hd__dfxtp_2 _40461_ (.CLK(clk),
    .D(_02955_),
    .Q(\mem_rdata_q[24] ));
 sky130_fd_sc_hd__dfxtp_2 _40462_ (.CLK(clk),
    .D(_02956_),
    .Q(\mem_rdata_q[25] ));
 sky130_fd_sc_hd__dfxtp_2 _40463_ (.CLK(clk),
    .D(_02957_),
    .Q(\mem_rdata_q[26] ));
 sky130_fd_sc_hd__dfxtp_2 _40464_ (.CLK(clk),
    .D(_02958_),
    .Q(\mem_rdata_q[27] ));
 sky130_fd_sc_hd__dfxtp_2 _40465_ (.CLK(clk),
    .D(_02959_),
    .Q(\mem_rdata_q[28] ));
 sky130_fd_sc_hd__dfxtp_2 _40466_ (.CLK(clk),
    .D(_02960_),
    .Q(\mem_rdata_q[29] ));
 sky130_fd_sc_hd__dfxtp_2 _40467_ (.CLK(clk),
    .D(_02961_),
    .Q(\mem_rdata_q[30] ));
 sky130_fd_sc_hd__dfxtp_2 _40468_ (.CLK(clk),
    .D(_02962_),
    .Q(\mem_rdata_q[31] ));
 sky130_fd_sc_hd__dfxtp_2 _40469_ (.CLK(clk),
    .D(_02963_),
    .Q(\cpuregs[2][0] ));
 sky130_fd_sc_hd__dfxtp_2 _40470_ (.CLK(clk),
    .D(_02964_),
    .Q(\cpuregs[2][1] ));
 sky130_fd_sc_hd__dfxtp_2 _40471_ (.CLK(clk),
    .D(_02965_),
    .Q(\cpuregs[2][2] ));
 sky130_fd_sc_hd__dfxtp_2 _40472_ (.CLK(clk),
    .D(_02966_),
    .Q(\cpuregs[2][3] ));
 sky130_fd_sc_hd__dfxtp_2 _40473_ (.CLK(clk),
    .D(_02967_),
    .Q(\cpuregs[2][4] ));
 sky130_fd_sc_hd__dfxtp_2 _40474_ (.CLK(clk),
    .D(_02968_),
    .Q(\cpuregs[2][5] ));
 sky130_fd_sc_hd__dfxtp_2 _40475_ (.CLK(clk),
    .D(_02969_),
    .Q(\cpuregs[2][6] ));
 sky130_fd_sc_hd__dfxtp_2 _40476_ (.CLK(clk),
    .D(_02970_),
    .Q(\cpuregs[2][7] ));
 sky130_fd_sc_hd__dfxtp_2 _40477_ (.CLK(clk),
    .D(_02971_),
    .Q(\cpuregs[2][8] ));
 sky130_fd_sc_hd__dfxtp_2 _40478_ (.CLK(clk),
    .D(_02972_),
    .Q(\cpuregs[2][9] ));
 sky130_fd_sc_hd__dfxtp_2 _40479_ (.CLK(clk),
    .D(_02973_),
    .Q(\cpuregs[2][10] ));
 sky130_fd_sc_hd__dfxtp_2 _40480_ (.CLK(clk),
    .D(_02974_),
    .Q(\cpuregs[2][11] ));
 sky130_fd_sc_hd__dfxtp_2 _40481_ (.CLK(clk),
    .D(_02975_),
    .Q(\cpuregs[2][12] ));
 sky130_fd_sc_hd__dfxtp_2 _40482_ (.CLK(clk),
    .D(_02976_),
    .Q(\cpuregs[2][13] ));
 sky130_fd_sc_hd__dfxtp_2 _40483_ (.CLK(clk),
    .D(_02977_),
    .Q(\cpuregs[2][14] ));
 sky130_fd_sc_hd__dfxtp_2 _40484_ (.CLK(clk),
    .D(_02978_),
    .Q(\cpuregs[2][15] ));
 sky130_fd_sc_hd__dfxtp_2 _40485_ (.CLK(clk),
    .D(_02979_),
    .Q(\cpuregs[2][16] ));
 sky130_fd_sc_hd__dfxtp_2 _40486_ (.CLK(clk),
    .D(_02980_),
    .Q(\cpuregs[2][17] ));
 sky130_fd_sc_hd__dfxtp_2 _40487_ (.CLK(clk),
    .D(_02981_),
    .Q(\cpuregs[2][18] ));
 sky130_fd_sc_hd__dfxtp_2 _40488_ (.CLK(clk),
    .D(_02982_),
    .Q(\cpuregs[2][19] ));
 sky130_fd_sc_hd__dfxtp_2 _40489_ (.CLK(clk),
    .D(_02983_),
    .Q(\cpuregs[2][20] ));
 sky130_fd_sc_hd__dfxtp_2 _40490_ (.CLK(clk),
    .D(_02984_),
    .Q(\cpuregs[2][21] ));
 sky130_fd_sc_hd__dfxtp_2 _40491_ (.CLK(clk),
    .D(_02985_),
    .Q(\cpuregs[2][22] ));
 sky130_fd_sc_hd__dfxtp_2 _40492_ (.CLK(clk),
    .D(_02986_),
    .Q(\cpuregs[2][23] ));
 sky130_fd_sc_hd__dfxtp_2 _40493_ (.CLK(clk),
    .D(_02987_),
    .Q(\cpuregs[2][24] ));
 sky130_fd_sc_hd__dfxtp_2 _40494_ (.CLK(clk),
    .D(_02988_),
    .Q(\cpuregs[2][25] ));
 sky130_fd_sc_hd__dfxtp_2 _40495_ (.CLK(clk),
    .D(_02989_),
    .Q(\cpuregs[2][26] ));
 sky130_fd_sc_hd__dfxtp_2 _40496_ (.CLK(clk),
    .D(_02990_),
    .Q(\cpuregs[2][27] ));
 sky130_fd_sc_hd__dfxtp_2 _40497_ (.CLK(clk),
    .D(_02991_),
    .Q(\cpuregs[2][28] ));
 sky130_fd_sc_hd__dfxtp_2 _40498_ (.CLK(clk),
    .D(_02992_),
    .Q(\cpuregs[2][29] ));
 sky130_fd_sc_hd__dfxtp_2 _40499_ (.CLK(clk),
    .D(_02993_),
    .Q(\cpuregs[2][30] ));
 sky130_fd_sc_hd__dfxtp_2 _40500_ (.CLK(clk),
    .D(_02994_),
    .Q(\cpuregs[2][31] ));
 sky130_fd_sc_hd__dfxtp_2 _40501_ (.CLK(clk),
    .D(_02995_),
    .Q(\cpuregs[5][0] ));
 sky130_fd_sc_hd__dfxtp_2 _40502_ (.CLK(clk),
    .D(_02996_),
    .Q(\cpuregs[5][1] ));
 sky130_fd_sc_hd__dfxtp_2 _40503_ (.CLK(clk),
    .D(_02997_),
    .Q(\cpuregs[5][2] ));
 sky130_fd_sc_hd__dfxtp_2 _40504_ (.CLK(clk),
    .D(_02998_),
    .Q(\cpuregs[5][3] ));
 sky130_fd_sc_hd__dfxtp_2 _40505_ (.CLK(clk),
    .D(_02999_),
    .Q(\cpuregs[5][4] ));
 sky130_fd_sc_hd__dfxtp_2 _40506_ (.CLK(clk),
    .D(_03000_),
    .Q(\cpuregs[5][5] ));
 sky130_fd_sc_hd__dfxtp_2 _40507_ (.CLK(clk),
    .D(_03001_),
    .Q(\cpuregs[5][6] ));
 sky130_fd_sc_hd__dfxtp_2 _40508_ (.CLK(clk),
    .D(_03002_),
    .Q(\cpuregs[5][7] ));
 sky130_fd_sc_hd__dfxtp_2 _40509_ (.CLK(clk),
    .D(_03003_),
    .Q(\cpuregs[5][8] ));
 sky130_fd_sc_hd__dfxtp_2 _40510_ (.CLK(clk),
    .D(_03004_),
    .Q(\cpuregs[5][9] ));
 sky130_fd_sc_hd__dfxtp_2 _40511_ (.CLK(clk),
    .D(_03005_),
    .Q(\cpuregs[5][10] ));
 sky130_fd_sc_hd__dfxtp_2 _40512_ (.CLK(clk),
    .D(_03006_),
    .Q(\cpuregs[5][11] ));
 sky130_fd_sc_hd__dfxtp_2 _40513_ (.CLK(clk),
    .D(_03007_),
    .Q(\cpuregs[5][12] ));
 sky130_fd_sc_hd__dfxtp_2 _40514_ (.CLK(clk),
    .D(_03008_),
    .Q(\cpuregs[5][13] ));
 sky130_fd_sc_hd__dfxtp_2 _40515_ (.CLK(clk),
    .D(_03009_),
    .Q(\cpuregs[5][14] ));
 sky130_fd_sc_hd__dfxtp_2 _40516_ (.CLK(clk),
    .D(_03010_),
    .Q(\cpuregs[5][15] ));
 sky130_fd_sc_hd__dfxtp_2 _40517_ (.CLK(clk),
    .D(_03011_),
    .Q(\cpuregs[5][16] ));
 sky130_fd_sc_hd__dfxtp_2 _40518_ (.CLK(clk),
    .D(_03012_),
    .Q(\cpuregs[5][17] ));
 sky130_fd_sc_hd__dfxtp_2 _40519_ (.CLK(clk),
    .D(_03013_),
    .Q(\cpuregs[5][18] ));
 sky130_fd_sc_hd__dfxtp_2 _40520_ (.CLK(clk),
    .D(_03014_),
    .Q(\cpuregs[5][19] ));
 sky130_fd_sc_hd__dfxtp_2 _40521_ (.CLK(clk),
    .D(_03015_),
    .Q(\cpuregs[5][20] ));
 sky130_fd_sc_hd__dfxtp_2 _40522_ (.CLK(clk),
    .D(_03016_),
    .Q(\cpuregs[5][21] ));
 sky130_fd_sc_hd__dfxtp_2 _40523_ (.CLK(clk),
    .D(_03017_),
    .Q(\cpuregs[5][22] ));
 sky130_fd_sc_hd__dfxtp_2 _40524_ (.CLK(clk),
    .D(_03018_),
    .Q(\cpuregs[5][23] ));
 sky130_fd_sc_hd__dfxtp_2 _40525_ (.CLK(clk),
    .D(_03019_),
    .Q(\cpuregs[5][24] ));
 sky130_fd_sc_hd__dfxtp_2 _40526_ (.CLK(clk),
    .D(_03020_),
    .Q(\cpuregs[5][25] ));
 sky130_fd_sc_hd__dfxtp_2 _40527_ (.CLK(clk),
    .D(_03021_),
    .Q(\cpuregs[5][26] ));
 sky130_fd_sc_hd__dfxtp_2 _40528_ (.CLK(clk),
    .D(_03022_),
    .Q(\cpuregs[5][27] ));
 sky130_fd_sc_hd__dfxtp_2 _40529_ (.CLK(clk),
    .D(_03023_),
    .Q(\cpuregs[5][28] ));
 sky130_fd_sc_hd__dfxtp_2 _40530_ (.CLK(clk),
    .D(_03024_),
    .Q(\cpuregs[5][29] ));
 sky130_fd_sc_hd__dfxtp_2 _40531_ (.CLK(clk),
    .D(_03025_),
    .Q(\cpuregs[5][30] ));
 sky130_fd_sc_hd__dfxtp_2 _40532_ (.CLK(clk),
    .D(_03026_),
    .Q(\cpuregs[5][31] ));
 sky130_fd_sc_hd__dfxtp_2 _40533_ (.CLK(clk),
    .D(_03027_),
    .Q(\pcpi_mul.rs1[0] ));
 sky130_fd_sc_hd__dfxtp_2 _40534_ (.CLK(clk),
    .D(_03028_),
    .Q(\pcpi_mul.rs1[1] ));
 sky130_fd_sc_hd__dfxtp_2 _40535_ (.CLK(clk),
    .D(_03029_),
    .Q(\pcpi_mul.rs1[2] ));
 sky130_fd_sc_hd__dfxtp_2 _40536_ (.CLK(clk),
    .D(_03030_),
    .Q(\pcpi_mul.rs1[3] ));
 sky130_fd_sc_hd__dfxtp_2 _40537_ (.CLK(clk),
    .D(_03031_),
    .Q(\pcpi_mul.rs1[4] ));
 sky130_fd_sc_hd__dfxtp_2 _40538_ (.CLK(clk),
    .D(_03032_),
    .Q(\pcpi_mul.rs1[5] ));
 sky130_fd_sc_hd__dfxtp_2 _40539_ (.CLK(clk),
    .D(_03033_),
    .Q(\pcpi_mul.rs1[6] ));
 sky130_fd_sc_hd__dfxtp_2 _40540_ (.CLK(clk),
    .D(_03034_),
    .Q(\pcpi_mul.rs1[7] ));
 sky130_fd_sc_hd__dfxtp_2 _40541_ (.CLK(clk),
    .D(_03035_),
    .Q(\pcpi_mul.rs1[8] ));
 sky130_fd_sc_hd__dfxtp_2 _40542_ (.CLK(clk),
    .D(_03036_),
    .Q(\pcpi_mul.rs1[9] ));
 sky130_fd_sc_hd__dfxtp_2 _40543_ (.CLK(clk),
    .D(_03037_),
    .Q(\pcpi_mul.rs1[10] ));
 sky130_fd_sc_hd__dfxtp_2 _40544_ (.CLK(clk),
    .D(_03038_),
    .Q(\pcpi_mul.rs1[11] ));
 sky130_fd_sc_hd__dfxtp_2 _40545_ (.CLK(clk),
    .D(_03039_),
    .Q(\pcpi_mul.rs1[12] ));
 sky130_fd_sc_hd__dfxtp_2 _40546_ (.CLK(clk),
    .D(_03040_),
    .Q(\pcpi_mul.rs1[13] ));
 sky130_fd_sc_hd__dfxtp_2 _40547_ (.CLK(clk),
    .D(_03041_),
    .Q(\pcpi_mul.rs1[14] ));
 sky130_fd_sc_hd__dfxtp_2 _40548_ (.CLK(clk),
    .D(_03042_),
    .Q(\pcpi_mul.rs1[15] ));
 sky130_fd_sc_hd__dfxtp_2 _40549_ (.CLK(clk),
    .D(_03043_),
    .Q(\pcpi_mul.rs1[16] ));
 sky130_fd_sc_hd__dfxtp_2 _40550_ (.CLK(clk),
    .D(_03044_),
    .Q(\pcpi_mul.rs1[17] ));
 sky130_fd_sc_hd__dfxtp_2 _40551_ (.CLK(clk),
    .D(_03045_),
    .Q(\pcpi_mul.rs1[18] ));
 sky130_fd_sc_hd__dfxtp_2 _40552_ (.CLK(clk),
    .D(_03046_),
    .Q(\pcpi_mul.rs1[19] ));
 sky130_fd_sc_hd__dfxtp_2 _40553_ (.CLK(clk),
    .D(_03047_),
    .Q(\pcpi_mul.rs1[20] ));
 sky130_fd_sc_hd__dfxtp_2 _40554_ (.CLK(clk),
    .D(_03048_),
    .Q(\pcpi_mul.rs1[21] ));
 sky130_fd_sc_hd__dfxtp_2 _40555_ (.CLK(clk),
    .D(_03049_),
    .Q(\pcpi_mul.rs1[22] ));
 sky130_fd_sc_hd__dfxtp_2 _40556_ (.CLK(clk),
    .D(_03050_),
    .Q(\pcpi_mul.rs1[23] ));
 sky130_fd_sc_hd__dfxtp_2 _40557_ (.CLK(clk),
    .D(_03051_),
    .Q(\pcpi_mul.rs1[24] ));
 sky130_fd_sc_hd__dfxtp_2 _40558_ (.CLK(clk),
    .D(_03052_),
    .Q(\pcpi_mul.rs1[25] ));
 sky130_fd_sc_hd__dfxtp_2 _40559_ (.CLK(clk),
    .D(_03053_),
    .Q(\pcpi_mul.rs1[26] ));
 sky130_fd_sc_hd__dfxtp_2 _40560_ (.CLK(clk),
    .D(_03054_),
    .Q(\pcpi_mul.rs1[27] ));
 sky130_fd_sc_hd__dfxtp_2 _40561_ (.CLK(clk),
    .D(_03055_),
    .Q(\pcpi_mul.rs1[28] ));
 sky130_fd_sc_hd__dfxtp_2 _40562_ (.CLK(clk),
    .D(_03056_),
    .Q(\pcpi_mul.rs1[29] ));
 sky130_fd_sc_hd__dfxtp_2 _40563_ (.CLK(clk),
    .D(_03057_),
    .Q(\pcpi_mul.rs1[30] ));
 sky130_fd_sc_hd__dfxtp_2 _40564_ (.CLK(clk),
    .D(_03058_),
    .Q(\pcpi_mul.rs1[31] ));
 sky130_fd_sc_hd__dfxtp_2 _40565_ (.CLK(clk),
    .D(_03059_),
    .Q(mem_addr[2]));
 sky130_fd_sc_hd__dfxtp_2 _40566_ (.CLK(clk),
    .D(_03060_),
    .Q(mem_addr[3]));
 sky130_fd_sc_hd__dfxtp_2 _40567_ (.CLK(clk),
    .D(_03061_),
    .Q(mem_addr[4]));
 sky130_fd_sc_hd__dfxtp_2 _40568_ (.CLK(clk),
    .D(_03062_),
    .Q(mem_addr[5]));
 sky130_fd_sc_hd__dfxtp_2 _40569_ (.CLK(clk),
    .D(_03063_),
    .Q(mem_addr[6]));
 sky130_fd_sc_hd__dfxtp_2 _40570_ (.CLK(clk),
    .D(_03064_),
    .Q(mem_addr[7]));
 sky130_fd_sc_hd__dfxtp_2 _40571_ (.CLK(clk),
    .D(_03065_),
    .Q(mem_addr[8]));
 sky130_fd_sc_hd__dfxtp_2 _40572_ (.CLK(clk),
    .D(_03066_),
    .Q(mem_addr[9]));
 sky130_fd_sc_hd__dfxtp_2 _40573_ (.CLK(clk),
    .D(_03067_),
    .Q(mem_addr[10]));
 sky130_fd_sc_hd__dfxtp_2 _40574_ (.CLK(clk),
    .D(_03068_),
    .Q(mem_addr[11]));
 sky130_fd_sc_hd__dfxtp_2 _40575_ (.CLK(clk),
    .D(_03069_),
    .Q(mem_addr[12]));
 sky130_fd_sc_hd__dfxtp_2 _40576_ (.CLK(clk),
    .D(_03070_),
    .Q(mem_addr[13]));
 sky130_fd_sc_hd__dfxtp_2 _40577_ (.CLK(clk),
    .D(_03071_),
    .Q(mem_addr[14]));
 sky130_fd_sc_hd__dfxtp_2 _40578_ (.CLK(clk),
    .D(_03072_),
    .Q(mem_addr[15]));
 sky130_fd_sc_hd__dfxtp_2 _40579_ (.CLK(clk),
    .D(_03073_),
    .Q(mem_addr[16]));
 sky130_fd_sc_hd__dfxtp_2 _40580_ (.CLK(clk),
    .D(_03074_),
    .Q(mem_addr[17]));
 sky130_fd_sc_hd__dfxtp_2 _40581_ (.CLK(clk),
    .D(_03075_),
    .Q(mem_addr[18]));
 sky130_fd_sc_hd__dfxtp_2 _40582_ (.CLK(clk),
    .D(_03076_),
    .Q(mem_addr[19]));
 sky130_fd_sc_hd__dfxtp_2 _40583_ (.CLK(clk),
    .D(_03077_),
    .Q(mem_addr[20]));
 sky130_fd_sc_hd__dfxtp_2 _40584_ (.CLK(clk),
    .D(_03078_),
    .Q(mem_addr[21]));
 sky130_fd_sc_hd__dfxtp_2 _40585_ (.CLK(clk),
    .D(_03079_),
    .Q(mem_addr[22]));
 sky130_fd_sc_hd__dfxtp_2 _40586_ (.CLK(clk),
    .D(_03080_),
    .Q(mem_addr[23]));
 sky130_fd_sc_hd__dfxtp_2 _40587_ (.CLK(clk),
    .D(_03081_),
    .Q(mem_addr[24]));
 sky130_fd_sc_hd__dfxtp_2 _40588_ (.CLK(clk),
    .D(_03082_),
    .Q(mem_addr[25]));
 sky130_fd_sc_hd__dfxtp_2 _40589_ (.CLK(clk),
    .D(_03083_),
    .Q(mem_addr[26]));
 sky130_fd_sc_hd__dfxtp_2 _40590_ (.CLK(clk),
    .D(_03084_),
    .Q(mem_addr[27]));
 sky130_fd_sc_hd__dfxtp_2 _40591_ (.CLK(clk),
    .D(_03085_),
    .Q(mem_addr[28]));
 sky130_fd_sc_hd__dfxtp_2 _40592_ (.CLK(clk),
    .D(_03086_),
    .Q(mem_addr[29]));
 sky130_fd_sc_hd__dfxtp_2 _40593_ (.CLK(clk),
    .D(_03087_),
    .Q(mem_addr[30]));
 sky130_fd_sc_hd__dfxtp_2 _40594_ (.CLK(clk),
    .D(_03088_),
    .Q(mem_addr[31]));
 sky130_fd_sc_hd__dfxtp_2 _40595_ (.CLK(clk),
    .D(_03089_),
    .Q(pcpi_rs1[0]));
 sky130_fd_sc_hd__dfxtp_2 _40596_ (.CLK(clk),
    .D(_03090_),
    .Q(pcpi_rs1[1]));
 sky130_fd_sc_hd__dfxtp_2 _40597_ (.CLK(clk),
    .D(_03091_),
    .Q(pcpi_rs1[2]));
 sky130_fd_sc_hd__dfxtp_2 _40598_ (.CLK(clk),
    .D(_03092_),
    .Q(pcpi_rs1[3]));
 sky130_fd_sc_hd__dfxtp_2 _40599_ (.CLK(clk),
    .D(_03093_),
    .Q(pcpi_rs1[4]));
 sky130_fd_sc_hd__dfxtp_2 _40600_ (.CLK(clk),
    .D(_03094_),
    .Q(pcpi_rs1[5]));
 sky130_fd_sc_hd__dfxtp_2 _40601_ (.CLK(clk),
    .D(_03095_),
    .Q(pcpi_rs1[6]));
 sky130_fd_sc_hd__dfxtp_2 _40602_ (.CLK(clk),
    .D(_03096_),
    .Q(pcpi_rs1[7]));
 sky130_fd_sc_hd__dfxtp_2 _40603_ (.CLK(clk),
    .D(_03097_),
    .Q(pcpi_rs1[8]));
 sky130_fd_sc_hd__dfxtp_2 _40604_ (.CLK(clk),
    .D(_03098_),
    .Q(pcpi_rs1[9]));
 sky130_fd_sc_hd__dfxtp_2 _40605_ (.CLK(clk),
    .D(_03099_),
    .Q(pcpi_rs1[10]));
 sky130_fd_sc_hd__dfxtp_2 _40606_ (.CLK(clk),
    .D(_03100_),
    .Q(pcpi_rs1[11]));
 sky130_fd_sc_hd__dfxtp_2 _40607_ (.CLK(clk),
    .D(_03101_),
    .Q(pcpi_rs1[12]));
 sky130_fd_sc_hd__dfxtp_2 _40608_ (.CLK(clk),
    .D(_03102_),
    .Q(pcpi_rs1[13]));
 sky130_fd_sc_hd__dfxtp_2 _40609_ (.CLK(clk),
    .D(_03103_),
    .Q(pcpi_rs1[14]));
 sky130_fd_sc_hd__dfxtp_2 _40610_ (.CLK(clk),
    .D(_03104_),
    .Q(pcpi_rs1[15]));
 sky130_fd_sc_hd__dfxtp_2 _40611_ (.CLK(clk),
    .D(_03105_),
    .Q(pcpi_rs1[16]));
 sky130_fd_sc_hd__dfxtp_2 _40612_ (.CLK(clk),
    .D(_03106_),
    .Q(pcpi_rs1[17]));
 sky130_fd_sc_hd__dfxtp_2 _40613_ (.CLK(clk),
    .D(_03107_),
    .Q(pcpi_rs1[18]));
 sky130_fd_sc_hd__dfxtp_2 _40614_ (.CLK(clk),
    .D(_03108_),
    .Q(pcpi_rs1[19]));
 sky130_fd_sc_hd__dfxtp_2 _40615_ (.CLK(clk),
    .D(_03109_),
    .Q(pcpi_rs1[20]));
 sky130_fd_sc_hd__dfxtp_2 _40616_ (.CLK(clk),
    .D(_03110_),
    .Q(pcpi_rs1[21]));
 sky130_fd_sc_hd__dfxtp_2 _40617_ (.CLK(clk),
    .D(_03111_),
    .Q(pcpi_rs1[22]));
 sky130_fd_sc_hd__dfxtp_2 _40618_ (.CLK(clk),
    .D(_03112_),
    .Q(pcpi_rs1[23]));
 sky130_fd_sc_hd__dfxtp_2 _40619_ (.CLK(clk),
    .D(_03113_),
    .Q(pcpi_rs1[24]));
 sky130_fd_sc_hd__dfxtp_2 _40620_ (.CLK(clk),
    .D(_03114_),
    .Q(pcpi_rs1[25]));
 sky130_fd_sc_hd__dfxtp_2 _40621_ (.CLK(clk),
    .D(_03115_),
    .Q(pcpi_rs1[26]));
 sky130_fd_sc_hd__dfxtp_2 _40622_ (.CLK(clk),
    .D(_03116_),
    .Q(pcpi_rs1[27]));
 sky130_fd_sc_hd__dfxtp_2 _40623_ (.CLK(clk),
    .D(_03117_),
    .Q(pcpi_rs1[28]));
 sky130_fd_sc_hd__dfxtp_2 _40624_ (.CLK(clk),
    .D(_03118_),
    .Q(pcpi_rs1[29]));
 sky130_fd_sc_hd__dfxtp_2 _40625_ (.CLK(clk),
    .D(_03119_),
    .Q(pcpi_rs1[30]));
 sky130_fd_sc_hd__dfxtp_2 _40626_ (.CLK(clk),
    .D(_03120_),
    .Q(pcpi_rs1[31]));
 sky130_fd_sc_hd__dfxtp_2 _40627_ (.CLK(clk),
    .D(_03121_),
    .Q(pcpi_insn[0]));
 sky130_fd_sc_hd__dfxtp_2 _40628_ (.CLK(clk),
    .D(_03122_),
    .Q(pcpi_insn[1]));
 sky130_fd_sc_hd__dfxtp_2 _40629_ (.CLK(clk),
    .D(_03123_),
    .Q(pcpi_insn[2]));
 sky130_fd_sc_hd__dfxtp_2 _40630_ (.CLK(clk),
    .D(_03124_),
    .Q(pcpi_insn[3]));
 sky130_fd_sc_hd__dfxtp_2 _40631_ (.CLK(clk),
    .D(_03125_),
    .Q(pcpi_insn[4]));
 sky130_fd_sc_hd__dfxtp_2 _40632_ (.CLK(clk),
    .D(_03126_),
    .Q(pcpi_insn[5]));
 sky130_fd_sc_hd__dfxtp_2 _40633_ (.CLK(clk),
    .D(_03127_),
    .Q(pcpi_insn[6]));
 sky130_fd_sc_hd__dfxtp_2 _40634_ (.CLK(clk),
    .D(_03128_),
    .Q(pcpi_insn[7]));
 sky130_fd_sc_hd__dfxtp_2 _40635_ (.CLK(clk),
    .D(_03129_),
    .Q(pcpi_insn[8]));
 sky130_fd_sc_hd__dfxtp_2 _40636_ (.CLK(clk),
    .D(_03130_),
    .Q(pcpi_insn[9]));
 sky130_fd_sc_hd__dfxtp_2 _40637_ (.CLK(clk),
    .D(_03131_),
    .Q(pcpi_insn[10]));
 sky130_fd_sc_hd__dfxtp_2 _40638_ (.CLK(clk),
    .D(_03132_),
    .Q(pcpi_insn[11]));
 sky130_fd_sc_hd__dfxtp_2 _40639_ (.CLK(clk),
    .D(_03133_),
    .Q(pcpi_insn[12]));
 sky130_fd_sc_hd__dfxtp_2 _40640_ (.CLK(clk),
    .D(_03134_),
    .Q(pcpi_insn[13]));
 sky130_fd_sc_hd__dfxtp_2 _40641_ (.CLK(clk),
    .D(_03135_),
    .Q(pcpi_insn[14]));
 sky130_fd_sc_hd__dfxtp_2 _40642_ (.CLK(clk),
    .D(_03136_),
    .Q(pcpi_insn[15]));
 sky130_fd_sc_hd__dfxtp_2 _40643_ (.CLK(clk),
    .D(_03137_),
    .Q(pcpi_insn[16]));
 sky130_fd_sc_hd__dfxtp_2 _40644_ (.CLK(clk),
    .D(_03138_),
    .Q(pcpi_insn[17]));
 sky130_fd_sc_hd__dfxtp_2 _40645_ (.CLK(clk),
    .D(_03139_),
    .Q(pcpi_insn[18]));
 sky130_fd_sc_hd__dfxtp_2 _40646_ (.CLK(clk),
    .D(_03140_),
    .Q(pcpi_insn[19]));
 sky130_fd_sc_hd__dfxtp_2 _40647_ (.CLK(clk),
    .D(_03141_),
    .Q(pcpi_insn[20]));
 sky130_fd_sc_hd__dfxtp_2 _40648_ (.CLK(clk),
    .D(_03142_),
    .Q(pcpi_insn[21]));
 sky130_fd_sc_hd__dfxtp_2 _40649_ (.CLK(clk),
    .D(_03143_),
    .Q(pcpi_insn[22]));
 sky130_fd_sc_hd__dfxtp_2 _40650_ (.CLK(clk),
    .D(_03144_),
    .Q(pcpi_insn[23]));
 sky130_fd_sc_hd__dfxtp_2 _40651_ (.CLK(clk),
    .D(_03145_),
    .Q(pcpi_insn[24]));
 sky130_fd_sc_hd__dfxtp_2 _40652_ (.CLK(clk),
    .D(_03146_),
    .Q(pcpi_insn[25]));
 sky130_fd_sc_hd__dfxtp_2 _40653_ (.CLK(clk),
    .D(_03147_),
    .Q(pcpi_insn[26]));
 sky130_fd_sc_hd__dfxtp_2 _40654_ (.CLK(clk),
    .D(_03148_),
    .Q(pcpi_insn[27]));
 sky130_fd_sc_hd__dfxtp_2 _40655_ (.CLK(clk),
    .D(_03149_),
    .Q(pcpi_insn[28]));
 sky130_fd_sc_hd__dfxtp_2 _40656_ (.CLK(clk),
    .D(_03150_),
    .Q(pcpi_insn[29]));
 sky130_fd_sc_hd__dfxtp_2 _40657_ (.CLK(clk),
    .D(_03151_),
    .Q(pcpi_insn[30]));
 sky130_fd_sc_hd__dfxtp_2 _40658_ (.CLK(clk),
    .D(_03152_),
    .Q(pcpi_insn[31]));
 sky130_fd_sc_hd__dfxtp_2 _40659_ (.CLK(clk),
    .D(_03153_),
    .Q(instr_lui));
 sky130_fd_sc_hd__dfxtp_2 _40660_ (.CLK(clk),
    .D(_03154_),
    .Q(instr_auipc));
 sky130_fd_sc_hd__dfxtp_2 _40661_ (.CLK(clk),
    .D(_03155_),
    .Q(instr_jal));
 sky130_fd_sc_hd__dfxtp_2 _40662_ (.CLK(clk),
    .D(_03156_),
    .Q(instr_jalr));
 sky130_fd_sc_hd__dfxtp_2 _40663_ (.CLK(clk),
    .D(_03157_),
    .Q(instr_lb));
 sky130_fd_sc_hd__dfxtp_2 _40664_ (.CLK(clk),
    .D(_03158_),
    .Q(instr_lh));
 sky130_fd_sc_hd__dfxtp_2 _40665_ (.CLK(clk),
    .D(_03159_),
    .Q(instr_lw));
 sky130_fd_sc_hd__dfxtp_2 _40666_ (.CLK(clk),
    .D(_03160_),
    .Q(instr_lbu));
 sky130_fd_sc_hd__dfxtp_2 _40667_ (.CLK(clk),
    .D(_03161_),
    .Q(instr_lhu));
 sky130_fd_sc_hd__dfxtp_2 _40668_ (.CLK(clk),
    .D(_03162_),
    .Q(instr_sb));
 sky130_fd_sc_hd__dfxtp_2 _40669_ (.CLK(clk),
    .D(_03163_),
    .Q(instr_sh));
 sky130_fd_sc_hd__dfxtp_2 _40670_ (.CLK(clk),
    .D(_03164_),
    .Q(instr_sw));
 sky130_fd_sc_hd__dfxtp_2 _40671_ (.CLK(clk),
    .D(_03165_),
    .Q(instr_slli));
 sky130_fd_sc_hd__dfxtp_2 _40672_ (.CLK(clk),
    .D(_03166_),
    .Q(instr_srli));
 sky130_fd_sc_hd__dfxtp_2 _40673_ (.CLK(clk),
    .D(_03167_),
    .Q(instr_srai));
 sky130_fd_sc_hd__dfxtp_2 _40674_ (.CLK(clk),
    .D(_03168_),
    .Q(instr_rdcycle));
 sky130_fd_sc_hd__dfxtp_2 _40675_ (.CLK(clk),
    .D(_03169_),
    .Q(instr_rdcycleh));
 sky130_fd_sc_hd__dfxtp_2 _40676_ (.CLK(clk),
    .D(_03170_),
    .Q(instr_rdinstr));
 sky130_fd_sc_hd__dfxtp_2 _40677_ (.CLK(clk),
    .D(_03171_),
    .Q(instr_rdinstrh));
 sky130_fd_sc_hd__dfxtp_2 _40678_ (.CLK(clk),
    .D(_03172_),
    .Q(instr_ecall_ebreak));
 sky130_fd_sc_hd__dfxtp_2 _40679_ (.CLK(clk),
    .D(_03173_),
    .Q(instr_getq));
 sky130_fd_sc_hd__dfxtp_2 _40680_ (.CLK(clk),
    .D(_03174_),
    .Q(instr_setq));
 sky130_fd_sc_hd__dfxtp_2 _40681_ (.CLK(clk),
    .D(_03175_),
    .Q(instr_retirq));
 sky130_fd_sc_hd__dfxtp_2 _40682_ (.CLK(clk),
    .D(_03176_),
    .Q(instr_maskirq));
 sky130_fd_sc_hd__dfxtp_2 _40683_ (.CLK(clk),
    .D(_03177_),
    .Q(instr_waitirq));
 sky130_fd_sc_hd__dfxtp_2 _40684_ (.CLK(clk),
    .D(_03178_),
    .Q(instr_timer));
 sky130_fd_sc_hd__dfxtp_2 _40685_ (.CLK(clk),
    .D(_03179_),
    .Q(\decoded_rd[0] ));
 sky130_fd_sc_hd__dfxtp_2 _40686_ (.CLK(clk),
    .D(_03180_),
    .Q(\decoded_rd[1] ));
 sky130_fd_sc_hd__dfxtp_2 _40687_ (.CLK(clk),
    .D(_03181_),
    .Q(\decoded_rd[2] ));
 sky130_fd_sc_hd__dfxtp_2 _40688_ (.CLK(clk),
    .D(_03182_),
    .Q(\decoded_rd[3] ));
 sky130_fd_sc_hd__dfxtp_2 _40689_ (.CLK(clk),
    .D(_03183_),
    .Q(\decoded_rd[4] ));
 sky130_fd_sc_hd__dfxtp_2 _40690_ (.CLK(clk),
    .D(_03184_),
    .Q(\decoded_imm[0] ));
 sky130_fd_sc_hd__dfxtp_2 _40691_ (.CLK(clk),
    .D(_03185_),
    .Q(\decoded_imm_uj[1] ));
 sky130_fd_sc_hd__dfxtp_2 _40692_ (.CLK(clk),
    .D(_03186_),
    .Q(\decoded_imm_uj[2] ));
 sky130_fd_sc_hd__dfxtp_2 _40693_ (.CLK(clk),
    .D(_03187_),
    .Q(\decoded_imm_uj[3] ));
 sky130_fd_sc_hd__dfxtp_2 _40694_ (.CLK(clk),
    .D(_03188_),
    .Q(\decoded_imm_uj[4] ));
 sky130_fd_sc_hd__dfxtp_2 _40695_ (.CLK(clk),
    .D(_03189_),
    .Q(\decoded_imm_uj[5] ));
 sky130_fd_sc_hd__dfxtp_2 _40696_ (.CLK(clk),
    .D(_03190_),
    .Q(\decoded_imm_uj[6] ));
 sky130_fd_sc_hd__dfxtp_2 _40697_ (.CLK(clk),
    .D(_03191_),
    .Q(\decoded_imm_uj[7] ));
 sky130_fd_sc_hd__dfxtp_2 _40698_ (.CLK(clk),
    .D(_03192_),
    .Q(\decoded_imm_uj[8] ));
 sky130_fd_sc_hd__dfxtp_2 _40699_ (.CLK(clk),
    .D(_03193_),
    .Q(\decoded_imm_uj[9] ));
 sky130_fd_sc_hd__dfxtp_2 _40700_ (.CLK(clk),
    .D(_03194_),
    .Q(\decoded_imm_uj[10] ));
 sky130_fd_sc_hd__dfxtp_2 _40701_ (.CLK(clk),
    .D(_03195_),
    .Q(\decoded_imm_uj[11] ));
 sky130_fd_sc_hd__dfxtp_2 _40702_ (.CLK(clk),
    .D(_03196_),
    .Q(\decoded_imm_uj[12] ));
 sky130_fd_sc_hd__dfxtp_2 _40703_ (.CLK(clk),
    .D(_03197_),
    .Q(\decoded_imm_uj[13] ));
 sky130_fd_sc_hd__dfxtp_2 _40704_ (.CLK(clk),
    .D(_03198_),
    .Q(\decoded_imm_uj[14] ));
 sky130_fd_sc_hd__dfxtp_2 _40705_ (.CLK(clk),
    .D(_03199_),
    .Q(\decoded_imm_uj[15] ));
 sky130_fd_sc_hd__dfxtp_2 _40706_ (.CLK(clk),
    .D(_03200_),
    .Q(\decoded_imm_uj[16] ));
 sky130_fd_sc_hd__dfxtp_2 _40707_ (.CLK(clk),
    .D(_03201_),
    .Q(\decoded_imm_uj[17] ));
 sky130_fd_sc_hd__dfxtp_2 _40708_ (.CLK(clk),
    .D(_03202_),
    .Q(\decoded_imm_uj[18] ));
 sky130_fd_sc_hd__dfxtp_2 _40709_ (.CLK(clk),
    .D(_03203_),
    .Q(\decoded_imm_uj[19] ));
 sky130_fd_sc_hd__dfxtp_2 _40710_ (.CLK(clk),
    .D(_03204_),
    .Q(\decoded_imm_uj[20] ));
 sky130_fd_sc_hd__dfxtp_2 _40711_ (.CLK(clk),
    .D(_03205_),
    .Q(is_lb_lh_lw_lbu_lhu));
 sky130_fd_sc_hd__dfxtp_2 _40712_ (.CLK(clk),
    .D(_03206_),
    .Q(is_slli_srli_srai));
 sky130_fd_sc_hd__dfxtp_2 _40713_ (.CLK(clk),
    .D(_03207_),
    .Q(is_jalr_addi_slti_sltiu_xori_ori_andi));
 sky130_fd_sc_hd__dfxtp_2 _40714_ (.CLK(clk),
    .D(_03208_),
    .Q(is_sb_sh_sw));
 sky130_fd_sc_hd__dfxtp_2 _40715_ (.CLK(clk),
    .D(_03209_),
    .Q(\cpuregs[13][0] ));
 sky130_fd_sc_hd__dfxtp_2 _40716_ (.CLK(clk),
    .D(_03210_),
    .Q(\cpuregs[13][1] ));
 sky130_fd_sc_hd__dfxtp_2 _40717_ (.CLK(clk),
    .D(_03211_),
    .Q(\cpuregs[13][2] ));
 sky130_fd_sc_hd__dfxtp_2 _40718_ (.CLK(clk),
    .D(_03212_),
    .Q(\cpuregs[13][3] ));
 sky130_fd_sc_hd__dfxtp_2 _40719_ (.CLK(clk),
    .D(_03213_),
    .Q(\cpuregs[13][4] ));
 sky130_fd_sc_hd__dfxtp_2 _40720_ (.CLK(clk),
    .D(_03214_),
    .Q(\cpuregs[13][5] ));
 sky130_fd_sc_hd__dfxtp_2 _40721_ (.CLK(clk),
    .D(_03215_),
    .Q(\cpuregs[13][6] ));
 sky130_fd_sc_hd__dfxtp_2 _40722_ (.CLK(clk),
    .D(_03216_),
    .Q(\cpuregs[13][7] ));
 sky130_fd_sc_hd__dfxtp_2 _40723_ (.CLK(clk),
    .D(_03217_),
    .Q(\cpuregs[13][8] ));
 sky130_fd_sc_hd__dfxtp_2 _40724_ (.CLK(clk),
    .D(_03218_),
    .Q(\cpuregs[13][9] ));
 sky130_fd_sc_hd__dfxtp_2 _40725_ (.CLK(clk),
    .D(_03219_),
    .Q(\cpuregs[13][10] ));
 sky130_fd_sc_hd__dfxtp_2 _40726_ (.CLK(clk),
    .D(_03220_),
    .Q(\cpuregs[13][11] ));
 sky130_fd_sc_hd__dfxtp_2 _40727_ (.CLK(clk),
    .D(_03221_),
    .Q(\cpuregs[13][12] ));
 sky130_fd_sc_hd__dfxtp_2 _40728_ (.CLK(clk),
    .D(_03222_),
    .Q(\cpuregs[13][13] ));
 sky130_fd_sc_hd__dfxtp_2 _40729_ (.CLK(clk),
    .D(_03223_),
    .Q(\cpuregs[13][14] ));
 sky130_fd_sc_hd__dfxtp_2 _40730_ (.CLK(clk),
    .D(_03224_),
    .Q(\cpuregs[13][15] ));
 sky130_fd_sc_hd__dfxtp_2 _40731_ (.CLK(clk),
    .D(_03225_),
    .Q(\cpuregs[13][16] ));
 sky130_fd_sc_hd__dfxtp_2 _40732_ (.CLK(clk),
    .D(_03226_),
    .Q(\cpuregs[13][17] ));
 sky130_fd_sc_hd__dfxtp_2 _40733_ (.CLK(clk),
    .D(_03227_),
    .Q(\cpuregs[13][18] ));
 sky130_fd_sc_hd__dfxtp_2 _40734_ (.CLK(clk),
    .D(_03228_),
    .Q(\cpuregs[13][19] ));
 sky130_fd_sc_hd__dfxtp_2 _40735_ (.CLK(clk),
    .D(_03229_),
    .Q(\cpuregs[13][20] ));
 sky130_fd_sc_hd__dfxtp_2 _40736_ (.CLK(clk),
    .D(_03230_),
    .Q(\cpuregs[13][21] ));
 sky130_fd_sc_hd__dfxtp_2 _40737_ (.CLK(clk),
    .D(_03231_),
    .Q(\cpuregs[13][22] ));
 sky130_fd_sc_hd__dfxtp_2 _40738_ (.CLK(clk),
    .D(_03232_),
    .Q(\cpuregs[13][23] ));
 sky130_fd_sc_hd__dfxtp_2 _40739_ (.CLK(clk),
    .D(_03233_),
    .Q(\cpuregs[13][24] ));
 sky130_fd_sc_hd__dfxtp_2 _40740_ (.CLK(clk),
    .D(_03234_),
    .Q(\cpuregs[13][25] ));
 sky130_fd_sc_hd__dfxtp_2 _40741_ (.CLK(clk),
    .D(_03235_),
    .Q(\cpuregs[13][26] ));
 sky130_fd_sc_hd__dfxtp_2 _40742_ (.CLK(clk),
    .D(_03236_),
    .Q(\cpuregs[13][27] ));
 sky130_fd_sc_hd__dfxtp_2 _40743_ (.CLK(clk),
    .D(_03237_),
    .Q(\cpuregs[13][28] ));
 sky130_fd_sc_hd__dfxtp_2 _40744_ (.CLK(clk),
    .D(_03238_),
    .Q(\cpuregs[13][29] ));
 sky130_fd_sc_hd__dfxtp_2 _40745_ (.CLK(clk),
    .D(_03239_),
    .Q(\cpuregs[13][30] ));
 sky130_fd_sc_hd__dfxtp_2 _40746_ (.CLK(clk),
    .D(_03240_),
    .Q(\cpuregs[13][31] ));
 sky130_fd_sc_hd__dfxtp_2 _40747_ (.CLK(clk),
    .D(_03241_),
    .Q(is_alu_reg_imm));
 sky130_fd_sc_hd__dfxtp_2 _40748_ (.CLK(clk),
    .D(_03242_),
    .Q(is_alu_reg_reg));
 sky130_fd_sc_hd__dfxtp_2 _40749_ (.CLK(clk),
    .D(_03243_),
    .Q(mem_wstrb[0]));
 sky130_fd_sc_hd__dfxtp_2 _40750_ (.CLK(clk),
    .D(_03244_),
    .Q(mem_wstrb[1]));
 sky130_fd_sc_hd__dfxtp_2 _40751_ (.CLK(clk),
    .D(_03245_),
    .Q(mem_wstrb[2]));
 sky130_fd_sc_hd__dfxtp_2 _40752_ (.CLK(clk),
    .D(_03246_),
    .Q(mem_wstrb[3]));
 sky130_fd_sc_hd__dfxtp_2 _40753_ (.CLK(clk),
    .D(_03247_),
    .Q(\pcpi_mul.rs2[0] ));
 sky130_fd_sc_hd__dfxtp_2 _40754_ (.CLK(clk),
    .D(_03248_),
    .Q(\pcpi_mul.rs2[1] ));
 sky130_fd_sc_hd__dfxtp_2 _40755_ (.CLK(clk),
    .D(_03249_),
    .Q(\pcpi_mul.rs2[2] ));
 sky130_fd_sc_hd__dfxtp_2 _40756_ (.CLK(clk),
    .D(_03250_),
    .Q(\pcpi_mul.rs2[3] ));
 sky130_fd_sc_hd__dfxtp_2 _40757_ (.CLK(clk),
    .D(_03251_),
    .Q(\pcpi_mul.rs2[4] ));
 sky130_fd_sc_hd__dfxtp_2 _40758_ (.CLK(clk),
    .D(_03252_),
    .Q(\pcpi_mul.rs2[5] ));
 sky130_fd_sc_hd__dfxtp_2 _40759_ (.CLK(clk),
    .D(_03253_),
    .Q(\pcpi_mul.rs2[6] ));
 sky130_fd_sc_hd__dfxtp_2 _40760_ (.CLK(clk),
    .D(_03254_),
    .Q(\pcpi_mul.rs2[7] ));
 sky130_fd_sc_hd__dfxtp_2 _40761_ (.CLK(clk),
    .D(_03255_),
    .Q(\pcpi_mul.rs2[8] ));
 sky130_fd_sc_hd__dfxtp_2 _40762_ (.CLK(clk),
    .D(_03256_),
    .Q(\pcpi_mul.rs2[9] ));
 sky130_fd_sc_hd__dfxtp_2 _40763_ (.CLK(clk),
    .D(_03257_),
    .Q(\pcpi_mul.rs2[10] ));
 sky130_fd_sc_hd__dfxtp_2 _40764_ (.CLK(clk),
    .D(_03258_),
    .Q(\pcpi_mul.rs2[11] ));
 sky130_fd_sc_hd__dfxtp_2 _40765_ (.CLK(clk),
    .D(_03259_),
    .Q(\pcpi_mul.rs2[12] ));
 sky130_fd_sc_hd__dfxtp_2 _40766_ (.CLK(clk),
    .D(_03260_),
    .Q(\pcpi_mul.rs2[13] ));
 sky130_fd_sc_hd__dfxtp_2 _40767_ (.CLK(clk),
    .D(_03261_),
    .Q(\pcpi_mul.rs2[14] ));
 sky130_fd_sc_hd__dfxtp_2 _40768_ (.CLK(clk),
    .D(_03262_),
    .Q(\pcpi_mul.rs2[15] ));
 sky130_fd_sc_hd__dfxtp_2 _40769_ (.CLK(clk),
    .D(_03263_),
    .Q(\pcpi_mul.rs2[16] ));
 sky130_fd_sc_hd__dfxtp_2 _40770_ (.CLK(clk),
    .D(_03264_),
    .Q(\pcpi_mul.rs2[17] ));
 sky130_fd_sc_hd__dfxtp_2 _40771_ (.CLK(clk),
    .D(_03265_),
    .Q(\pcpi_mul.rs2[18] ));
 sky130_fd_sc_hd__dfxtp_2 _40772_ (.CLK(clk),
    .D(_03266_),
    .Q(\pcpi_mul.rs2[19] ));
 sky130_fd_sc_hd__dfxtp_2 _40773_ (.CLK(clk),
    .D(_03267_),
    .Q(\pcpi_mul.rs2[20] ));
 sky130_fd_sc_hd__dfxtp_2 _40774_ (.CLK(clk),
    .D(_03268_),
    .Q(\pcpi_mul.rs2[21] ));
 sky130_fd_sc_hd__dfxtp_2 _40775_ (.CLK(clk),
    .D(_03269_),
    .Q(\pcpi_mul.rs2[22] ));
 sky130_fd_sc_hd__dfxtp_2 _40776_ (.CLK(clk),
    .D(_03270_),
    .Q(\pcpi_mul.rs2[23] ));
 sky130_fd_sc_hd__dfxtp_2 _40777_ (.CLK(clk),
    .D(_03271_),
    .Q(\pcpi_mul.rs2[24] ));
 sky130_fd_sc_hd__dfxtp_2 _40778_ (.CLK(clk),
    .D(_03272_),
    .Q(\pcpi_mul.rs2[25] ));
 sky130_fd_sc_hd__dfxtp_2 _40779_ (.CLK(clk),
    .D(_03273_),
    .Q(\pcpi_mul.rs2[26] ));
 sky130_fd_sc_hd__dfxtp_2 _40780_ (.CLK(clk),
    .D(_03274_),
    .Q(\pcpi_mul.rs2[27] ));
 sky130_fd_sc_hd__dfxtp_2 _40781_ (.CLK(clk),
    .D(_03275_),
    .Q(\pcpi_mul.rs2[28] ));
 sky130_fd_sc_hd__dfxtp_2 _40782_ (.CLK(clk),
    .D(_03276_),
    .Q(\pcpi_mul.rs2[29] ));
 sky130_fd_sc_hd__dfxtp_2 _40783_ (.CLK(clk),
    .D(_03277_),
    .Q(\pcpi_mul.rs2[30] ));
 sky130_fd_sc_hd__dfxtp_2 _40784_ (.CLK(clk),
    .D(_03278_),
    .Q(\pcpi_mul.rs2[31] ));
 sky130_fd_sc_hd__dfxtp_2 _40785_ (.CLK(clk),
    .D(_03279_),
    .Q(\cpuregs[17][0] ));
 sky130_fd_sc_hd__dfxtp_2 _40786_ (.CLK(clk),
    .D(_03280_),
    .Q(\cpuregs[17][1] ));
 sky130_fd_sc_hd__dfxtp_2 _40787_ (.CLK(clk),
    .D(_03281_),
    .Q(\cpuregs[17][2] ));
 sky130_fd_sc_hd__dfxtp_2 _40788_ (.CLK(clk),
    .D(_03282_),
    .Q(\cpuregs[17][3] ));
 sky130_fd_sc_hd__dfxtp_2 _40789_ (.CLK(clk),
    .D(_03283_),
    .Q(\cpuregs[17][4] ));
 sky130_fd_sc_hd__dfxtp_2 _40790_ (.CLK(clk),
    .D(_03284_),
    .Q(\cpuregs[17][5] ));
 sky130_fd_sc_hd__dfxtp_2 _40791_ (.CLK(clk),
    .D(_03285_),
    .Q(\cpuregs[17][6] ));
 sky130_fd_sc_hd__dfxtp_2 _40792_ (.CLK(clk),
    .D(_03286_),
    .Q(\cpuregs[17][7] ));
 sky130_fd_sc_hd__dfxtp_2 _40793_ (.CLK(clk),
    .D(_03287_),
    .Q(\cpuregs[17][8] ));
 sky130_fd_sc_hd__dfxtp_2 _40794_ (.CLK(clk),
    .D(_03288_),
    .Q(\cpuregs[17][9] ));
 sky130_fd_sc_hd__dfxtp_2 _40795_ (.CLK(clk),
    .D(_03289_),
    .Q(\cpuregs[17][10] ));
 sky130_fd_sc_hd__dfxtp_2 _40796_ (.CLK(clk),
    .D(_03290_),
    .Q(\cpuregs[17][11] ));
 sky130_fd_sc_hd__dfxtp_2 _40797_ (.CLK(clk),
    .D(_03291_),
    .Q(\cpuregs[17][12] ));
 sky130_fd_sc_hd__dfxtp_2 _40798_ (.CLK(clk),
    .D(_03292_),
    .Q(\cpuregs[17][13] ));
 sky130_fd_sc_hd__dfxtp_2 _40799_ (.CLK(clk),
    .D(_03293_),
    .Q(\cpuregs[17][14] ));
 sky130_fd_sc_hd__dfxtp_2 _40800_ (.CLK(clk),
    .D(_03294_),
    .Q(\cpuregs[17][15] ));
 sky130_fd_sc_hd__dfxtp_2 _40801_ (.CLK(clk),
    .D(_03295_),
    .Q(\cpuregs[17][16] ));
 sky130_fd_sc_hd__dfxtp_2 _40802_ (.CLK(clk),
    .D(_03296_),
    .Q(\cpuregs[17][17] ));
 sky130_fd_sc_hd__dfxtp_2 _40803_ (.CLK(clk),
    .D(_03297_),
    .Q(\cpuregs[17][18] ));
 sky130_fd_sc_hd__dfxtp_2 _40804_ (.CLK(clk),
    .D(_03298_),
    .Q(\cpuregs[17][19] ));
 sky130_fd_sc_hd__dfxtp_2 _40805_ (.CLK(clk),
    .D(_03299_),
    .Q(\cpuregs[17][20] ));
 sky130_fd_sc_hd__dfxtp_2 _40806_ (.CLK(clk),
    .D(_03300_),
    .Q(\cpuregs[17][21] ));
 sky130_fd_sc_hd__dfxtp_2 _40807_ (.CLK(clk),
    .D(_03301_),
    .Q(\cpuregs[17][22] ));
 sky130_fd_sc_hd__dfxtp_2 _40808_ (.CLK(clk),
    .D(_03302_),
    .Q(\cpuregs[17][23] ));
 sky130_fd_sc_hd__dfxtp_2 _40809_ (.CLK(clk),
    .D(_03303_),
    .Q(\cpuregs[17][24] ));
 sky130_fd_sc_hd__dfxtp_2 _40810_ (.CLK(clk),
    .D(_03304_),
    .Q(\cpuregs[17][25] ));
 sky130_fd_sc_hd__dfxtp_2 _40811_ (.CLK(clk),
    .D(_03305_),
    .Q(\cpuregs[17][26] ));
 sky130_fd_sc_hd__dfxtp_2 _40812_ (.CLK(clk),
    .D(_03306_),
    .Q(\cpuregs[17][27] ));
 sky130_fd_sc_hd__dfxtp_2 _40813_ (.CLK(clk),
    .D(_03307_),
    .Q(\cpuregs[17][28] ));
 sky130_fd_sc_hd__dfxtp_2 _40814_ (.CLK(clk),
    .D(_03308_),
    .Q(\cpuregs[17][29] ));
 sky130_fd_sc_hd__dfxtp_2 _40815_ (.CLK(clk),
    .D(_03309_),
    .Q(\cpuregs[17][30] ));
 sky130_fd_sc_hd__dfxtp_2 _40816_ (.CLK(clk),
    .D(_03310_),
    .Q(\cpuregs[17][31] ));
 sky130_fd_sc_hd__dfxtp_2 _40817_ (.CLK(clk),
    .D(_03311_),
    .Q(\cpuregs[16][0] ));
 sky130_fd_sc_hd__dfxtp_2 _40818_ (.CLK(clk),
    .D(_03312_),
    .Q(\cpuregs[16][1] ));
 sky130_fd_sc_hd__dfxtp_2 _40819_ (.CLK(clk),
    .D(_03313_),
    .Q(\cpuregs[16][2] ));
 sky130_fd_sc_hd__dfxtp_2 _40820_ (.CLK(clk),
    .D(_03314_),
    .Q(\cpuregs[16][3] ));
 sky130_fd_sc_hd__dfxtp_2 _40821_ (.CLK(clk),
    .D(_03315_),
    .Q(\cpuregs[16][4] ));
 sky130_fd_sc_hd__dfxtp_2 _40822_ (.CLK(clk),
    .D(_03316_),
    .Q(\cpuregs[16][5] ));
 sky130_fd_sc_hd__dfxtp_2 _40823_ (.CLK(clk),
    .D(_03317_),
    .Q(\cpuregs[16][6] ));
 sky130_fd_sc_hd__dfxtp_2 _40824_ (.CLK(clk),
    .D(_03318_),
    .Q(\cpuregs[16][7] ));
 sky130_fd_sc_hd__dfxtp_2 _40825_ (.CLK(clk),
    .D(_03319_),
    .Q(\cpuregs[16][8] ));
 sky130_fd_sc_hd__dfxtp_2 _40826_ (.CLK(clk),
    .D(_03320_),
    .Q(\cpuregs[16][9] ));
 sky130_fd_sc_hd__dfxtp_2 _40827_ (.CLK(clk),
    .D(_03321_),
    .Q(\cpuregs[16][10] ));
 sky130_fd_sc_hd__dfxtp_2 _40828_ (.CLK(clk),
    .D(_03322_),
    .Q(\cpuregs[16][11] ));
 sky130_fd_sc_hd__dfxtp_2 _40829_ (.CLK(clk),
    .D(_03323_),
    .Q(\cpuregs[16][12] ));
 sky130_fd_sc_hd__dfxtp_2 _40830_ (.CLK(clk),
    .D(_03324_),
    .Q(\cpuregs[16][13] ));
 sky130_fd_sc_hd__dfxtp_2 _40831_ (.CLK(clk),
    .D(_03325_),
    .Q(\cpuregs[16][14] ));
 sky130_fd_sc_hd__dfxtp_2 _40832_ (.CLK(clk),
    .D(_03326_),
    .Q(\cpuregs[16][15] ));
 sky130_fd_sc_hd__dfxtp_2 _40833_ (.CLK(clk),
    .D(_03327_),
    .Q(\cpuregs[16][16] ));
 sky130_fd_sc_hd__dfxtp_2 _40834_ (.CLK(clk),
    .D(_03328_),
    .Q(\cpuregs[16][17] ));
 sky130_fd_sc_hd__dfxtp_2 _40835_ (.CLK(clk),
    .D(_03329_),
    .Q(\cpuregs[16][18] ));
 sky130_fd_sc_hd__dfxtp_2 _40836_ (.CLK(clk),
    .D(_03330_),
    .Q(\cpuregs[16][19] ));
 sky130_fd_sc_hd__dfxtp_2 _40837_ (.CLK(clk),
    .D(_03331_),
    .Q(\cpuregs[16][20] ));
 sky130_fd_sc_hd__dfxtp_2 _40838_ (.CLK(clk),
    .D(_03332_),
    .Q(\cpuregs[16][21] ));
 sky130_fd_sc_hd__dfxtp_2 _40839_ (.CLK(clk),
    .D(_03333_),
    .Q(\cpuregs[16][22] ));
 sky130_fd_sc_hd__dfxtp_2 _40840_ (.CLK(clk),
    .D(_03334_),
    .Q(\cpuregs[16][23] ));
 sky130_fd_sc_hd__dfxtp_2 _40841_ (.CLK(clk),
    .D(_03335_),
    .Q(\cpuregs[16][24] ));
 sky130_fd_sc_hd__dfxtp_2 _40842_ (.CLK(clk),
    .D(_03336_),
    .Q(\cpuregs[16][25] ));
 sky130_fd_sc_hd__dfxtp_2 _40843_ (.CLK(clk),
    .D(_03337_),
    .Q(\cpuregs[16][26] ));
 sky130_fd_sc_hd__dfxtp_2 _40844_ (.CLK(clk),
    .D(_03338_),
    .Q(\cpuregs[16][27] ));
 sky130_fd_sc_hd__dfxtp_2 _40845_ (.CLK(clk),
    .D(_03339_),
    .Q(\cpuregs[16][28] ));
 sky130_fd_sc_hd__dfxtp_2 _40846_ (.CLK(clk),
    .D(_03340_),
    .Q(\cpuregs[16][29] ));
 sky130_fd_sc_hd__dfxtp_2 _40847_ (.CLK(clk),
    .D(_03341_),
    .Q(\cpuregs[16][30] ));
 sky130_fd_sc_hd__dfxtp_2 _40848_ (.CLK(clk),
    .D(_03342_),
    .Q(\cpuregs[16][31] ));
 sky130_fd_sc_hd__dfxtp_2 _40849_ (.CLK(clk),
    .D(_03343_),
    .Q(\cpuregs[12][0] ));
 sky130_fd_sc_hd__dfxtp_2 _40850_ (.CLK(clk),
    .D(_03344_),
    .Q(\cpuregs[12][1] ));
 sky130_fd_sc_hd__dfxtp_2 _40851_ (.CLK(clk),
    .D(_03345_),
    .Q(\cpuregs[12][2] ));
 sky130_fd_sc_hd__dfxtp_2 _40852_ (.CLK(clk),
    .D(_03346_),
    .Q(\cpuregs[12][3] ));
 sky130_fd_sc_hd__dfxtp_2 _40853_ (.CLK(clk),
    .D(_03347_),
    .Q(\cpuregs[12][4] ));
 sky130_fd_sc_hd__dfxtp_2 _40854_ (.CLK(clk),
    .D(_03348_),
    .Q(\cpuregs[12][5] ));
 sky130_fd_sc_hd__dfxtp_2 _40855_ (.CLK(clk),
    .D(_03349_),
    .Q(\cpuregs[12][6] ));
 sky130_fd_sc_hd__dfxtp_2 _40856_ (.CLK(clk),
    .D(_03350_),
    .Q(\cpuregs[12][7] ));
 sky130_fd_sc_hd__dfxtp_2 _40857_ (.CLK(clk),
    .D(_03351_),
    .Q(\cpuregs[12][8] ));
 sky130_fd_sc_hd__dfxtp_2 _40858_ (.CLK(clk),
    .D(_03352_),
    .Q(\cpuregs[12][9] ));
 sky130_fd_sc_hd__dfxtp_2 _40859_ (.CLK(clk),
    .D(_03353_),
    .Q(\cpuregs[12][10] ));
 sky130_fd_sc_hd__dfxtp_2 _40860_ (.CLK(clk),
    .D(_03354_),
    .Q(\cpuregs[12][11] ));
 sky130_fd_sc_hd__dfxtp_2 _40861_ (.CLK(clk),
    .D(_03355_),
    .Q(\cpuregs[12][12] ));
 sky130_fd_sc_hd__dfxtp_2 _40862_ (.CLK(clk),
    .D(_03356_),
    .Q(\cpuregs[12][13] ));
 sky130_fd_sc_hd__dfxtp_2 _40863_ (.CLK(clk),
    .D(_03357_),
    .Q(\cpuregs[12][14] ));
 sky130_fd_sc_hd__dfxtp_2 _40864_ (.CLK(clk),
    .D(_03358_),
    .Q(\cpuregs[12][15] ));
 sky130_fd_sc_hd__dfxtp_2 _40865_ (.CLK(clk),
    .D(_03359_),
    .Q(\cpuregs[12][16] ));
 sky130_fd_sc_hd__dfxtp_2 _40866_ (.CLK(clk),
    .D(_03360_),
    .Q(\cpuregs[12][17] ));
 sky130_fd_sc_hd__dfxtp_2 _40867_ (.CLK(clk),
    .D(_03361_),
    .Q(\cpuregs[12][18] ));
 sky130_fd_sc_hd__dfxtp_2 _40868_ (.CLK(clk),
    .D(_03362_),
    .Q(\cpuregs[12][19] ));
 sky130_fd_sc_hd__dfxtp_2 _40869_ (.CLK(clk),
    .D(_03363_),
    .Q(\cpuregs[12][20] ));
 sky130_fd_sc_hd__dfxtp_2 _40870_ (.CLK(clk),
    .D(_03364_),
    .Q(\cpuregs[12][21] ));
 sky130_fd_sc_hd__dfxtp_2 _40871_ (.CLK(clk),
    .D(_03365_),
    .Q(\cpuregs[12][22] ));
 sky130_fd_sc_hd__dfxtp_2 _40872_ (.CLK(clk),
    .D(_03366_),
    .Q(\cpuregs[12][23] ));
 sky130_fd_sc_hd__dfxtp_2 _40873_ (.CLK(clk),
    .D(_03367_),
    .Q(\cpuregs[12][24] ));
 sky130_fd_sc_hd__dfxtp_2 _40874_ (.CLK(clk),
    .D(_03368_),
    .Q(\cpuregs[12][25] ));
 sky130_fd_sc_hd__dfxtp_2 _40875_ (.CLK(clk),
    .D(_03369_),
    .Q(\cpuregs[12][26] ));
 sky130_fd_sc_hd__dfxtp_2 _40876_ (.CLK(clk),
    .D(_03370_),
    .Q(\cpuregs[12][27] ));
 sky130_fd_sc_hd__dfxtp_2 _40877_ (.CLK(clk),
    .D(_03371_),
    .Q(\cpuregs[12][28] ));
 sky130_fd_sc_hd__dfxtp_2 _40878_ (.CLK(clk),
    .D(_03372_),
    .Q(\cpuregs[12][29] ));
 sky130_fd_sc_hd__dfxtp_2 _40879_ (.CLK(clk),
    .D(_03373_),
    .Q(\cpuregs[12][30] ));
 sky130_fd_sc_hd__dfxtp_2 _40880_ (.CLK(clk),
    .D(_03374_),
    .Q(\cpuregs[12][31] ));
 sky130_fd_sc_hd__dfxtp_2 _40881_ (.CLK(clk),
    .D(_03375_),
    .Q(\cpuregs[1][0] ));
 sky130_fd_sc_hd__dfxtp_2 _40882_ (.CLK(clk),
    .D(_03376_),
    .Q(\cpuregs[1][1] ));
 sky130_fd_sc_hd__dfxtp_2 _40883_ (.CLK(clk),
    .D(_03377_),
    .Q(\cpuregs[1][2] ));
 sky130_fd_sc_hd__dfxtp_2 _40884_ (.CLK(clk),
    .D(_03378_),
    .Q(\cpuregs[1][3] ));
 sky130_fd_sc_hd__dfxtp_2 _40885_ (.CLK(clk),
    .D(_03379_),
    .Q(\cpuregs[1][4] ));
 sky130_fd_sc_hd__dfxtp_2 _40886_ (.CLK(clk),
    .D(_03380_),
    .Q(\cpuregs[1][5] ));
 sky130_fd_sc_hd__dfxtp_2 _40887_ (.CLK(clk),
    .D(_03381_),
    .Q(\cpuregs[1][6] ));
 sky130_fd_sc_hd__dfxtp_2 _40888_ (.CLK(clk),
    .D(_03382_),
    .Q(\cpuregs[1][7] ));
 sky130_fd_sc_hd__dfxtp_2 _40889_ (.CLK(clk),
    .D(_03383_),
    .Q(\cpuregs[1][8] ));
 sky130_fd_sc_hd__dfxtp_2 _40890_ (.CLK(clk),
    .D(_03384_),
    .Q(\cpuregs[1][9] ));
 sky130_fd_sc_hd__dfxtp_2 _40891_ (.CLK(clk),
    .D(_03385_),
    .Q(\cpuregs[1][10] ));
 sky130_fd_sc_hd__dfxtp_2 _40892_ (.CLK(clk),
    .D(_03386_),
    .Q(\cpuregs[1][11] ));
 sky130_fd_sc_hd__dfxtp_2 _40893_ (.CLK(clk),
    .D(_03387_),
    .Q(\cpuregs[1][12] ));
 sky130_fd_sc_hd__dfxtp_2 _40894_ (.CLK(clk),
    .D(_03388_),
    .Q(\cpuregs[1][13] ));
 sky130_fd_sc_hd__dfxtp_2 _40895_ (.CLK(clk),
    .D(_03389_),
    .Q(\cpuregs[1][14] ));
 sky130_fd_sc_hd__dfxtp_2 _40896_ (.CLK(clk),
    .D(_03390_),
    .Q(\cpuregs[1][15] ));
 sky130_fd_sc_hd__dfxtp_2 _40897_ (.CLK(clk),
    .D(_03391_),
    .Q(\cpuregs[1][16] ));
 sky130_fd_sc_hd__dfxtp_2 _40898_ (.CLK(clk),
    .D(_03392_),
    .Q(\cpuregs[1][17] ));
 sky130_fd_sc_hd__dfxtp_2 _40899_ (.CLK(clk),
    .D(_03393_),
    .Q(\cpuregs[1][18] ));
 sky130_fd_sc_hd__dfxtp_2 _40900_ (.CLK(clk),
    .D(_03394_),
    .Q(\cpuregs[1][19] ));
 sky130_fd_sc_hd__dfxtp_2 _40901_ (.CLK(clk),
    .D(_03395_),
    .Q(\cpuregs[1][20] ));
 sky130_fd_sc_hd__dfxtp_2 _40902_ (.CLK(clk),
    .D(_03396_),
    .Q(\cpuregs[1][21] ));
 sky130_fd_sc_hd__dfxtp_2 _40903_ (.CLK(clk),
    .D(_03397_),
    .Q(\cpuregs[1][22] ));
 sky130_fd_sc_hd__dfxtp_2 _40904_ (.CLK(clk),
    .D(_03398_),
    .Q(\cpuregs[1][23] ));
 sky130_fd_sc_hd__dfxtp_2 _40905_ (.CLK(clk),
    .D(_03399_),
    .Q(\cpuregs[1][24] ));
 sky130_fd_sc_hd__dfxtp_2 _40906_ (.CLK(clk),
    .D(_03400_),
    .Q(\cpuregs[1][25] ));
 sky130_fd_sc_hd__dfxtp_2 _40907_ (.CLK(clk),
    .D(_03401_),
    .Q(\cpuregs[1][26] ));
 sky130_fd_sc_hd__dfxtp_2 _40908_ (.CLK(clk),
    .D(_03402_),
    .Q(\cpuregs[1][27] ));
 sky130_fd_sc_hd__dfxtp_2 _40909_ (.CLK(clk),
    .D(_03403_),
    .Q(\cpuregs[1][28] ));
 sky130_fd_sc_hd__dfxtp_2 _40910_ (.CLK(clk),
    .D(_03404_),
    .Q(\cpuregs[1][29] ));
 sky130_fd_sc_hd__dfxtp_2 _40911_ (.CLK(clk),
    .D(_03405_),
    .Q(\cpuregs[1][30] ));
 sky130_fd_sc_hd__dfxtp_2 _40912_ (.CLK(clk),
    .D(_03406_),
    .Q(\cpuregs[1][31] ));
 sky130_fd_sc_hd__dfxtp_2 _40913_ (.CLK(clk),
    .D(_03407_),
    .Q(\cpuregs[3][0] ));
 sky130_fd_sc_hd__dfxtp_2 _40914_ (.CLK(clk),
    .D(_03408_),
    .Q(\cpuregs[3][1] ));
 sky130_fd_sc_hd__dfxtp_2 _40915_ (.CLK(clk),
    .D(_03409_),
    .Q(\cpuregs[3][2] ));
 sky130_fd_sc_hd__dfxtp_2 _40916_ (.CLK(clk),
    .D(_03410_),
    .Q(\cpuregs[3][3] ));
 sky130_fd_sc_hd__dfxtp_2 _40917_ (.CLK(clk),
    .D(_03411_),
    .Q(\cpuregs[3][4] ));
 sky130_fd_sc_hd__dfxtp_2 _40918_ (.CLK(clk),
    .D(_03412_),
    .Q(\cpuregs[3][5] ));
 sky130_fd_sc_hd__dfxtp_2 _40919_ (.CLK(clk),
    .D(_03413_),
    .Q(\cpuregs[3][6] ));
 sky130_fd_sc_hd__dfxtp_2 _40920_ (.CLK(clk),
    .D(_03414_),
    .Q(\cpuregs[3][7] ));
 sky130_fd_sc_hd__dfxtp_2 _40921_ (.CLK(clk),
    .D(_03415_),
    .Q(\cpuregs[3][8] ));
 sky130_fd_sc_hd__dfxtp_2 _40922_ (.CLK(clk),
    .D(_03416_),
    .Q(\cpuregs[3][9] ));
 sky130_fd_sc_hd__dfxtp_2 _40923_ (.CLK(clk),
    .D(_03417_),
    .Q(\cpuregs[3][10] ));
 sky130_fd_sc_hd__dfxtp_2 _40924_ (.CLK(clk),
    .D(_03418_),
    .Q(\cpuregs[3][11] ));
 sky130_fd_sc_hd__dfxtp_2 _40925_ (.CLK(clk),
    .D(_03419_),
    .Q(\cpuregs[3][12] ));
 sky130_fd_sc_hd__dfxtp_2 _40926_ (.CLK(clk),
    .D(_03420_),
    .Q(\cpuregs[3][13] ));
 sky130_fd_sc_hd__dfxtp_2 _40927_ (.CLK(clk),
    .D(_03421_),
    .Q(\cpuregs[3][14] ));
 sky130_fd_sc_hd__dfxtp_2 _40928_ (.CLK(clk),
    .D(_03422_),
    .Q(\cpuregs[3][15] ));
 sky130_fd_sc_hd__dfxtp_2 _40929_ (.CLK(clk),
    .D(_03423_),
    .Q(\cpuregs[3][16] ));
 sky130_fd_sc_hd__dfxtp_2 _40930_ (.CLK(clk),
    .D(_03424_),
    .Q(\cpuregs[3][17] ));
 sky130_fd_sc_hd__dfxtp_2 _40931_ (.CLK(clk),
    .D(_03425_),
    .Q(\cpuregs[3][18] ));
 sky130_fd_sc_hd__dfxtp_2 _40932_ (.CLK(clk),
    .D(_03426_),
    .Q(\cpuregs[3][19] ));
 sky130_fd_sc_hd__dfxtp_2 _40933_ (.CLK(clk),
    .D(_03427_),
    .Q(\cpuregs[3][20] ));
 sky130_fd_sc_hd__dfxtp_2 _40934_ (.CLK(clk),
    .D(_03428_),
    .Q(\cpuregs[3][21] ));
 sky130_fd_sc_hd__dfxtp_2 _40935_ (.CLK(clk),
    .D(_03429_),
    .Q(\cpuregs[3][22] ));
 sky130_fd_sc_hd__dfxtp_2 _40936_ (.CLK(clk),
    .D(_03430_),
    .Q(\cpuregs[3][23] ));
 sky130_fd_sc_hd__dfxtp_2 _40937_ (.CLK(clk),
    .D(_03431_),
    .Q(\cpuregs[3][24] ));
 sky130_fd_sc_hd__dfxtp_2 _40938_ (.CLK(clk),
    .D(_03432_),
    .Q(\cpuregs[3][25] ));
 sky130_fd_sc_hd__dfxtp_2 _40939_ (.CLK(clk),
    .D(_03433_),
    .Q(\cpuregs[3][26] ));
 sky130_fd_sc_hd__dfxtp_2 _40940_ (.CLK(clk),
    .D(_03434_),
    .Q(\cpuregs[3][27] ));
 sky130_fd_sc_hd__dfxtp_2 _40941_ (.CLK(clk),
    .D(_03435_),
    .Q(\cpuregs[3][28] ));
 sky130_fd_sc_hd__dfxtp_2 _40942_ (.CLK(clk),
    .D(_03436_),
    .Q(\cpuregs[3][29] ));
 sky130_fd_sc_hd__dfxtp_2 _40943_ (.CLK(clk),
    .D(_03437_),
    .Q(\cpuregs[3][30] ));
 sky130_fd_sc_hd__dfxtp_2 _40944_ (.CLK(clk),
    .D(_03438_),
    .Q(\cpuregs[3][31] ));
 sky130_fd_sc_hd__dfxtp_2 _40945_ (.CLK(clk),
    .D(_03439_),
    .Q(\cpuregs[11][0] ));
 sky130_fd_sc_hd__dfxtp_2 _40946_ (.CLK(clk),
    .D(_03440_),
    .Q(\cpuregs[11][1] ));
 sky130_fd_sc_hd__dfxtp_2 _40947_ (.CLK(clk),
    .D(_03441_),
    .Q(\cpuregs[11][2] ));
 sky130_fd_sc_hd__dfxtp_2 _40948_ (.CLK(clk),
    .D(_03442_),
    .Q(\cpuregs[11][3] ));
 sky130_fd_sc_hd__dfxtp_2 _40949_ (.CLK(clk),
    .D(_03443_),
    .Q(\cpuregs[11][4] ));
 sky130_fd_sc_hd__dfxtp_2 _40950_ (.CLK(clk),
    .D(_03444_),
    .Q(\cpuregs[11][5] ));
 sky130_fd_sc_hd__dfxtp_2 _40951_ (.CLK(clk),
    .D(_03445_),
    .Q(\cpuregs[11][6] ));
 sky130_fd_sc_hd__dfxtp_2 _40952_ (.CLK(clk),
    .D(_03446_),
    .Q(\cpuregs[11][7] ));
 sky130_fd_sc_hd__dfxtp_2 _40953_ (.CLK(clk),
    .D(_03447_),
    .Q(\cpuregs[11][8] ));
 sky130_fd_sc_hd__dfxtp_2 _40954_ (.CLK(clk),
    .D(_03448_),
    .Q(\cpuregs[11][9] ));
 sky130_fd_sc_hd__dfxtp_2 _40955_ (.CLK(clk),
    .D(_03449_),
    .Q(\cpuregs[11][10] ));
 sky130_fd_sc_hd__dfxtp_2 _40956_ (.CLK(clk),
    .D(_03450_),
    .Q(\cpuregs[11][11] ));
 sky130_fd_sc_hd__dfxtp_2 _40957_ (.CLK(clk),
    .D(_03451_),
    .Q(\cpuregs[11][12] ));
 sky130_fd_sc_hd__dfxtp_2 _40958_ (.CLK(clk),
    .D(_03452_),
    .Q(\cpuregs[11][13] ));
 sky130_fd_sc_hd__dfxtp_2 _40959_ (.CLK(clk),
    .D(_03453_),
    .Q(\cpuregs[11][14] ));
 sky130_fd_sc_hd__dfxtp_2 _40960_ (.CLK(clk),
    .D(_03454_),
    .Q(\cpuregs[11][15] ));
 sky130_fd_sc_hd__dfxtp_2 _40961_ (.CLK(clk),
    .D(_03455_),
    .Q(\cpuregs[11][16] ));
 sky130_fd_sc_hd__dfxtp_2 _40962_ (.CLK(clk),
    .D(_03456_),
    .Q(\cpuregs[11][17] ));
 sky130_fd_sc_hd__dfxtp_2 _40963_ (.CLK(clk),
    .D(_03457_),
    .Q(\cpuregs[11][18] ));
 sky130_fd_sc_hd__dfxtp_2 _40964_ (.CLK(clk),
    .D(_03458_),
    .Q(\cpuregs[11][19] ));
 sky130_fd_sc_hd__dfxtp_2 _40965_ (.CLK(clk),
    .D(_03459_),
    .Q(\cpuregs[11][20] ));
 sky130_fd_sc_hd__dfxtp_2 _40966_ (.CLK(clk),
    .D(_03460_),
    .Q(\cpuregs[11][21] ));
 sky130_fd_sc_hd__dfxtp_2 _40967_ (.CLK(clk),
    .D(_03461_),
    .Q(\cpuregs[11][22] ));
 sky130_fd_sc_hd__dfxtp_2 _40968_ (.CLK(clk),
    .D(_03462_),
    .Q(\cpuregs[11][23] ));
 sky130_fd_sc_hd__dfxtp_2 _40969_ (.CLK(clk),
    .D(_03463_),
    .Q(\cpuregs[11][24] ));
 sky130_fd_sc_hd__dfxtp_2 _40970_ (.CLK(clk),
    .D(_03464_),
    .Q(\cpuregs[11][25] ));
 sky130_fd_sc_hd__dfxtp_2 _40971_ (.CLK(clk),
    .D(_03465_),
    .Q(\cpuregs[11][26] ));
 sky130_fd_sc_hd__dfxtp_2 _40972_ (.CLK(clk),
    .D(_03466_),
    .Q(\cpuregs[11][27] ));
 sky130_fd_sc_hd__dfxtp_2 _40973_ (.CLK(clk),
    .D(_03467_),
    .Q(\cpuregs[11][28] ));
 sky130_fd_sc_hd__dfxtp_2 _40974_ (.CLK(clk),
    .D(_03468_),
    .Q(\cpuregs[11][29] ));
 sky130_fd_sc_hd__dfxtp_2 _40975_ (.CLK(clk),
    .D(_03469_),
    .Q(\cpuregs[11][30] ));
 sky130_fd_sc_hd__dfxtp_2 _40976_ (.CLK(clk),
    .D(_03470_),
    .Q(\cpuregs[11][31] ));
 sky130_fd_sc_hd__dfxtp_2 _40977_ (.CLK(clk),
    .D(_03471_),
    .Q(\cpuregs[15][0] ));
 sky130_fd_sc_hd__dfxtp_2 _40978_ (.CLK(clk),
    .D(_03472_),
    .Q(\cpuregs[15][1] ));
 sky130_fd_sc_hd__dfxtp_2 _40979_ (.CLK(clk),
    .D(_03473_),
    .Q(\cpuregs[15][2] ));
 sky130_fd_sc_hd__dfxtp_2 _40980_ (.CLK(clk),
    .D(_03474_),
    .Q(\cpuregs[15][3] ));
 sky130_fd_sc_hd__dfxtp_2 _40981_ (.CLK(clk),
    .D(_03475_),
    .Q(\cpuregs[15][4] ));
 sky130_fd_sc_hd__dfxtp_2 _40982_ (.CLK(clk),
    .D(_03476_),
    .Q(\cpuregs[15][5] ));
 sky130_fd_sc_hd__dfxtp_2 _40983_ (.CLK(clk),
    .D(_03477_),
    .Q(\cpuregs[15][6] ));
 sky130_fd_sc_hd__dfxtp_2 _40984_ (.CLK(clk),
    .D(_03478_),
    .Q(\cpuregs[15][7] ));
 sky130_fd_sc_hd__dfxtp_2 _40985_ (.CLK(clk),
    .D(_03479_),
    .Q(\cpuregs[15][8] ));
 sky130_fd_sc_hd__dfxtp_2 _40986_ (.CLK(clk),
    .D(_03480_),
    .Q(\cpuregs[15][9] ));
 sky130_fd_sc_hd__dfxtp_2 _40987_ (.CLK(clk),
    .D(_03481_),
    .Q(\cpuregs[15][10] ));
 sky130_fd_sc_hd__dfxtp_2 _40988_ (.CLK(clk),
    .D(_03482_),
    .Q(\cpuregs[15][11] ));
 sky130_fd_sc_hd__dfxtp_2 _40989_ (.CLK(clk),
    .D(_03483_),
    .Q(\cpuregs[15][12] ));
 sky130_fd_sc_hd__dfxtp_2 _40990_ (.CLK(clk),
    .D(_03484_),
    .Q(\cpuregs[15][13] ));
 sky130_fd_sc_hd__dfxtp_2 _40991_ (.CLK(clk),
    .D(_03485_),
    .Q(\cpuregs[15][14] ));
 sky130_fd_sc_hd__dfxtp_2 _40992_ (.CLK(clk),
    .D(_03486_),
    .Q(\cpuregs[15][15] ));
 sky130_fd_sc_hd__dfxtp_2 _40993_ (.CLK(clk),
    .D(_03487_),
    .Q(\cpuregs[15][16] ));
 sky130_fd_sc_hd__dfxtp_2 _40994_ (.CLK(clk),
    .D(_03488_),
    .Q(\cpuregs[15][17] ));
 sky130_fd_sc_hd__dfxtp_2 _40995_ (.CLK(clk),
    .D(_03489_),
    .Q(\cpuregs[15][18] ));
 sky130_fd_sc_hd__dfxtp_2 _40996_ (.CLK(clk),
    .D(_03490_),
    .Q(\cpuregs[15][19] ));
 sky130_fd_sc_hd__dfxtp_2 _40997_ (.CLK(clk),
    .D(_03491_),
    .Q(\cpuregs[15][20] ));
 sky130_fd_sc_hd__dfxtp_2 _40998_ (.CLK(clk),
    .D(_03492_),
    .Q(\cpuregs[15][21] ));
 sky130_fd_sc_hd__dfxtp_2 _40999_ (.CLK(clk),
    .D(_03493_),
    .Q(\cpuregs[15][22] ));
 sky130_fd_sc_hd__dfxtp_2 _41000_ (.CLK(clk),
    .D(_03494_),
    .Q(\cpuregs[15][23] ));
 sky130_fd_sc_hd__dfxtp_2 _41001_ (.CLK(clk),
    .D(_03495_),
    .Q(\cpuregs[15][24] ));
 sky130_fd_sc_hd__dfxtp_2 _41002_ (.CLK(clk),
    .D(_03496_),
    .Q(\cpuregs[15][25] ));
 sky130_fd_sc_hd__dfxtp_2 _41003_ (.CLK(clk),
    .D(_03497_),
    .Q(\cpuregs[15][26] ));
 sky130_fd_sc_hd__dfxtp_2 _41004_ (.CLK(clk),
    .D(_03498_),
    .Q(\cpuregs[15][27] ));
 sky130_fd_sc_hd__dfxtp_2 _41005_ (.CLK(clk),
    .D(_03499_),
    .Q(\cpuregs[15][28] ));
 sky130_fd_sc_hd__dfxtp_2 _41006_ (.CLK(clk),
    .D(_03500_),
    .Q(\cpuregs[15][29] ));
 sky130_fd_sc_hd__dfxtp_2 _41007_ (.CLK(clk),
    .D(_03501_),
    .Q(\cpuregs[15][30] ));
 sky130_fd_sc_hd__dfxtp_2 _41008_ (.CLK(clk),
    .D(_03502_),
    .Q(\cpuregs[15][31] ));
 sky130_fd_sc_hd__dfxtp_2 _41009_ (.CLK(clk),
    .D(_03503_),
    .Q(\latched_rd[4] ));
 sky130_fd_sc_hd__dfxtp_2 _41010_ (.CLK(clk),
    .D(_03504_),
    .Q(\cpuregs[7][0] ));
 sky130_fd_sc_hd__dfxtp_2 _41011_ (.CLK(clk),
    .D(_03505_),
    .Q(\cpuregs[7][1] ));
 sky130_fd_sc_hd__dfxtp_2 _41012_ (.CLK(clk),
    .D(_03506_),
    .Q(\cpuregs[7][2] ));
 sky130_fd_sc_hd__dfxtp_2 _41013_ (.CLK(clk),
    .D(_03507_),
    .Q(\cpuregs[7][3] ));
 sky130_fd_sc_hd__dfxtp_2 _41014_ (.CLK(clk),
    .D(_03508_),
    .Q(\cpuregs[7][4] ));
 sky130_fd_sc_hd__dfxtp_2 _41015_ (.CLK(clk),
    .D(_03509_),
    .Q(\cpuregs[7][5] ));
 sky130_fd_sc_hd__dfxtp_2 _41016_ (.CLK(clk),
    .D(_03510_),
    .Q(\cpuregs[7][6] ));
 sky130_fd_sc_hd__dfxtp_2 _41017_ (.CLK(clk),
    .D(_03511_),
    .Q(\cpuregs[7][7] ));
 sky130_fd_sc_hd__dfxtp_2 _41018_ (.CLK(clk),
    .D(_03512_),
    .Q(\cpuregs[7][8] ));
 sky130_fd_sc_hd__dfxtp_2 _41019_ (.CLK(clk),
    .D(_03513_),
    .Q(\cpuregs[7][9] ));
 sky130_fd_sc_hd__dfxtp_2 _41020_ (.CLK(clk),
    .D(_03514_),
    .Q(\cpuregs[7][10] ));
 sky130_fd_sc_hd__dfxtp_2 _41021_ (.CLK(clk),
    .D(_03515_),
    .Q(\cpuregs[7][11] ));
 sky130_fd_sc_hd__dfxtp_2 _41022_ (.CLK(clk),
    .D(_03516_),
    .Q(\cpuregs[7][12] ));
 sky130_fd_sc_hd__dfxtp_2 _41023_ (.CLK(clk),
    .D(_03517_),
    .Q(\cpuregs[7][13] ));
 sky130_fd_sc_hd__dfxtp_2 _41024_ (.CLK(clk),
    .D(_03518_),
    .Q(\cpuregs[7][14] ));
 sky130_fd_sc_hd__dfxtp_2 _41025_ (.CLK(clk),
    .D(_03519_),
    .Q(\cpuregs[7][15] ));
 sky130_fd_sc_hd__dfxtp_2 _41026_ (.CLK(clk),
    .D(_03520_),
    .Q(\cpuregs[7][16] ));
 sky130_fd_sc_hd__dfxtp_2 _41027_ (.CLK(clk),
    .D(_03521_),
    .Q(\cpuregs[7][17] ));
 sky130_fd_sc_hd__dfxtp_2 _41028_ (.CLK(clk),
    .D(_03522_),
    .Q(\cpuregs[7][18] ));
 sky130_fd_sc_hd__dfxtp_2 _41029_ (.CLK(clk),
    .D(_03523_),
    .Q(\cpuregs[7][19] ));
 sky130_fd_sc_hd__dfxtp_2 _41030_ (.CLK(clk),
    .D(_03524_),
    .Q(\cpuregs[7][20] ));
 sky130_fd_sc_hd__dfxtp_2 _41031_ (.CLK(clk),
    .D(_03525_),
    .Q(\cpuregs[7][21] ));
 sky130_fd_sc_hd__dfxtp_2 _41032_ (.CLK(clk),
    .D(_03526_),
    .Q(\cpuregs[7][22] ));
 sky130_fd_sc_hd__dfxtp_2 _41033_ (.CLK(clk),
    .D(_03527_),
    .Q(\cpuregs[7][23] ));
 sky130_fd_sc_hd__dfxtp_2 _41034_ (.CLK(clk),
    .D(_03528_),
    .Q(\cpuregs[7][24] ));
 sky130_fd_sc_hd__dfxtp_2 _41035_ (.CLK(clk),
    .D(_03529_),
    .Q(\cpuregs[7][25] ));
 sky130_fd_sc_hd__dfxtp_2 _41036_ (.CLK(clk),
    .D(_03530_),
    .Q(\cpuregs[7][26] ));
 sky130_fd_sc_hd__dfxtp_2 _41037_ (.CLK(clk),
    .D(_03531_),
    .Q(\cpuregs[7][27] ));
 sky130_fd_sc_hd__dfxtp_2 _41038_ (.CLK(clk),
    .D(_03532_),
    .Q(\cpuregs[7][28] ));
 sky130_fd_sc_hd__dfxtp_2 _41039_ (.CLK(clk),
    .D(_03533_),
    .Q(\cpuregs[7][29] ));
 sky130_fd_sc_hd__dfxtp_2 _41040_ (.CLK(clk),
    .D(_03534_),
    .Q(\cpuregs[7][30] ));
 sky130_fd_sc_hd__dfxtp_2 _41041_ (.CLK(clk),
    .D(_03535_),
    .Q(\cpuregs[7][31] ));
 sky130_fd_sc_hd__dfxtp_2 _41042_ (.CLK(clk),
    .D(_03536_),
    .Q(mem_wdata[0]));
 sky130_fd_sc_hd__dfxtp_2 _41043_ (.CLK(clk),
    .D(_03537_),
    .Q(mem_wdata[1]));
 sky130_fd_sc_hd__dfxtp_2 _41044_ (.CLK(clk),
    .D(_03538_),
    .Q(mem_wdata[2]));
 sky130_fd_sc_hd__dfxtp_2 _41045_ (.CLK(clk),
    .D(_03539_),
    .Q(mem_wdata[3]));
 sky130_fd_sc_hd__dfxtp_2 _41046_ (.CLK(clk),
    .D(_03540_),
    .Q(mem_wdata[4]));
 sky130_fd_sc_hd__dfxtp_2 _41047_ (.CLK(clk),
    .D(_03541_),
    .Q(mem_wdata[5]));
 sky130_fd_sc_hd__dfxtp_2 _41048_ (.CLK(clk),
    .D(_03542_),
    .Q(mem_wdata[6]));
 sky130_fd_sc_hd__dfxtp_2 _41049_ (.CLK(clk),
    .D(_03543_),
    .Q(mem_wdata[7]));
 sky130_fd_sc_hd__dfxtp_2 _41050_ (.CLK(clk),
    .D(_03544_),
    .Q(mem_wdata[8]));
 sky130_fd_sc_hd__dfxtp_2 _41051_ (.CLK(clk),
    .D(_03545_),
    .Q(mem_wdata[9]));
 sky130_fd_sc_hd__dfxtp_2 _41052_ (.CLK(clk),
    .D(_03546_),
    .Q(mem_wdata[10]));
 sky130_fd_sc_hd__dfxtp_2 _41053_ (.CLK(clk),
    .D(_03547_),
    .Q(mem_wdata[11]));
 sky130_fd_sc_hd__dfxtp_2 _41054_ (.CLK(clk),
    .D(_03548_),
    .Q(mem_wdata[12]));
 sky130_fd_sc_hd__dfxtp_2 _41055_ (.CLK(clk),
    .D(_03549_),
    .Q(mem_wdata[13]));
 sky130_fd_sc_hd__dfxtp_2 _41056_ (.CLK(clk),
    .D(_03550_),
    .Q(mem_wdata[14]));
 sky130_fd_sc_hd__dfxtp_2 _41057_ (.CLK(clk),
    .D(_03551_),
    .Q(mem_wdata[15]));
 sky130_fd_sc_hd__dfxtp_2 _41058_ (.CLK(clk),
    .D(_03552_),
    .Q(mem_wdata[16]));
 sky130_fd_sc_hd__dfxtp_2 _41059_ (.CLK(clk),
    .D(_03553_),
    .Q(mem_wdata[17]));
 sky130_fd_sc_hd__dfxtp_2 _41060_ (.CLK(clk),
    .D(_03554_),
    .Q(mem_wdata[18]));
 sky130_fd_sc_hd__dfxtp_2 _41061_ (.CLK(clk),
    .D(_03555_),
    .Q(mem_wdata[19]));
 sky130_fd_sc_hd__dfxtp_2 _41062_ (.CLK(clk),
    .D(_03556_),
    .Q(mem_wdata[20]));
 sky130_fd_sc_hd__dfxtp_2 _41063_ (.CLK(clk),
    .D(_03557_),
    .Q(mem_wdata[21]));
 sky130_fd_sc_hd__dfxtp_2 _41064_ (.CLK(clk),
    .D(_03558_),
    .Q(mem_wdata[22]));
 sky130_fd_sc_hd__dfxtp_2 _41065_ (.CLK(clk),
    .D(_03559_),
    .Q(mem_wdata[23]));
 sky130_fd_sc_hd__dfxtp_2 _41066_ (.CLK(clk),
    .D(_03560_),
    .Q(mem_wdata[24]));
 sky130_fd_sc_hd__dfxtp_2 _41067_ (.CLK(clk),
    .D(_03561_),
    .Q(mem_wdata[25]));
 sky130_fd_sc_hd__dfxtp_2 _41068_ (.CLK(clk),
    .D(_03562_),
    .Q(mem_wdata[26]));
 sky130_fd_sc_hd__dfxtp_2 _41069_ (.CLK(clk),
    .D(_03563_),
    .Q(mem_wdata[27]));
 sky130_fd_sc_hd__dfxtp_2 _41070_ (.CLK(clk),
    .D(_03564_),
    .Q(mem_wdata[28]));
 sky130_fd_sc_hd__dfxtp_2 _41071_ (.CLK(clk),
    .D(_03565_),
    .Q(mem_wdata[29]));
 sky130_fd_sc_hd__dfxtp_2 _41072_ (.CLK(clk),
    .D(_03566_),
    .Q(mem_wdata[30]));
 sky130_fd_sc_hd__dfxtp_2 _41073_ (.CLK(clk),
    .D(_03567_),
    .Q(mem_wdata[31]));
 sky130_fd_sc_hd__dfxtp_2 _41074_ (.CLK(clk),
    .D(_03568_),
    .Q(\cpuregs[19][0] ));
 sky130_fd_sc_hd__dfxtp_2 _41075_ (.CLK(clk),
    .D(_03569_),
    .Q(\cpuregs[19][1] ));
 sky130_fd_sc_hd__dfxtp_2 _41076_ (.CLK(clk),
    .D(_03570_),
    .Q(\cpuregs[19][2] ));
 sky130_fd_sc_hd__dfxtp_2 _41077_ (.CLK(clk),
    .D(_03571_),
    .Q(\cpuregs[19][3] ));
 sky130_fd_sc_hd__dfxtp_2 _41078_ (.CLK(clk),
    .D(_03572_),
    .Q(\cpuregs[19][4] ));
 sky130_fd_sc_hd__dfxtp_2 _41079_ (.CLK(clk),
    .D(_03573_),
    .Q(\cpuregs[19][5] ));
 sky130_fd_sc_hd__dfxtp_2 _41080_ (.CLK(clk),
    .D(_03574_),
    .Q(\cpuregs[19][6] ));
 sky130_fd_sc_hd__dfxtp_2 _41081_ (.CLK(clk),
    .D(_03575_),
    .Q(\cpuregs[19][7] ));
 sky130_fd_sc_hd__dfxtp_2 _41082_ (.CLK(clk),
    .D(_03576_),
    .Q(\cpuregs[19][8] ));
 sky130_fd_sc_hd__dfxtp_2 _41083_ (.CLK(clk),
    .D(_03577_),
    .Q(\cpuregs[19][9] ));
 sky130_fd_sc_hd__dfxtp_2 _41084_ (.CLK(clk),
    .D(_03578_),
    .Q(\cpuregs[19][10] ));
 sky130_fd_sc_hd__dfxtp_2 _41085_ (.CLK(clk),
    .D(_03579_),
    .Q(\cpuregs[19][11] ));
 sky130_fd_sc_hd__dfxtp_2 _41086_ (.CLK(clk),
    .D(_03580_),
    .Q(\cpuregs[19][12] ));
 sky130_fd_sc_hd__dfxtp_2 _41087_ (.CLK(clk),
    .D(_03581_),
    .Q(\cpuregs[19][13] ));
 sky130_fd_sc_hd__dfxtp_2 _41088_ (.CLK(clk),
    .D(_03582_),
    .Q(\cpuregs[19][14] ));
 sky130_fd_sc_hd__dfxtp_2 _41089_ (.CLK(clk),
    .D(_03583_),
    .Q(\cpuregs[19][15] ));
 sky130_fd_sc_hd__dfxtp_2 _41090_ (.CLK(clk),
    .D(_03584_),
    .Q(\cpuregs[19][16] ));
 sky130_fd_sc_hd__dfxtp_2 _41091_ (.CLK(clk),
    .D(_03585_),
    .Q(\cpuregs[19][17] ));
 sky130_fd_sc_hd__dfxtp_2 _41092_ (.CLK(clk),
    .D(_03586_),
    .Q(\cpuregs[19][18] ));
 sky130_fd_sc_hd__dfxtp_2 _41093_ (.CLK(clk),
    .D(_03587_),
    .Q(\cpuregs[19][19] ));
 sky130_fd_sc_hd__dfxtp_2 _41094_ (.CLK(clk),
    .D(_03588_),
    .Q(\cpuregs[19][20] ));
 sky130_fd_sc_hd__dfxtp_2 _41095_ (.CLK(clk),
    .D(_03589_),
    .Q(\cpuregs[19][21] ));
 sky130_fd_sc_hd__dfxtp_2 _41096_ (.CLK(clk),
    .D(_03590_),
    .Q(\cpuregs[19][22] ));
 sky130_fd_sc_hd__dfxtp_2 _41097_ (.CLK(clk),
    .D(_03591_),
    .Q(\cpuregs[19][23] ));
 sky130_fd_sc_hd__dfxtp_2 _41098_ (.CLK(clk),
    .D(_03592_),
    .Q(\cpuregs[19][24] ));
 sky130_fd_sc_hd__dfxtp_2 _41099_ (.CLK(clk),
    .D(_03593_),
    .Q(\cpuregs[19][25] ));
 sky130_fd_sc_hd__dfxtp_2 _41100_ (.CLK(clk),
    .D(_03594_),
    .Q(\cpuregs[19][26] ));
 sky130_fd_sc_hd__dfxtp_2 _41101_ (.CLK(clk),
    .D(_03595_),
    .Q(\cpuregs[19][27] ));
 sky130_fd_sc_hd__dfxtp_2 _41102_ (.CLK(clk),
    .D(_03596_),
    .Q(\cpuregs[19][28] ));
 sky130_fd_sc_hd__dfxtp_2 _41103_ (.CLK(clk),
    .D(_03597_),
    .Q(\cpuregs[19][29] ));
 sky130_fd_sc_hd__dfxtp_2 _41104_ (.CLK(clk),
    .D(_03598_),
    .Q(\cpuregs[19][30] ));
 sky130_fd_sc_hd__dfxtp_2 _41105_ (.CLK(clk),
    .D(_03599_),
    .Q(\cpuregs[19][31] ));
 sky130_fd_sc_hd__dfxtp_2 _41106_ (.CLK(clk),
    .D(_03600_),
    .Q(\cpuregs[4][0] ));
 sky130_fd_sc_hd__dfxtp_2 _41107_ (.CLK(clk),
    .D(_03601_),
    .Q(\cpuregs[4][1] ));
 sky130_fd_sc_hd__dfxtp_2 _41108_ (.CLK(clk),
    .D(_03602_),
    .Q(\cpuregs[4][2] ));
 sky130_fd_sc_hd__dfxtp_2 _41109_ (.CLK(clk),
    .D(_03603_),
    .Q(\cpuregs[4][3] ));
 sky130_fd_sc_hd__dfxtp_2 _41110_ (.CLK(clk),
    .D(_03604_),
    .Q(\cpuregs[4][4] ));
 sky130_fd_sc_hd__dfxtp_2 _41111_ (.CLK(clk),
    .D(_03605_),
    .Q(\cpuregs[4][5] ));
 sky130_fd_sc_hd__dfxtp_2 _41112_ (.CLK(clk),
    .D(_03606_),
    .Q(\cpuregs[4][6] ));
 sky130_fd_sc_hd__dfxtp_2 _41113_ (.CLK(clk),
    .D(_03607_),
    .Q(\cpuregs[4][7] ));
 sky130_fd_sc_hd__dfxtp_2 _41114_ (.CLK(clk),
    .D(_03608_),
    .Q(\cpuregs[4][8] ));
 sky130_fd_sc_hd__dfxtp_2 _41115_ (.CLK(clk),
    .D(_03609_),
    .Q(\cpuregs[4][9] ));
 sky130_fd_sc_hd__dfxtp_2 _41116_ (.CLK(clk),
    .D(_03610_),
    .Q(\cpuregs[4][10] ));
 sky130_fd_sc_hd__dfxtp_2 _41117_ (.CLK(clk),
    .D(_03611_),
    .Q(\cpuregs[4][11] ));
 sky130_fd_sc_hd__dfxtp_2 _41118_ (.CLK(clk),
    .D(_03612_),
    .Q(\cpuregs[4][12] ));
 sky130_fd_sc_hd__dfxtp_2 _41119_ (.CLK(clk),
    .D(_03613_),
    .Q(\cpuregs[4][13] ));
 sky130_fd_sc_hd__dfxtp_2 _41120_ (.CLK(clk),
    .D(_03614_),
    .Q(\cpuregs[4][14] ));
 sky130_fd_sc_hd__dfxtp_2 _41121_ (.CLK(clk),
    .D(_03615_),
    .Q(\cpuregs[4][15] ));
 sky130_fd_sc_hd__dfxtp_2 _41122_ (.CLK(clk),
    .D(_03616_),
    .Q(\cpuregs[4][16] ));
 sky130_fd_sc_hd__dfxtp_2 _41123_ (.CLK(clk),
    .D(_03617_),
    .Q(\cpuregs[4][17] ));
 sky130_fd_sc_hd__dfxtp_2 _41124_ (.CLK(clk),
    .D(_03618_),
    .Q(\cpuregs[4][18] ));
 sky130_fd_sc_hd__dfxtp_2 _41125_ (.CLK(clk),
    .D(_03619_),
    .Q(\cpuregs[4][19] ));
 sky130_fd_sc_hd__dfxtp_2 _41126_ (.CLK(clk),
    .D(_03620_),
    .Q(\cpuregs[4][20] ));
 sky130_fd_sc_hd__dfxtp_2 _41127_ (.CLK(clk),
    .D(_03621_),
    .Q(\cpuregs[4][21] ));
 sky130_fd_sc_hd__dfxtp_2 _41128_ (.CLK(clk),
    .D(_03622_),
    .Q(\cpuregs[4][22] ));
 sky130_fd_sc_hd__dfxtp_2 _41129_ (.CLK(clk),
    .D(_03623_),
    .Q(\cpuregs[4][23] ));
 sky130_fd_sc_hd__dfxtp_2 _41130_ (.CLK(clk),
    .D(_03624_),
    .Q(\cpuregs[4][24] ));
 sky130_fd_sc_hd__dfxtp_2 _41131_ (.CLK(clk),
    .D(_03625_),
    .Q(\cpuregs[4][25] ));
 sky130_fd_sc_hd__dfxtp_2 _41132_ (.CLK(clk),
    .D(_03626_),
    .Q(\cpuregs[4][26] ));
 sky130_fd_sc_hd__dfxtp_2 _41133_ (.CLK(clk),
    .D(_03627_),
    .Q(\cpuregs[4][27] ));
 sky130_fd_sc_hd__dfxtp_2 _41134_ (.CLK(clk),
    .D(_03628_),
    .Q(\cpuregs[4][28] ));
 sky130_fd_sc_hd__dfxtp_2 _41135_ (.CLK(clk),
    .D(_03629_),
    .Q(\cpuregs[4][29] ));
 sky130_fd_sc_hd__dfxtp_2 _41136_ (.CLK(clk),
    .D(_03630_),
    .Q(\cpuregs[4][30] ));
 sky130_fd_sc_hd__dfxtp_2 _41137_ (.CLK(clk),
    .D(_03631_),
    .Q(\cpuregs[4][31] ));
 sky130_fd_sc_hd__dfxtp_2 _41138_ (.CLK(clk),
    .D(_03632_),
    .Q(mem_la_wdata[0]));
 sky130_fd_sc_hd__dfxtp_2 _41139_ (.CLK(clk),
    .D(_03633_),
    .Q(mem_la_wdata[1]));
 sky130_fd_sc_hd__dfxtp_2 _41140_ (.CLK(clk),
    .D(_03634_),
    .Q(mem_la_wdata[2]));
 sky130_fd_sc_hd__dfxtp_2 _41141_ (.CLK(clk),
    .D(_03635_),
    .Q(mem_la_wdata[3]));
 sky130_fd_sc_hd__dfxtp_2 _41142_ (.CLK(clk),
    .D(_03636_),
    .Q(mem_la_wdata[4]));
 sky130_fd_sc_hd__dfxtp_2 _41143_ (.CLK(clk),
    .D(_03637_),
    .Q(mem_la_wdata[5]));
 sky130_fd_sc_hd__dfxtp_2 _41144_ (.CLK(clk),
    .D(_03638_),
    .Q(mem_la_wdata[6]));
 sky130_fd_sc_hd__dfxtp_2 _41145_ (.CLK(clk),
    .D(_03639_),
    .Q(mem_la_wdata[7]));
 sky130_fd_sc_hd__dfxtp_2 _41146_ (.CLK(clk),
    .D(_03640_),
    .Q(pcpi_rs2[8]));
 sky130_fd_sc_hd__dfxtp_2 _41147_ (.CLK(clk),
    .D(_03641_),
    .Q(pcpi_rs2[9]));
 sky130_fd_sc_hd__dfxtp_2 _41148_ (.CLK(clk),
    .D(_03642_),
    .Q(pcpi_rs2[10]));
 sky130_fd_sc_hd__dfxtp_2 _41149_ (.CLK(clk),
    .D(_03643_),
    .Q(pcpi_rs2[11]));
 sky130_fd_sc_hd__dfxtp_2 _41150_ (.CLK(clk),
    .D(_03644_),
    .Q(pcpi_rs2[12]));
 sky130_fd_sc_hd__dfxtp_2 _41151_ (.CLK(clk),
    .D(_03645_),
    .Q(pcpi_rs2[13]));
 sky130_fd_sc_hd__dfxtp_2 _41152_ (.CLK(clk),
    .D(_03646_),
    .Q(pcpi_rs2[14]));
 sky130_fd_sc_hd__dfxtp_2 _41153_ (.CLK(clk),
    .D(_03647_),
    .Q(pcpi_rs2[15]));
 sky130_fd_sc_hd__dfxtp_2 _41154_ (.CLK(clk),
    .D(_03648_),
    .Q(pcpi_rs2[16]));
 sky130_fd_sc_hd__dfxtp_2 _41155_ (.CLK(clk),
    .D(_03649_),
    .Q(pcpi_rs2[17]));
 sky130_fd_sc_hd__dfxtp_2 _41156_ (.CLK(clk),
    .D(_03650_),
    .Q(pcpi_rs2[18]));
 sky130_fd_sc_hd__dfxtp_2 _41157_ (.CLK(clk),
    .D(_03651_),
    .Q(pcpi_rs2[19]));
 sky130_fd_sc_hd__dfxtp_2 _41158_ (.CLK(clk),
    .D(_03652_),
    .Q(pcpi_rs2[20]));
 sky130_fd_sc_hd__dfxtp_2 _41159_ (.CLK(clk),
    .D(_03653_),
    .Q(pcpi_rs2[21]));
 sky130_fd_sc_hd__dfxtp_2 _41160_ (.CLK(clk),
    .D(_03654_),
    .Q(pcpi_rs2[22]));
 sky130_fd_sc_hd__dfxtp_2 _41161_ (.CLK(clk),
    .D(_03655_),
    .Q(pcpi_rs2[23]));
 sky130_fd_sc_hd__dfxtp_2 _41162_ (.CLK(clk),
    .D(_03656_),
    .Q(pcpi_rs2[24]));
 sky130_fd_sc_hd__dfxtp_2 _41163_ (.CLK(clk),
    .D(_03657_),
    .Q(pcpi_rs2[25]));
 sky130_fd_sc_hd__dfxtp_2 _41164_ (.CLK(clk),
    .D(_03658_),
    .Q(pcpi_rs2[26]));
 sky130_fd_sc_hd__dfxtp_2 _41165_ (.CLK(clk),
    .D(_03659_),
    .Q(pcpi_rs2[27]));
 sky130_fd_sc_hd__dfxtp_2 _41166_ (.CLK(clk),
    .D(_03660_),
    .Q(pcpi_rs2[28]));
 sky130_fd_sc_hd__dfxtp_2 _41167_ (.CLK(clk),
    .D(_03661_),
    .Q(pcpi_rs2[29]));
 sky130_fd_sc_hd__dfxtp_2 _41168_ (.CLK(clk),
    .D(_03662_),
    .Q(pcpi_rs2[30]));
 sky130_fd_sc_hd__dfxtp_2 _41169_ (.CLK(clk),
    .D(_03663_),
    .Q(pcpi_rs2[31]));
 sky130_fd_sc_hd__dfxtp_2 _41170_ (.CLK(clk),
    .D(_03664_),
    .Q(\cpuregs[9][0] ));
 sky130_fd_sc_hd__dfxtp_2 _41171_ (.CLK(clk),
    .D(_03665_),
    .Q(\cpuregs[9][1] ));
 sky130_fd_sc_hd__dfxtp_2 _41172_ (.CLK(clk),
    .D(_03666_),
    .Q(\cpuregs[9][2] ));
 sky130_fd_sc_hd__dfxtp_2 _41173_ (.CLK(clk),
    .D(_03667_),
    .Q(\cpuregs[9][3] ));
 sky130_fd_sc_hd__dfxtp_2 _41174_ (.CLK(clk),
    .D(_03668_),
    .Q(\cpuregs[9][4] ));
 sky130_fd_sc_hd__dfxtp_2 _41175_ (.CLK(clk),
    .D(_03669_),
    .Q(\cpuregs[9][5] ));
 sky130_fd_sc_hd__dfxtp_2 _41176_ (.CLK(clk),
    .D(_03670_),
    .Q(\cpuregs[9][6] ));
 sky130_fd_sc_hd__dfxtp_2 _41177_ (.CLK(clk),
    .D(_03671_),
    .Q(\cpuregs[9][7] ));
 sky130_fd_sc_hd__dfxtp_2 _41178_ (.CLK(clk),
    .D(_03672_),
    .Q(\cpuregs[9][8] ));
 sky130_fd_sc_hd__dfxtp_2 _41179_ (.CLK(clk),
    .D(_03673_),
    .Q(\cpuregs[9][9] ));
 sky130_fd_sc_hd__dfxtp_2 _41180_ (.CLK(clk),
    .D(_03674_),
    .Q(\cpuregs[9][10] ));
 sky130_fd_sc_hd__dfxtp_2 _41181_ (.CLK(clk),
    .D(_03675_),
    .Q(\cpuregs[9][11] ));
 sky130_fd_sc_hd__dfxtp_2 _41182_ (.CLK(clk),
    .D(_03676_),
    .Q(\cpuregs[9][12] ));
 sky130_fd_sc_hd__dfxtp_2 _41183_ (.CLK(clk),
    .D(_03677_),
    .Q(\cpuregs[9][13] ));
 sky130_fd_sc_hd__dfxtp_2 _41184_ (.CLK(clk),
    .D(_03678_),
    .Q(\cpuregs[9][14] ));
 sky130_fd_sc_hd__dfxtp_2 _41185_ (.CLK(clk),
    .D(_03679_),
    .Q(\cpuregs[9][15] ));
 sky130_fd_sc_hd__dfxtp_2 _41186_ (.CLK(clk),
    .D(_03680_),
    .Q(\cpuregs[9][16] ));
 sky130_fd_sc_hd__dfxtp_2 _41187_ (.CLK(clk),
    .D(_03681_),
    .Q(\cpuregs[9][17] ));
 sky130_fd_sc_hd__dfxtp_2 _41188_ (.CLK(clk),
    .D(_03682_),
    .Q(\cpuregs[9][18] ));
 sky130_fd_sc_hd__dfxtp_2 _41189_ (.CLK(clk),
    .D(_03683_),
    .Q(\cpuregs[9][19] ));
 sky130_fd_sc_hd__dfxtp_2 _41190_ (.CLK(clk),
    .D(_03684_),
    .Q(\cpuregs[9][20] ));
 sky130_fd_sc_hd__dfxtp_2 _41191_ (.CLK(clk),
    .D(_03685_),
    .Q(\cpuregs[9][21] ));
 sky130_fd_sc_hd__dfxtp_2 _41192_ (.CLK(clk),
    .D(_03686_),
    .Q(\cpuregs[9][22] ));
 sky130_fd_sc_hd__dfxtp_2 _41193_ (.CLK(clk),
    .D(_03687_),
    .Q(\cpuregs[9][23] ));
 sky130_fd_sc_hd__dfxtp_2 _41194_ (.CLK(clk),
    .D(_03688_),
    .Q(\cpuregs[9][24] ));
 sky130_fd_sc_hd__dfxtp_2 _41195_ (.CLK(clk),
    .D(_03689_),
    .Q(\cpuregs[9][25] ));
 sky130_fd_sc_hd__dfxtp_2 _41196_ (.CLK(clk),
    .D(_03690_),
    .Q(\cpuregs[9][26] ));
 sky130_fd_sc_hd__dfxtp_2 _41197_ (.CLK(clk),
    .D(_03691_),
    .Q(\cpuregs[9][27] ));
 sky130_fd_sc_hd__dfxtp_2 _41198_ (.CLK(clk),
    .D(_03692_),
    .Q(\cpuregs[9][28] ));
 sky130_fd_sc_hd__dfxtp_2 _41199_ (.CLK(clk),
    .D(_03693_),
    .Q(\cpuregs[9][29] ));
 sky130_fd_sc_hd__dfxtp_2 _41200_ (.CLK(clk),
    .D(_03694_),
    .Q(\cpuregs[9][30] ));
 sky130_fd_sc_hd__dfxtp_2 _41201_ (.CLK(clk),
    .D(_03695_),
    .Q(\cpuregs[9][31] ));
 sky130_fd_sc_hd__dfxtp_2 _41202_ (.CLK(clk),
    .D(_03696_),
    .Q(\cpuregs[6][0] ));
 sky130_fd_sc_hd__dfxtp_2 _41203_ (.CLK(clk),
    .D(_03697_),
    .Q(\cpuregs[6][1] ));
 sky130_fd_sc_hd__dfxtp_2 _41204_ (.CLK(clk),
    .D(_03698_),
    .Q(\cpuregs[6][2] ));
 sky130_fd_sc_hd__dfxtp_2 _41205_ (.CLK(clk),
    .D(_03699_),
    .Q(\cpuregs[6][3] ));
 sky130_fd_sc_hd__dfxtp_2 _41206_ (.CLK(clk),
    .D(_03700_),
    .Q(\cpuregs[6][4] ));
 sky130_fd_sc_hd__dfxtp_2 _41207_ (.CLK(clk),
    .D(_03701_),
    .Q(\cpuregs[6][5] ));
 sky130_fd_sc_hd__dfxtp_2 _41208_ (.CLK(clk),
    .D(_03702_),
    .Q(\cpuregs[6][6] ));
 sky130_fd_sc_hd__dfxtp_2 _41209_ (.CLK(clk),
    .D(_03703_),
    .Q(\cpuregs[6][7] ));
 sky130_fd_sc_hd__dfxtp_2 _41210_ (.CLK(clk),
    .D(_03704_),
    .Q(\cpuregs[6][8] ));
 sky130_fd_sc_hd__dfxtp_2 _41211_ (.CLK(clk),
    .D(_03705_),
    .Q(\cpuregs[6][9] ));
 sky130_fd_sc_hd__dfxtp_2 _41212_ (.CLK(clk),
    .D(_03706_),
    .Q(\cpuregs[6][10] ));
 sky130_fd_sc_hd__dfxtp_2 _41213_ (.CLK(clk),
    .D(_03707_),
    .Q(\cpuregs[6][11] ));
 sky130_fd_sc_hd__dfxtp_2 _41214_ (.CLK(clk),
    .D(_03708_),
    .Q(\cpuregs[6][12] ));
 sky130_fd_sc_hd__dfxtp_2 _41215_ (.CLK(clk),
    .D(_03709_),
    .Q(\cpuregs[6][13] ));
 sky130_fd_sc_hd__dfxtp_2 _41216_ (.CLK(clk),
    .D(_03710_),
    .Q(\cpuregs[6][14] ));
 sky130_fd_sc_hd__dfxtp_2 _41217_ (.CLK(clk),
    .D(_03711_),
    .Q(\cpuregs[6][15] ));
 sky130_fd_sc_hd__dfxtp_2 _41218_ (.CLK(clk),
    .D(_03712_),
    .Q(\cpuregs[6][16] ));
 sky130_fd_sc_hd__dfxtp_2 _41219_ (.CLK(clk),
    .D(_03713_),
    .Q(\cpuregs[6][17] ));
 sky130_fd_sc_hd__dfxtp_2 _41220_ (.CLK(clk),
    .D(_03714_),
    .Q(\cpuregs[6][18] ));
 sky130_fd_sc_hd__dfxtp_2 _41221_ (.CLK(clk),
    .D(_03715_),
    .Q(\cpuregs[6][19] ));
 sky130_fd_sc_hd__dfxtp_2 _41222_ (.CLK(clk),
    .D(_03716_),
    .Q(\cpuregs[6][20] ));
 sky130_fd_sc_hd__dfxtp_2 _41223_ (.CLK(clk),
    .D(_03717_),
    .Q(\cpuregs[6][21] ));
 sky130_fd_sc_hd__dfxtp_2 _41224_ (.CLK(clk),
    .D(_03718_),
    .Q(\cpuregs[6][22] ));
 sky130_fd_sc_hd__dfxtp_2 _41225_ (.CLK(clk),
    .D(_03719_),
    .Q(\cpuregs[6][23] ));
 sky130_fd_sc_hd__dfxtp_2 _41226_ (.CLK(clk),
    .D(_03720_),
    .Q(\cpuregs[6][24] ));
 sky130_fd_sc_hd__dfxtp_2 _41227_ (.CLK(clk),
    .D(_03721_),
    .Q(\cpuregs[6][25] ));
 sky130_fd_sc_hd__dfxtp_2 _41228_ (.CLK(clk),
    .D(_03722_),
    .Q(\cpuregs[6][26] ));
 sky130_fd_sc_hd__dfxtp_2 _41229_ (.CLK(clk),
    .D(_03723_),
    .Q(\cpuregs[6][27] ));
 sky130_fd_sc_hd__dfxtp_2 _41230_ (.CLK(clk),
    .D(_03724_),
    .Q(\cpuregs[6][28] ));
 sky130_fd_sc_hd__dfxtp_2 _41231_ (.CLK(clk),
    .D(_03725_),
    .Q(\cpuregs[6][29] ));
 sky130_fd_sc_hd__dfxtp_2 _41232_ (.CLK(clk),
    .D(_03726_),
    .Q(\cpuregs[6][30] ));
 sky130_fd_sc_hd__dfxtp_2 _41233_ (.CLK(clk),
    .D(_03727_),
    .Q(\cpuregs[6][31] ));
 sky130_fd_sc_hd__dfxtp_2 _41234_ (.CLK(clk),
    .D(_03728_),
    .Q(\pcpi_mul.active[0] ));
 sky130_fd_sc_hd__dfxtp_2 _41235_ (.CLK(clk),
    .D(_03729_),
    .Q(\pcpi_mul.active[1] ));
 sky130_fd_sc_hd__dfxtp_2 _41236_ (.CLK(clk),
    .D(_03730_),
    .Q(trap));
 sky130_fd_sc_hd__dfxtp_2 _41237_ (.CLK(clk),
    .D(_03731_),
    .Q(\count_cycle[0] ));
 sky130_fd_sc_hd__dfxtp_2 _41238_ (.CLK(clk),
    .D(_03732_),
    .Q(\count_cycle[1] ));
 sky130_fd_sc_hd__dfxtp_2 _41239_ (.CLK(clk),
    .D(_03733_),
    .Q(\count_cycle[2] ));
 sky130_fd_sc_hd__dfxtp_2 _41240_ (.CLK(clk),
    .D(_03734_),
    .Q(\count_cycle[3] ));
 sky130_fd_sc_hd__dfxtp_2 _41241_ (.CLK(clk),
    .D(_03735_),
    .Q(\count_cycle[4] ));
 sky130_fd_sc_hd__dfxtp_2 _41242_ (.CLK(clk),
    .D(_03736_),
    .Q(\count_cycle[5] ));
 sky130_fd_sc_hd__dfxtp_2 _41243_ (.CLK(clk),
    .D(_03737_),
    .Q(\count_cycle[6] ));
 sky130_fd_sc_hd__dfxtp_2 _41244_ (.CLK(clk),
    .D(_03738_),
    .Q(\count_cycle[7] ));
 sky130_fd_sc_hd__dfxtp_2 _41245_ (.CLK(clk),
    .D(_03739_),
    .Q(\count_cycle[8] ));
 sky130_fd_sc_hd__dfxtp_2 _41246_ (.CLK(clk),
    .D(_03740_),
    .Q(\count_cycle[9] ));
 sky130_fd_sc_hd__dfxtp_2 _41247_ (.CLK(clk),
    .D(_03741_),
    .Q(\count_cycle[10] ));
 sky130_fd_sc_hd__dfxtp_2 _41248_ (.CLK(clk),
    .D(_03742_),
    .Q(\count_cycle[11] ));
 sky130_fd_sc_hd__dfxtp_2 _41249_ (.CLK(clk),
    .D(_03743_),
    .Q(\count_cycle[12] ));
 sky130_fd_sc_hd__dfxtp_2 _41250_ (.CLK(clk),
    .D(_03744_),
    .Q(\count_cycle[13] ));
 sky130_fd_sc_hd__dfxtp_2 _41251_ (.CLK(clk),
    .D(_03745_),
    .Q(\count_cycle[14] ));
 sky130_fd_sc_hd__dfxtp_2 _41252_ (.CLK(clk),
    .D(_03746_),
    .Q(\count_cycle[15] ));
 sky130_fd_sc_hd__dfxtp_2 _41253_ (.CLK(clk),
    .D(_03747_),
    .Q(\count_cycle[16] ));
 sky130_fd_sc_hd__dfxtp_2 _41254_ (.CLK(clk),
    .D(_03748_),
    .Q(\count_cycle[17] ));
 sky130_fd_sc_hd__dfxtp_2 _41255_ (.CLK(clk),
    .D(_03749_),
    .Q(\count_cycle[18] ));
 sky130_fd_sc_hd__dfxtp_2 _41256_ (.CLK(clk),
    .D(_03750_),
    .Q(\count_cycle[19] ));
 sky130_fd_sc_hd__dfxtp_2 _41257_ (.CLK(clk),
    .D(_03751_),
    .Q(\count_cycle[20] ));
 sky130_fd_sc_hd__dfxtp_2 _41258_ (.CLK(clk),
    .D(_03752_),
    .Q(\count_cycle[21] ));
 sky130_fd_sc_hd__dfxtp_2 _41259_ (.CLK(clk),
    .D(_03753_),
    .Q(\count_cycle[22] ));
 sky130_fd_sc_hd__dfxtp_2 _41260_ (.CLK(clk),
    .D(_03754_),
    .Q(\count_cycle[23] ));
 sky130_fd_sc_hd__dfxtp_2 _41261_ (.CLK(clk),
    .D(_03755_),
    .Q(\count_cycle[24] ));
 sky130_fd_sc_hd__dfxtp_2 _41262_ (.CLK(clk),
    .D(_03756_),
    .Q(\count_cycle[25] ));
 sky130_fd_sc_hd__dfxtp_2 _41263_ (.CLK(clk),
    .D(_03757_),
    .Q(\count_cycle[26] ));
 sky130_fd_sc_hd__dfxtp_2 _41264_ (.CLK(clk),
    .D(_03758_),
    .Q(\count_cycle[27] ));
 sky130_fd_sc_hd__dfxtp_2 _41265_ (.CLK(clk),
    .D(_03759_),
    .Q(\count_cycle[28] ));
 sky130_fd_sc_hd__dfxtp_2 _41266_ (.CLK(clk),
    .D(_03760_),
    .Q(\count_cycle[29] ));
 sky130_fd_sc_hd__dfxtp_2 _41267_ (.CLK(clk),
    .D(_03761_),
    .Q(\count_cycle[30] ));
 sky130_fd_sc_hd__dfxtp_2 _41268_ (.CLK(clk),
    .D(_03762_),
    .Q(\count_cycle[31] ));
 sky130_fd_sc_hd__dfxtp_2 _41269_ (.CLK(clk),
    .D(_03763_),
    .Q(\count_cycle[32] ));
 sky130_fd_sc_hd__dfxtp_2 _41270_ (.CLK(clk),
    .D(_03764_),
    .Q(\count_cycle[33] ));
 sky130_fd_sc_hd__dfxtp_2 _41271_ (.CLK(clk),
    .D(_03765_),
    .Q(\count_cycle[34] ));
 sky130_fd_sc_hd__dfxtp_2 _41272_ (.CLK(clk),
    .D(_03766_),
    .Q(\count_cycle[35] ));
 sky130_fd_sc_hd__dfxtp_2 _41273_ (.CLK(clk),
    .D(_03767_),
    .Q(\count_cycle[36] ));
 sky130_fd_sc_hd__dfxtp_2 _41274_ (.CLK(clk),
    .D(_03768_),
    .Q(\count_cycle[37] ));
 sky130_fd_sc_hd__dfxtp_2 _41275_ (.CLK(clk),
    .D(_03769_),
    .Q(\count_cycle[38] ));
 sky130_fd_sc_hd__dfxtp_2 _41276_ (.CLK(clk),
    .D(_03770_),
    .Q(\count_cycle[39] ));
 sky130_fd_sc_hd__dfxtp_2 _41277_ (.CLK(clk),
    .D(_03771_),
    .Q(\count_cycle[40] ));
 sky130_fd_sc_hd__dfxtp_2 _41278_ (.CLK(clk),
    .D(_03772_),
    .Q(\count_cycle[41] ));
 sky130_fd_sc_hd__dfxtp_2 _41279_ (.CLK(clk),
    .D(_03773_),
    .Q(\count_cycle[42] ));
 sky130_fd_sc_hd__dfxtp_2 _41280_ (.CLK(clk),
    .D(_03774_),
    .Q(\count_cycle[43] ));
 sky130_fd_sc_hd__dfxtp_2 _41281_ (.CLK(clk),
    .D(_03775_),
    .Q(\count_cycle[44] ));
 sky130_fd_sc_hd__dfxtp_2 _41282_ (.CLK(clk),
    .D(_03776_),
    .Q(\count_cycle[45] ));
 sky130_fd_sc_hd__dfxtp_2 _41283_ (.CLK(clk),
    .D(_03777_),
    .Q(\count_cycle[46] ));
 sky130_fd_sc_hd__dfxtp_2 _41284_ (.CLK(clk),
    .D(_03778_),
    .Q(\count_cycle[47] ));
 sky130_fd_sc_hd__dfxtp_2 _41285_ (.CLK(clk),
    .D(_03779_),
    .Q(\count_cycle[48] ));
 sky130_fd_sc_hd__dfxtp_2 _41286_ (.CLK(clk),
    .D(_03780_),
    .Q(\count_cycle[49] ));
 sky130_fd_sc_hd__dfxtp_2 _41287_ (.CLK(clk),
    .D(_03781_),
    .Q(\count_cycle[50] ));
 sky130_fd_sc_hd__dfxtp_2 _41288_ (.CLK(clk),
    .D(_03782_),
    .Q(\count_cycle[51] ));
 sky130_fd_sc_hd__dfxtp_2 _41289_ (.CLK(clk),
    .D(_03783_),
    .Q(\count_cycle[52] ));
 sky130_fd_sc_hd__dfxtp_2 _41290_ (.CLK(clk),
    .D(_03784_),
    .Q(\count_cycle[53] ));
 sky130_fd_sc_hd__dfxtp_2 _41291_ (.CLK(clk),
    .D(_03785_),
    .Q(\count_cycle[54] ));
 sky130_fd_sc_hd__dfxtp_2 _41292_ (.CLK(clk),
    .D(_03786_),
    .Q(\count_cycle[55] ));
 sky130_fd_sc_hd__dfxtp_2 _41293_ (.CLK(clk),
    .D(_03787_),
    .Q(\count_cycle[56] ));
 sky130_fd_sc_hd__dfxtp_2 _41294_ (.CLK(clk),
    .D(_03788_),
    .Q(\count_cycle[57] ));
 sky130_fd_sc_hd__dfxtp_2 _41295_ (.CLK(clk),
    .D(_03789_),
    .Q(\count_cycle[58] ));
 sky130_fd_sc_hd__dfxtp_2 _41296_ (.CLK(clk),
    .D(_03790_),
    .Q(\count_cycle[59] ));
 sky130_fd_sc_hd__dfxtp_2 _41297_ (.CLK(clk),
    .D(_03791_),
    .Q(\count_cycle[60] ));
 sky130_fd_sc_hd__dfxtp_2 _41298_ (.CLK(clk),
    .D(_03792_),
    .Q(\count_cycle[61] ));
 sky130_fd_sc_hd__dfxtp_2 _41299_ (.CLK(clk),
    .D(_03793_),
    .Q(\count_cycle[62] ));
 sky130_fd_sc_hd__dfxtp_2 _41300_ (.CLK(clk),
    .D(_03794_),
    .Q(\count_cycle[63] ));
 sky130_fd_sc_hd__dfxtp_2 _41301_ (.CLK(clk),
    .D(_03795_),
    .Q(\timer[0] ));
 sky130_fd_sc_hd__dfxtp_2 _41302_ (.CLK(clk),
    .D(_03796_),
    .Q(\timer[1] ));
 sky130_fd_sc_hd__dfxtp_2 _41303_ (.CLK(clk),
    .D(_03797_),
    .Q(\timer[2] ));
 sky130_fd_sc_hd__dfxtp_2 _41304_ (.CLK(clk),
    .D(_03798_),
    .Q(\timer[3] ));
 sky130_fd_sc_hd__dfxtp_2 _41305_ (.CLK(clk),
    .D(_03799_),
    .Q(\timer[4] ));
 sky130_fd_sc_hd__dfxtp_2 _41306_ (.CLK(clk),
    .D(_03800_),
    .Q(\timer[5] ));
 sky130_fd_sc_hd__dfxtp_2 _41307_ (.CLK(clk),
    .D(_03801_),
    .Q(\timer[6] ));
 sky130_fd_sc_hd__dfxtp_2 _41308_ (.CLK(clk),
    .D(_03802_),
    .Q(\timer[7] ));
 sky130_fd_sc_hd__dfxtp_2 _41309_ (.CLK(clk),
    .D(_03803_),
    .Q(\timer[8] ));
 sky130_fd_sc_hd__dfxtp_2 _41310_ (.CLK(clk),
    .D(_03804_),
    .Q(\timer[9] ));
 sky130_fd_sc_hd__dfxtp_2 _41311_ (.CLK(clk),
    .D(_03805_),
    .Q(\timer[10] ));
 sky130_fd_sc_hd__dfxtp_2 _41312_ (.CLK(clk),
    .D(_03806_),
    .Q(\timer[11] ));
 sky130_fd_sc_hd__dfxtp_2 _41313_ (.CLK(clk),
    .D(_03807_),
    .Q(\timer[12] ));
 sky130_fd_sc_hd__dfxtp_2 _41314_ (.CLK(clk),
    .D(_03808_),
    .Q(\timer[13] ));
 sky130_fd_sc_hd__dfxtp_2 _41315_ (.CLK(clk),
    .D(_03809_),
    .Q(\timer[14] ));
 sky130_fd_sc_hd__dfxtp_2 _41316_ (.CLK(clk),
    .D(_03810_),
    .Q(\timer[15] ));
 sky130_fd_sc_hd__dfxtp_2 _41317_ (.CLK(clk),
    .D(_03811_),
    .Q(\timer[16] ));
 sky130_fd_sc_hd__dfxtp_2 _41318_ (.CLK(clk),
    .D(_03812_),
    .Q(\timer[17] ));
 sky130_fd_sc_hd__dfxtp_2 _41319_ (.CLK(clk),
    .D(_03813_),
    .Q(\timer[18] ));
 sky130_fd_sc_hd__dfxtp_2 _41320_ (.CLK(clk),
    .D(_03814_),
    .Q(\timer[19] ));
 sky130_fd_sc_hd__dfxtp_2 _41321_ (.CLK(clk),
    .D(_03815_),
    .Q(\timer[20] ));
 sky130_fd_sc_hd__dfxtp_2 _41322_ (.CLK(clk),
    .D(_03816_),
    .Q(\timer[21] ));
 sky130_fd_sc_hd__dfxtp_2 _41323_ (.CLK(clk),
    .D(_03817_),
    .Q(\timer[22] ));
 sky130_fd_sc_hd__dfxtp_2 _41324_ (.CLK(clk),
    .D(_03818_),
    .Q(\timer[23] ));
 sky130_fd_sc_hd__dfxtp_2 _41325_ (.CLK(clk),
    .D(_03819_),
    .Q(\timer[24] ));
 sky130_fd_sc_hd__dfxtp_2 _41326_ (.CLK(clk),
    .D(_03820_),
    .Q(\timer[25] ));
 sky130_fd_sc_hd__dfxtp_2 _41327_ (.CLK(clk),
    .D(_03821_),
    .Q(\timer[26] ));
 sky130_fd_sc_hd__dfxtp_2 _41328_ (.CLK(clk),
    .D(_03822_),
    .Q(\timer[27] ));
 sky130_fd_sc_hd__dfxtp_2 _41329_ (.CLK(clk),
    .D(_03823_),
    .Q(\timer[28] ));
 sky130_fd_sc_hd__dfxtp_2 _41330_ (.CLK(clk),
    .D(_03824_),
    .Q(\timer[29] ));
 sky130_fd_sc_hd__dfxtp_2 _41331_ (.CLK(clk),
    .D(_03825_),
    .Q(\timer[30] ));
 sky130_fd_sc_hd__dfxtp_2 _41332_ (.CLK(clk),
    .D(_03826_),
    .Q(\timer[31] ));
 sky130_fd_sc_hd__dfxtp_2 _41333_ (.CLK(clk),
    .D(_03827_),
    .Q(pcpi_timeout));
 sky130_fd_sc_hd__dfxtp_2 _41334_ (.CLK(clk),
    .D(_03828_),
    .Q(decoder_pseudo_trigger));
 sky130_fd_sc_hd__dfxtp_2 _41335_ (.CLK(clk),
    .D(_03829_),
    .Q(is_compare));
 sky130_fd_sc_hd__dfxtp_2 _41336_ (.CLK(clk),
    .D(_03830_),
    .Q(do_waitirq));
 sky130_fd_sc_hd__dfxtp_2 _41337_ (.CLK(clk),
    .D(_03831_),
    .Q(mem_valid));
 sky130_fd_sc_hd__dfxtp_2 _41338_ (.CLK(clk),
    .D(_03832_),
    .Q(pcpi_valid));
 sky130_fd_sc_hd__dfxtp_2 _41339_ (.CLK(clk),
    .D(_03833_),
    .Q(eoi[0]));
 sky130_fd_sc_hd__dfxtp_2 _41340_ (.CLK(clk),
    .D(_03834_),
    .Q(eoi[1]));
 sky130_fd_sc_hd__dfxtp_2 _41341_ (.CLK(clk),
    .D(_03835_),
    .Q(eoi[2]));
 sky130_fd_sc_hd__dfxtp_2 _41342_ (.CLK(clk),
    .D(_03836_),
    .Q(eoi[3]));
 sky130_fd_sc_hd__dfxtp_2 _41343_ (.CLK(clk),
    .D(_03837_),
    .Q(eoi[4]));
 sky130_fd_sc_hd__dfxtp_2 _41344_ (.CLK(clk),
    .D(_03838_),
    .Q(eoi[5]));
 sky130_fd_sc_hd__dfxtp_2 _41345_ (.CLK(clk),
    .D(_03839_),
    .Q(eoi[6]));
 sky130_fd_sc_hd__dfxtp_2 _41346_ (.CLK(clk),
    .D(_03840_),
    .Q(eoi[7]));
 sky130_fd_sc_hd__dfxtp_2 _41347_ (.CLK(clk),
    .D(_03841_),
    .Q(eoi[8]));
 sky130_fd_sc_hd__dfxtp_2 _41348_ (.CLK(clk),
    .D(_03842_),
    .Q(eoi[9]));
 sky130_fd_sc_hd__dfxtp_2 _41349_ (.CLK(clk),
    .D(_03843_),
    .Q(eoi[10]));
 sky130_fd_sc_hd__dfxtp_2 _41350_ (.CLK(clk),
    .D(_03844_),
    .Q(eoi[11]));
 sky130_fd_sc_hd__dfxtp_2 _41351_ (.CLK(clk),
    .D(_03845_),
    .Q(eoi[12]));
 sky130_fd_sc_hd__dfxtp_2 _41352_ (.CLK(clk),
    .D(_03846_),
    .Q(eoi[13]));
 sky130_fd_sc_hd__dfxtp_2 _41353_ (.CLK(clk),
    .D(_03847_),
    .Q(eoi[14]));
 sky130_fd_sc_hd__dfxtp_2 _41354_ (.CLK(clk),
    .D(_03848_),
    .Q(eoi[15]));
 sky130_fd_sc_hd__dfxtp_2 _41355_ (.CLK(clk),
    .D(_03849_),
    .Q(eoi[16]));
 sky130_fd_sc_hd__dfxtp_2 _41356_ (.CLK(clk),
    .D(_03850_),
    .Q(eoi[17]));
 sky130_fd_sc_hd__dfxtp_2 _41357_ (.CLK(clk),
    .D(_03851_),
    .Q(eoi[18]));
 sky130_fd_sc_hd__dfxtp_2 _41358_ (.CLK(clk),
    .D(_03852_),
    .Q(eoi[19]));
 sky130_fd_sc_hd__dfxtp_2 _41359_ (.CLK(clk),
    .D(_03853_),
    .Q(eoi[20]));
 sky130_fd_sc_hd__dfxtp_2 _41360_ (.CLK(clk),
    .D(_03854_),
    .Q(eoi[21]));
 sky130_fd_sc_hd__dfxtp_2 _41361_ (.CLK(clk),
    .D(_03855_),
    .Q(eoi[22]));
 sky130_fd_sc_hd__dfxtp_2 _41362_ (.CLK(clk),
    .D(_03856_),
    .Q(eoi[23]));
 sky130_fd_sc_hd__dfxtp_2 _41363_ (.CLK(clk),
    .D(_03857_),
    .Q(eoi[24]));
 sky130_fd_sc_hd__dfxtp_2 _41364_ (.CLK(clk),
    .D(_03858_),
    .Q(eoi[25]));
 sky130_fd_sc_hd__dfxtp_2 _41365_ (.CLK(clk),
    .D(_03859_),
    .Q(eoi[26]));
 sky130_fd_sc_hd__dfxtp_2 _41366_ (.CLK(clk),
    .D(_03860_),
    .Q(eoi[27]));
 sky130_fd_sc_hd__dfxtp_2 _41367_ (.CLK(clk),
    .D(_03861_),
    .Q(eoi[28]));
 sky130_fd_sc_hd__dfxtp_2 _41368_ (.CLK(clk),
    .D(_03862_),
    .Q(eoi[29]));
 sky130_fd_sc_hd__dfxtp_2 _41369_ (.CLK(clk),
    .D(_03863_),
    .Q(eoi[30]));
 sky130_fd_sc_hd__dfxtp_2 _41370_ (.CLK(clk),
    .D(_03864_),
    .Q(eoi[31]));
 sky130_fd_sc_hd__dfxtp_2 _41371_ (.CLK(clk),
    .D(_03865_),
    .Q(\count_instr[0] ));
 sky130_fd_sc_hd__dfxtp_2 _41372_ (.CLK(clk),
    .D(_03866_),
    .Q(\count_instr[1] ));
 sky130_fd_sc_hd__dfxtp_2 _41373_ (.CLK(clk),
    .D(_03867_),
    .Q(\count_instr[2] ));
 sky130_fd_sc_hd__dfxtp_2 _41374_ (.CLK(clk),
    .D(_03868_),
    .Q(\count_instr[3] ));
 sky130_fd_sc_hd__dfxtp_2 _41375_ (.CLK(clk),
    .D(_03869_),
    .Q(\count_instr[4] ));
 sky130_fd_sc_hd__dfxtp_2 _41376_ (.CLK(clk),
    .D(_03870_),
    .Q(\count_instr[5] ));
 sky130_fd_sc_hd__dfxtp_2 _41377_ (.CLK(clk),
    .D(_03871_),
    .Q(\count_instr[6] ));
 sky130_fd_sc_hd__dfxtp_2 _41378_ (.CLK(clk),
    .D(_03872_),
    .Q(\count_instr[7] ));
 sky130_fd_sc_hd__dfxtp_2 _41379_ (.CLK(clk),
    .D(_03873_),
    .Q(\count_instr[8] ));
 sky130_fd_sc_hd__dfxtp_2 _41380_ (.CLK(clk),
    .D(_03874_),
    .Q(\count_instr[9] ));
 sky130_fd_sc_hd__dfxtp_2 _41381_ (.CLK(clk),
    .D(_03875_),
    .Q(\count_instr[10] ));
 sky130_fd_sc_hd__dfxtp_2 _41382_ (.CLK(clk),
    .D(_03876_),
    .Q(\count_instr[11] ));
 sky130_fd_sc_hd__dfxtp_2 _41383_ (.CLK(clk),
    .D(_03877_),
    .Q(\count_instr[12] ));
 sky130_fd_sc_hd__dfxtp_2 _41384_ (.CLK(clk),
    .D(_03878_),
    .Q(\count_instr[13] ));
 sky130_fd_sc_hd__dfxtp_2 _41385_ (.CLK(clk),
    .D(_03879_),
    .Q(\count_instr[14] ));
 sky130_fd_sc_hd__dfxtp_2 _41386_ (.CLK(clk),
    .D(_03880_),
    .Q(\count_instr[15] ));
 sky130_fd_sc_hd__dfxtp_2 _41387_ (.CLK(clk),
    .D(_03881_),
    .Q(\count_instr[16] ));
 sky130_fd_sc_hd__dfxtp_2 _41388_ (.CLK(clk),
    .D(_03882_),
    .Q(\count_instr[17] ));
 sky130_fd_sc_hd__dfxtp_2 _41389_ (.CLK(clk),
    .D(_03883_),
    .Q(\count_instr[18] ));
 sky130_fd_sc_hd__dfxtp_2 _41390_ (.CLK(clk),
    .D(_03884_),
    .Q(\count_instr[19] ));
 sky130_fd_sc_hd__dfxtp_2 _41391_ (.CLK(clk),
    .D(_03885_),
    .Q(\count_instr[20] ));
 sky130_fd_sc_hd__dfxtp_2 _41392_ (.CLK(clk),
    .D(_03886_),
    .Q(\count_instr[21] ));
 sky130_fd_sc_hd__dfxtp_2 _41393_ (.CLK(clk),
    .D(_03887_),
    .Q(\count_instr[22] ));
 sky130_fd_sc_hd__dfxtp_2 _41394_ (.CLK(clk),
    .D(_03888_),
    .Q(\count_instr[23] ));
 sky130_fd_sc_hd__dfxtp_2 _41395_ (.CLK(clk),
    .D(_03889_),
    .Q(\count_instr[24] ));
 sky130_fd_sc_hd__dfxtp_2 _41396_ (.CLK(clk),
    .D(_03890_),
    .Q(\count_instr[25] ));
 sky130_fd_sc_hd__dfxtp_2 _41397_ (.CLK(clk),
    .D(_03891_),
    .Q(\count_instr[26] ));
 sky130_fd_sc_hd__dfxtp_2 _41398_ (.CLK(clk),
    .D(_03892_),
    .Q(\count_instr[27] ));
 sky130_fd_sc_hd__dfxtp_2 _41399_ (.CLK(clk),
    .D(_03893_),
    .Q(\count_instr[28] ));
 sky130_fd_sc_hd__dfxtp_2 _41400_ (.CLK(clk),
    .D(_03894_),
    .Q(\count_instr[29] ));
 sky130_fd_sc_hd__dfxtp_2 _41401_ (.CLK(clk),
    .D(_03895_),
    .Q(\count_instr[30] ));
 sky130_fd_sc_hd__dfxtp_2 _41402_ (.CLK(clk),
    .D(_03896_),
    .Q(\count_instr[31] ));
 sky130_fd_sc_hd__dfxtp_2 _41403_ (.CLK(clk),
    .D(_03897_),
    .Q(\count_instr[32] ));
 sky130_fd_sc_hd__dfxtp_2 _41404_ (.CLK(clk),
    .D(_03898_),
    .Q(\count_instr[33] ));
 sky130_fd_sc_hd__dfxtp_2 _41405_ (.CLK(clk),
    .D(_03899_),
    .Q(\count_instr[34] ));
 sky130_fd_sc_hd__dfxtp_2 _41406_ (.CLK(clk),
    .D(_03900_),
    .Q(\count_instr[35] ));
 sky130_fd_sc_hd__dfxtp_2 _41407_ (.CLK(clk),
    .D(_03901_),
    .Q(\count_instr[36] ));
 sky130_fd_sc_hd__dfxtp_2 _41408_ (.CLK(clk),
    .D(_03902_),
    .Q(\count_instr[37] ));
 sky130_fd_sc_hd__dfxtp_2 _41409_ (.CLK(clk),
    .D(_03903_),
    .Q(\count_instr[38] ));
 sky130_fd_sc_hd__dfxtp_2 _41410_ (.CLK(clk),
    .D(_03904_),
    .Q(\count_instr[39] ));
 sky130_fd_sc_hd__dfxtp_2 _41411_ (.CLK(clk),
    .D(_03905_),
    .Q(\count_instr[40] ));
 sky130_fd_sc_hd__dfxtp_2 _41412_ (.CLK(clk),
    .D(_03906_),
    .Q(\count_instr[41] ));
 sky130_fd_sc_hd__dfxtp_2 _41413_ (.CLK(clk),
    .D(_03907_),
    .Q(\count_instr[42] ));
 sky130_fd_sc_hd__dfxtp_2 _41414_ (.CLK(clk),
    .D(_03908_),
    .Q(\count_instr[43] ));
 sky130_fd_sc_hd__dfxtp_2 _41415_ (.CLK(clk),
    .D(_03909_),
    .Q(\count_instr[44] ));
 sky130_fd_sc_hd__dfxtp_2 _41416_ (.CLK(clk),
    .D(_03910_),
    .Q(\count_instr[45] ));
 sky130_fd_sc_hd__dfxtp_2 _41417_ (.CLK(clk),
    .D(_03911_),
    .Q(\count_instr[46] ));
 sky130_fd_sc_hd__dfxtp_2 _41418_ (.CLK(clk),
    .D(_03912_),
    .Q(\count_instr[47] ));
 sky130_fd_sc_hd__dfxtp_2 _41419_ (.CLK(clk),
    .D(_03913_),
    .Q(\count_instr[48] ));
 sky130_fd_sc_hd__dfxtp_2 _41420_ (.CLK(clk),
    .D(_03914_),
    .Q(\count_instr[49] ));
 sky130_fd_sc_hd__dfxtp_2 _41421_ (.CLK(clk),
    .D(_03915_),
    .Q(\count_instr[50] ));
 sky130_fd_sc_hd__dfxtp_2 _41422_ (.CLK(clk),
    .D(_03916_),
    .Q(\count_instr[51] ));
 sky130_fd_sc_hd__dfxtp_2 _41423_ (.CLK(clk),
    .D(_03917_),
    .Q(\count_instr[52] ));
 sky130_fd_sc_hd__dfxtp_2 _41424_ (.CLK(clk),
    .D(_03918_),
    .Q(\count_instr[53] ));
 sky130_fd_sc_hd__dfxtp_2 _41425_ (.CLK(clk),
    .D(_03919_),
    .Q(\count_instr[54] ));
 sky130_fd_sc_hd__dfxtp_2 _41426_ (.CLK(clk),
    .D(_03920_),
    .Q(\count_instr[55] ));
 sky130_fd_sc_hd__dfxtp_2 _41427_ (.CLK(clk),
    .D(_03921_),
    .Q(\count_instr[56] ));
 sky130_fd_sc_hd__dfxtp_2 _41428_ (.CLK(clk),
    .D(_03922_),
    .Q(\count_instr[57] ));
 sky130_fd_sc_hd__dfxtp_2 _41429_ (.CLK(clk),
    .D(_03923_),
    .Q(\count_instr[58] ));
 sky130_fd_sc_hd__dfxtp_2 _41430_ (.CLK(clk),
    .D(_03924_),
    .Q(\count_instr[59] ));
 sky130_fd_sc_hd__dfxtp_2 _41431_ (.CLK(clk),
    .D(_03925_),
    .Q(\count_instr[60] ));
 sky130_fd_sc_hd__dfxtp_2 _41432_ (.CLK(clk),
    .D(_03926_),
    .Q(\count_instr[61] ));
 sky130_fd_sc_hd__dfxtp_2 _41433_ (.CLK(clk),
    .D(_03927_),
    .Q(\count_instr[62] ));
 sky130_fd_sc_hd__dfxtp_2 _41434_ (.CLK(clk),
    .D(_03928_),
    .Q(\count_instr[63] ));
 sky130_fd_sc_hd__dfxtp_2 _41435_ (.CLK(clk),
    .D(_03929_),
    .Q(\reg_pc[1] ));
 sky130_fd_sc_hd__dfxtp_2 _41436_ (.CLK(clk),
    .D(_03930_),
    .Q(\reg_pc[2] ));
 sky130_fd_sc_hd__dfxtp_2 _41437_ (.CLK(clk),
    .D(_03931_),
    .Q(\reg_pc[3] ));
 sky130_fd_sc_hd__dfxtp_2 _41438_ (.CLK(clk),
    .D(_03932_),
    .Q(\reg_pc[4] ));
 sky130_fd_sc_hd__dfxtp_2 _41439_ (.CLK(clk),
    .D(_03933_),
    .Q(\reg_pc[5] ));
 sky130_fd_sc_hd__dfxtp_2 _41440_ (.CLK(clk),
    .D(_03934_),
    .Q(\reg_pc[6] ));
 sky130_fd_sc_hd__dfxtp_2 _41441_ (.CLK(clk),
    .D(_03935_),
    .Q(\reg_pc[7] ));
 sky130_fd_sc_hd__dfxtp_2 _41442_ (.CLK(clk),
    .D(_03936_),
    .Q(\reg_pc[8] ));
 sky130_fd_sc_hd__dfxtp_2 _41443_ (.CLK(clk),
    .D(_03937_),
    .Q(\reg_pc[9] ));
 sky130_fd_sc_hd__dfxtp_2 _41444_ (.CLK(clk),
    .D(_03938_),
    .Q(\reg_pc[10] ));
 sky130_fd_sc_hd__dfxtp_2 _41445_ (.CLK(clk),
    .D(_03939_),
    .Q(\reg_pc[11] ));
 sky130_fd_sc_hd__dfxtp_2 _41446_ (.CLK(clk),
    .D(_03940_),
    .Q(\reg_pc[12] ));
 sky130_fd_sc_hd__dfxtp_2 _41447_ (.CLK(clk),
    .D(_03941_),
    .Q(\reg_pc[13] ));
 sky130_fd_sc_hd__dfxtp_2 _41448_ (.CLK(clk),
    .D(_03942_),
    .Q(\reg_pc[14] ));
 sky130_fd_sc_hd__dfxtp_2 _41449_ (.CLK(clk),
    .D(_03943_),
    .Q(\reg_pc[15] ));
 sky130_fd_sc_hd__dfxtp_2 _41450_ (.CLK(clk),
    .D(_03944_),
    .Q(\reg_pc[16] ));
 sky130_fd_sc_hd__dfxtp_2 _41451_ (.CLK(clk),
    .D(_03945_),
    .Q(\reg_pc[17] ));
 sky130_fd_sc_hd__dfxtp_2 _41452_ (.CLK(clk),
    .D(_03946_),
    .Q(\reg_pc[18] ));
 sky130_fd_sc_hd__dfxtp_2 _41453_ (.CLK(clk),
    .D(_03947_),
    .Q(\reg_pc[19] ));
 sky130_fd_sc_hd__dfxtp_2 _41454_ (.CLK(clk),
    .D(_03948_),
    .Q(\reg_pc[20] ));
 sky130_fd_sc_hd__dfxtp_2 _41455_ (.CLK(clk),
    .D(_03949_),
    .Q(\reg_pc[21] ));
 sky130_fd_sc_hd__dfxtp_2 _41456_ (.CLK(clk),
    .D(_03950_),
    .Q(\reg_pc[22] ));
 sky130_fd_sc_hd__dfxtp_2 _41457_ (.CLK(clk),
    .D(_03951_),
    .Q(\reg_pc[23] ));
 sky130_fd_sc_hd__dfxtp_2 _41458_ (.CLK(clk),
    .D(_03952_),
    .Q(\reg_pc[24] ));
 sky130_fd_sc_hd__dfxtp_2 _41459_ (.CLK(clk),
    .D(_03953_),
    .Q(\reg_pc[25] ));
 sky130_fd_sc_hd__dfxtp_2 _41460_ (.CLK(clk),
    .D(_03954_),
    .Q(\reg_pc[26] ));
 sky130_fd_sc_hd__dfxtp_2 _41461_ (.CLK(clk),
    .D(_03955_),
    .Q(\reg_pc[27] ));
 sky130_fd_sc_hd__dfxtp_2 _41462_ (.CLK(clk),
    .D(_03956_),
    .Q(\reg_pc[28] ));
 sky130_fd_sc_hd__dfxtp_2 _41463_ (.CLK(clk),
    .D(_03957_),
    .Q(\reg_pc[29] ));
 sky130_fd_sc_hd__dfxtp_2 _41464_ (.CLK(clk),
    .D(_03958_),
    .Q(\reg_pc[30] ));
 sky130_fd_sc_hd__dfxtp_2 _41465_ (.CLK(clk),
    .D(_03959_),
    .Q(\reg_pc[31] ));
 sky130_fd_sc_hd__dfxtp_2 _41466_ (.CLK(clk),
    .D(_03960_),
    .Q(\reg_next_pc[1] ));
 sky130_fd_sc_hd__dfxtp_2 _41467_ (.CLK(clk),
    .D(_03961_),
    .Q(\reg_next_pc[2] ));
 sky130_fd_sc_hd__dfxtp_2 _41468_ (.CLK(clk),
    .D(_03962_),
    .Q(\reg_next_pc[3] ));
 sky130_fd_sc_hd__dfxtp_2 _41469_ (.CLK(clk),
    .D(_03963_),
    .Q(\reg_next_pc[4] ));
 sky130_fd_sc_hd__dfxtp_2 _41470_ (.CLK(clk),
    .D(_03964_),
    .Q(\reg_next_pc[5] ));
 sky130_fd_sc_hd__dfxtp_2 _41471_ (.CLK(clk),
    .D(_03965_),
    .Q(\reg_next_pc[6] ));
 sky130_fd_sc_hd__dfxtp_2 _41472_ (.CLK(clk),
    .D(_03966_),
    .Q(\reg_next_pc[7] ));
 sky130_fd_sc_hd__dfxtp_2 _41473_ (.CLK(clk),
    .D(_03967_),
    .Q(\reg_next_pc[8] ));
 sky130_fd_sc_hd__dfxtp_2 _41474_ (.CLK(clk),
    .D(_03968_),
    .Q(\reg_next_pc[9] ));
 sky130_fd_sc_hd__dfxtp_2 _41475_ (.CLK(clk),
    .D(_03969_),
    .Q(\reg_next_pc[10] ));
 sky130_fd_sc_hd__dfxtp_2 _41476_ (.CLK(clk),
    .D(_03970_),
    .Q(\reg_next_pc[11] ));
 sky130_fd_sc_hd__dfxtp_2 _41477_ (.CLK(clk),
    .D(_03971_),
    .Q(\reg_next_pc[12] ));
 sky130_fd_sc_hd__dfxtp_2 _41478_ (.CLK(clk),
    .D(_03972_),
    .Q(\reg_next_pc[13] ));
 sky130_fd_sc_hd__dfxtp_2 _41479_ (.CLK(clk),
    .D(_03973_),
    .Q(\reg_next_pc[14] ));
 sky130_fd_sc_hd__dfxtp_2 _41480_ (.CLK(clk),
    .D(_03974_),
    .Q(\reg_next_pc[15] ));
 sky130_fd_sc_hd__dfxtp_2 _41481_ (.CLK(clk),
    .D(_03975_),
    .Q(\reg_next_pc[16] ));
 sky130_fd_sc_hd__dfxtp_2 _41482_ (.CLK(clk),
    .D(_03976_),
    .Q(\reg_next_pc[17] ));
 sky130_fd_sc_hd__dfxtp_2 _41483_ (.CLK(clk),
    .D(_03977_),
    .Q(\reg_next_pc[18] ));
 sky130_fd_sc_hd__dfxtp_2 _41484_ (.CLK(clk),
    .D(_03978_),
    .Q(\reg_next_pc[19] ));
 sky130_fd_sc_hd__dfxtp_2 _41485_ (.CLK(clk),
    .D(_03979_),
    .Q(\reg_next_pc[20] ));
 sky130_fd_sc_hd__dfxtp_2 _41486_ (.CLK(clk),
    .D(_03980_),
    .Q(\reg_next_pc[21] ));
 sky130_fd_sc_hd__dfxtp_2 _41487_ (.CLK(clk),
    .D(_03981_),
    .Q(\reg_next_pc[22] ));
 sky130_fd_sc_hd__dfxtp_2 _41488_ (.CLK(clk),
    .D(_03982_),
    .Q(\reg_next_pc[23] ));
 sky130_fd_sc_hd__dfxtp_2 _41489_ (.CLK(clk),
    .D(_03983_),
    .Q(\reg_next_pc[24] ));
 sky130_fd_sc_hd__dfxtp_2 _41490_ (.CLK(clk),
    .D(_03984_),
    .Q(\reg_next_pc[25] ));
 sky130_fd_sc_hd__dfxtp_2 _41491_ (.CLK(clk),
    .D(_03985_),
    .Q(\reg_next_pc[26] ));
 sky130_fd_sc_hd__dfxtp_2 _41492_ (.CLK(clk),
    .D(_03986_),
    .Q(\reg_next_pc[27] ));
 sky130_fd_sc_hd__dfxtp_2 _41493_ (.CLK(clk),
    .D(_03987_),
    .Q(\reg_next_pc[28] ));
 sky130_fd_sc_hd__dfxtp_2 _41494_ (.CLK(clk),
    .D(_03988_),
    .Q(\reg_next_pc[29] ));
 sky130_fd_sc_hd__dfxtp_2 _41495_ (.CLK(clk),
    .D(_03989_),
    .Q(\reg_next_pc[30] ));
 sky130_fd_sc_hd__dfxtp_2 _41496_ (.CLK(clk),
    .D(_03990_),
    .Q(\reg_next_pc[31] ));
 sky130_fd_sc_hd__dfxtp_2 _41497_ (.CLK(clk),
    .D(_03991_),
    .Q(mem_do_rdata));
 sky130_fd_sc_hd__dfxtp_2 _41498_ (.CLK(clk),
    .D(_03992_),
    .Q(mem_do_wdata));
 sky130_fd_sc_hd__dfxtp_2 _41499_ (.CLK(clk),
    .D(_03993_),
    .Q(\pcpi_timeout_counter[0] ));
 sky130_fd_sc_hd__dfxtp_2 _41500_ (.CLK(clk),
    .D(_03994_),
    .Q(\pcpi_timeout_counter[1] ));
 sky130_fd_sc_hd__dfxtp_2 _41501_ (.CLK(clk),
    .D(_03995_),
    .Q(\pcpi_timeout_counter[2] ));
 sky130_fd_sc_hd__dfxtp_2 _41502_ (.CLK(clk),
    .D(_03996_),
    .Q(\pcpi_timeout_counter[3] ));
 sky130_fd_sc_hd__dfxtp_2 _41503_ (.CLK(clk),
    .D(_03997_),
    .Q(instr_beq));
 sky130_fd_sc_hd__dfxtp_2 _41504_ (.CLK(clk),
    .D(_03998_),
    .Q(instr_bne));
 sky130_fd_sc_hd__dfxtp_2 _41505_ (.CLK(clk),
    .D(_03999_),
    .Q(instr_blt));
 sky130_fd_sc_hd__dfxtp_2 _41506_ (.CLK(clk),
    .D(_04000_),
    .Q(instr_bge));
 sky130_fd_sc_hd__dfxtp_2 _41507_ (.CLK(clk),
    .D(_04001_),
    .Q(instr_bltu));
 sky130_fd_sc_hd__dfxtp_2 _41508_ (.CLK(clk),
    .D(_04002_),
    .Q(instr_bgeu));
 sky130_fd_sc_hd__dfxtp_2 _41509_ (.CLK(clk),
    .D(_04003_),
    .Q(instr_addi));
 sky130_fd_sc_hd__dfxtp_2 _41510_ (.CLK(clk),
    .D(_04004_),
    .Q(instr_slti));
 sky130_fd_sc_hd__dfxtp_2 _41511_ (.CLK(clk),
    .D(_04005_),
    .Q(instr_sltiu));
 sky130_fd_sc_hd__dfxtp_2 _41512_ (.CLK(clk),
    .D(_04006_),
    .Q(instr_xori));
 sky130_fd_sc_hd__dfxtp_2 _41513_ (.CLK(clk),
    .D(_04007_),
    .Q(instr_ori));
 sky130_fd_sc_hd__dfxtp_2 _41514_ (.CLK(clk),
    .D(_04008_),
    .Q(instr_andi));
 sky130_fd_sc_hd__dfxtp_2 _41515_ (.CLK(clk),
    .D(_04009_),
    .Q(instr_add));
 sky130_fd_sc_hd__dfxtp_2 _41516_ (.CLK(clk),
    .D(_04010_),
    .Q(instr_sub));
 sky130_fd_sc_hd__dfxtp_2 _41517_ (.CLK(clk),
    .D(_04011_),
    .Q(instr_sll));
 sky130_fd_sc_hd__dfxtp_2 _41518_ (.CLK(clk),
    .D(_04012_),
    .Q(instr_slt));
 sky130_fd_sc_hd__dfxtp_2 _41519_ (.CLK(clk),
    .D(_04013_),
    .Q(instr_sltu));
 sky130_fd_sc_hd__dfxtp_2 _41520_ (.CLK(clk),
    .D(_04014_),
    .Q(instr_xor));
 sky130_fd_sc_hd__dfxtp_2 _41521_ (.CLK(clk),
    .D(_04015_),
    .Q(instr_srl));
 sky130_fd_sc_hd__dfxtp_2 _41522_ (.CLK(clk),
    .D(_04016_),
    .Q(instr_sra));
 sky130_fd_sc_hd__dfxtp_2 _41523_ (.CLK(clk),
    .D(_04017_),
    .Q(instr_or));
 sky130_fd_sc_hd__dfxtp_2 _41524_ (.CLK(clk),
    .D(_04018_),
    .Q(instr_and));
 sky130_fd_sc_hd__dfxtp_2 _41525_ (.CLK(clk),
    .D(_04019_),
    .Q(\decoded_rs1[0] ));
 sky130_fd_sc_hd__dfxtp_2 _41526_ (.CLK(clk),
    .D(_04020_),
    .Q(\decoded_rs1[1] ));
 sky130_fd_sc_hd__dfxtp_2 _41527_ (.CLK(clk),
    .D(_04021_),
    .Q(\decoded_rs1[2] ));
 sky130_fd_sc_hd__dfxtp_2 _41528_ (.CLK(clk),
    .D(_04022_),
    .Q(\decoded_rs1[3] ));
 sky130_fd_sc_hd__dfxtp_2 _41529_ (.CLK(clk),
    .D(_04023_),
    .Q(is_beq_bne_blt_bge_bltu_bgeu));
 sky130_fd_sc_hd__dfxtp_2 _41530_ (.CLK(clk),
    .D(_04024_),
    .Q(mem_instr));
 sky130_fd_sc_hd__dfxtp_2 _41531_ (.CLK(clk),
    .D(_04025_),
    .Q(\irq_mask[0] ));
 sky130_fd_sc_hd__dfxtp_2 _41532_ (.CLK(clk),
    .D(_04026_),
    .Q(\irq_mask[1] ));
 sky130_fd_sc_hd__dfxtp_2 _41533_ (.CLK(clk),
    .D(_04027_),
    .Q(\irq_mask[2] ));
 sky130_fd_sc_hd__dfxtp_2 _41534_ (.CLK(clk),
    .D(_04028_),
    .Q(\irq_mask[3] ));
 sky130_fd_sc_hd__dfxtp_2 _41535_ (.CLK(clk),
    .D(_04029_),
    .Q(\irq_mask[4] ));
 sky130_fd_sc_hd__dfxtp_2 _41536_ (.CLK(clk),
    .D(_04030_),
    .Q(\irq_mask[5] ));
 sky130_fd_sc_hd__dfxtp_2 _41537_ (.CLK(clk),
    .D(_04031_),
    .Q(\irq_mask[6] ));
 sky130_fd_sc_hd__dfxtp_2 _41538_ (.CLK(clk),
    .D(_04032_),
    .Q(\irq_mask[7] ));
 sky130_fd_sc_hd__dfxtp_2 _41539_ (.CLK(clk),
    .D(_04033_),
    .Q(\irq_mask[8] ));
 sky130_fd_sc_hd__dfxtp_2 _41540_ (.CLK(clk),
    .D(_04034_),
    .Q(\irq_mask[9] ));
 sky130_fd_sc_hd__dfxtp_2 _41541_ (.CLK(clk),
    .D(_04035_),
    .Q(\irq_mask[10] ));
 sky130_fd_sc_hd__dfxtp_2 _41542_ (.CLK(clk),
    .D(_04036_),
    .Q(\irq_mask[11] ));
 sky130_fd_sc_hd__dfxtp_2 _41543_ (.CLK(clk),
    .D(_04037_),
    .Q(\irq_mask[12] ));
 sky130_fd_sc_hd__dfxtp_2 _41544_ (.CLK(clk),
    .D(_04038_),
    .Q(\irq_mask[13] ));
 sky130_fd_sc_hd__dfxtp_2 _41545_ (.CLK(clk),
    .D(_04039_),
    .Q(\irq_mask[14] ));
 sky130_fd_sc_hd__dfxtp_2 _41546_ (.CLK(clk),
    .D(_04040_),
    .Q(\irq_mask[15] ));
 sky130_fd_sc_hd__dfxtp_2 _41547_ (.CLK(clk),
    .D(_04041_),
    .Q(\irq_mask[16] ));
 sky130_fd_sc_hd__dfxtp_2 _41548_ (.CLK(clk),
    .D(_04042_),
    .Q(\irq_mask[17] ));
 sky130_fd_sc_hd__dfxtp_2 _41549_ (.CLK(clk),
    .D(_04043_),
    .Q(\irq_mask[18] ));
 sky130_fd_sc_hd__dfxtp_2 _41550_ (.CLK(clk),
    .D(_04044_),
    .Q(\irq_mask[19] ));
 sky130_fd_sc_hd__dfxtp_2 _41551_ (.CLK(clk),
    .D(_04045_),
    .Q(\irq_mask[20] ));
 sky130_fd_sc_hd__dfxtp_2 _41552_ (.CLK(clk),
    .D(_04046_),
    .Q(\irq_mask[21] ));
 sky130_fd_sc_hd__dfxtp_2 _41553_ (.CLK(clk),
    .D(_04047_),
    .Q(\irq_mask[22] ));
 sky130_fd_sc_hd__dfxtp_2 _41554_ (.CLK(clk),
    .D(_04048_),
    .Q(\irq_mask[23] ));
 sky130_fd_sc_hd__dfxtp_2 _41555_ (.CLK(clk),
    .D(_04049_),
    .Q(\irq_mask[24] ));
 sky130_fd_sc_hd__dfxtp_2 _41556_ (.CLK(clk),
    .D(_04050_),
    .Q(\irq_mask[25] ));
 sky130_fd_sc_hd__dfxtp_2 _41557_ (.CLK(clk),
    .D(_04051_),
    .Q(\irq_mask[26] ));
 sky130_fd_sc_hd__dfxtp_2 _41558_ (.CLK(clk),
    .D(_04052_),
    .Q(\irq_mask[27] ));
 sky130_fd_sc_hd__dfxtp_2 _41559_ (.CLK(clk),
    .D(_04053_),
    .Q(\irq_mask[28] ));
 sky130_fd_sc_hd__dfxtp_2 _41560_ (.CLK(clk),
    .D(_04054_),
    .Q(\irq_mask[29] ));
 sky130_fd_sc_hd__dfxtp_2 _41561_ (.CLK(clk),
    .D(_04055_),
    .Q(\irq_mask[30] ));
 sky130_fd_sc_hd__dfxtp_2 _41562_ (.CLK(clk),
    .D(_04056_),
    .Q(\irq_mask[31] ));
 sky130_fd_sc_hd__dfxtp_2 _41563_ (.CLK(clk),
    .D(_04057_),
    .Q(mem_do_prefetch));
 sky130_fd_sc_hd__dfxtp_2 _41564_ (.CLK(clk),
    .D(_04058_),
    .Q(mem_do_rinst));
 sky130_fd_sc_hd__dfxtp_2 _41565_ (.CLK(clk),
    .D(_04059_),
    .Q(\irq_state[0] ));
 sky130_fd_sc_hd__dfxtp_2 _41566_ (.CLK(clk),
    .D(_04060_),
    .Q(\irq_state[1] ));
 sky130_fd_sc_hd__dfxtp_2 _41567_ (.CLK(clk),
    .D(_04061_),
    .Q(latched_store));
 sky130_fd_sc_hd__dfxtp_2 _41568_ (.CLK(clk),
    .D(_04062_),
    .Q(latched_stalu));
 sky130_fd_sc_hd__dfxtp_2 _41569_ (.CLK(clk),
    .D(_04063_),
    .Q(\pcpi_mul.rs2[32] ));
 sky130_fd_sc_hd__dfxtp_2 _41570_ (.CLK(clk),
    .D(_04064_),
    .Q(\pcpi_mul.rs1[32] ));
 sky130_fd_sc_hd__dfxtp_2 _41571_ (.CLK(clk),
    .D(_04065_),
    .Q(irq_delay));
 sky130_fd_sc_hd__dfxtp_2 _41572_ (.CLK(clk),
    .D(_04066_),
    .Q(\decoded_rs1[4] ));
 sky130_fd_sc_hd__dfxtp_2 _41573_ (.CLK(clk),
    .D(_04067_),
    .Q(\mem_state[0] ));
 sky130_fd_sc_hd__dfxtp_2 _41574_ (.CLK(clk),
    .D(_04068_),
    .Q(\mem_state[1] ));
 sky130_fd_sc_hd__dfxtp_2 _41575_ (.CLK(clk),
    .D(_04069_),
    .Q(latched_branch));
 sky130_fd_sc_hd__dfxtp_2 _41576_ (.CLK(clk),
    .D(_04070_),
    .Q(latched_is_lh));
 sky130_fd_sc_hd__dfxtp_2 _41577_ (.CLK(clk),
    .D(_04071_),
    .Q(latched_is_lb));
 sky130_fd_sc_hd__dfxtp_2 _41578_ (.CLK(clk),
    .D(_04072_),
    .Q(irq_active));
endmodule
