module picorv32a (clk,
    mem_instr,
    mem_la_read,
    mem_la_write,
    mem_ready,
    mem_valid,
    pcpi_ready,
    pcpi_valid,
    pcpi_wait,
    pcpi_wr,
    resetn,
    trace_valid,
    trap,
    eoi,
    irq,
    mem_addr,
    mem_la_addr,
    mem_la_wdata,
    mem_la_wstrb,
    mem_rdata,
    mem_wdata,
    mem_wstrb,
    pcpi_insn,
    pcpi_rd,
    pcpi_rs1,
    pcpi_rs2,
    trace_data);
 input clk;
 output mem_instr;
 output mem_la_read;
 output mem_la_write;
 input mem_ready;
 output mem_valid;
 input pcpi_ready;
 output pcpi_valid;
 input pcpi_wait;
 input pcpi_wr;
 input resetn;
 output trace_valid;
 output trap;
 output [31:0] eoi;
 input [31:0] irq;
 output [31:0] mem_addr;
 output [31:0] mem_la_addr;
 output [31:0] mem_la_wdata;
 output [3:0] mem_la_wstrb;
 input [31:0] mem_rdata;
 output [31:0] mem_wdata;
 output [3:0] mem_wstrb;
 output [31:0] pcpi_insn;
 input [31:0] pcpi_rd;
 output [31:0] pcpi_rs1;
 output [31:0] pcpi_rs2;
 output [35:0] trace_data;

 sky130_fd_sc_hd__clkbuf_2 _14370_ (.A(net101),
    .X(_11542_));
 sky130_fd_sc_hd__clkbuf_4 _14371_ (.A(_11542_),
    .X(_11543_));
 sky130_fd_sc_hd__clkbuf_2 _14372_ (.A(_11543_),
    .X(_11544_));
 sky130_fd_sc_hd__buf_1 _14373_ (.A(mem_do_prefetch),
    .X(_11545_));
 sky130_fd_sc_hd__nand2_2 _14374_ (.A(net237),
    .B(net65),
    .Y(_11546_));
 sky130_vsdinv _14375_ (.A(_11546_),
    .Y(_11547_));
 sky130_vsdinv _14376_ (.A(\mem_state[1] ),
    .Y(_11548_));
 sky130_vsdinv _14377_ (.A(\mem_state[0] ),
    .Y(_11549_));
 sky130_fd_sc_hd__nor2_1 _14378_ (.A(_11548_),
    .B(_11549_),
    .Y(_11550_));
 sky130_fd_sc_hd__buf_1 _14379_ (.A(mem_do_rinst),
    .X(_11551_));
 sky130_fd_sc_hd__o21a_1 _14380_ (.A1(mem_do_wdata),
    .A2(mem_do_rdata),
    .B1(_11547_),
    .X(_11552_));
 sky130_fd_sc_hd__or2_1 _14381_ (.A(\mem_state[1] ),
    .B(\mem_state[0] ),
    .X(_11553_));
 sky130_fd_sc_hd__o221a_1 _14382_ (.A1(_11547_),
    .A2(_11550_),
    .B1(_11551_),
    .B2(_11552_),
    .C1(_11553_),
    .X(_11554_));
 sky130_fd_sc_hd__nand2_2 _14383_ (.A(_11542_),
    .B(_11554_),
    .Y(_11555_));
 sky130_fd_sc_hd__nand2_1 _14384_ (.A(_11545_),
    .B(_11555_),
    .Y(_11556_));
 sky130_fd_sc_hd__buf_1 _14385_ (.A(mem_do_rdata),
    .X(_11557_));
 sky130_vsdinv _14386_ (.A(_11557_),
    .Y(_11558_));
 sky130_vsdinv _14387_ (.A(\cpu_state[6] ),
    .Y(_11559_));
 sky130_fd_sc_hd__buf_2 _14388_ (.A(_11559_),
    .X(_11560_));
 sky130_fd_sc_hd__nor2_1 _14389_ (.A(_11558_),
    .B(_11560_),
    .Y(_00319_));
 sky130_fd_sc_hd__a31o_1 _14390_ (.A1(_11544_),
    .A2(_11556_),
    .A3(_00319_),
    .B1(_00332_),
    .X(_11561_));
 sky130_vsdinv _14391_ (.A(_11561_),
    .Y(_11562_));
 sky130_fd_sc_hd__buf_1 _14392_ (.A(\cpu_state[6] ),
    .X(_11563_));
 sky130_fd_sc_hd__and2_1 _14393_ (.A(instr_lb),
    .B(_11563_),
    .X(_11564_));
 sky130_fd_sc_hd__buf_1 _14394_ (.A(_11544_),
    .X(_11565_));
 sky130_fd_sc_hd__buf_2 _14395_ (.A(_11565_),
    .X(_11566_));
 sky130_fd_sc_hd__o221a_1 _14396_ (.A1(latched_is_lb),
    .A2(_11562_),
    .B1(_11561_),
    .B2(_11564_),
    .C1(_11566_),
    .X(_04071_));
 sky130_fd_sc_hd__and2_1 _14397_ (.A(instr_lh),
    .B(_11563_),
    .X(_11567_));
 sky130_fd_sc_hd__o221a_1 _14398_ (.A1(latched_is_lh),
    .A2(_11562_),
    .B1(_11561_),
    .B2(_11567_),
    .C1(_11566_),
    .X(_04070_));
 sky130_fd_sc_hd__clkbuf_2 _14399_ (.A(instr_retirq),
    .X(_11568_));
 sky130_vsdinv _14400_ (.A(\cpu_state[2] ),
    .Y(_11569_));
 sky130_fd_sc_hd__buf_2 _14401_ (.A(_11569_),
    .X(_11570_));
 sky130_fd_sc_hd__buf_1 _14402_ (.A(_11570_),
    .X(_11571_));
 sky130_fd_sc_hd__clkbuf_2 _14403_ (.A(_11571_),
    .X(_11572_));
 sky130_fd_sc_hd__o21ba_1 _14404_ (.A1(_11568_),
    .A2(_11572_),
    .B1_N(_00331_),
    .X(_11573_));
 sky130_vsdinv _14405_ (.A(_11573_),
    .Y(_11574_));
 sky130_fd_sc_hd__buf_1 _14406_ (.A(latched_branch),
    .X(_11575_));
 sky130_fd_sc_hd__buf_1 _14407_ (.A(_11575_),
    .X(_11576_));
 sky130_fd_sc_hd__o221a_1 _14408_ (.A1(_14319_),
    .A2(_11574_),
    .B1(_11576_),
    .B2(_11573_),
    .C1(_11566_),
    .X(_04069_));
 sky130_vsdinv _14409_ (.A(net101),
    .Y(_11577_));
 sky130_fd_sc_hd__clkbuf_2 _14410_ (.A(_11577_),
    .X(_11578_));
 sky130_fd_sc_hd__buf_1 _14411_ (.A(_11578_),
    .X(_11579_));
 sky130_fd_sc_hd__buf_1 _14412_ (.A(_11579_),
    .X(_11580_));
 sky130_fd_sc_hd__clkbuf_2 _14413_ (.A(_11580_),
    .X(_11581_));
 sky130_fd_sc_hd__buf_1 _14414_ (.A(net408),
    .X(_11582_));
 sky130_fd_sc_hd__or2_1 _14415_ (.A(_11581_),
    .B(_11582_),
    .X(_11583_));
 sky130_vsdinv _14416_ (.A(_11583_),
    .Y(_11584_));
 sky130_fd_sc_hd__buf_1 _14417_ (.A(_11579_),
    .X(_11585_));
 sky130_fd_sc_hd__clkbuf_2 _14418_ (.A(_11585_),
    .X(_11586_));
 sky130_fd_sc_hd__clkbuf_2 _14419_ (.A(_11586_),
    .X(_11587_));
 sky130_fd_sc_hd__buf_1 _14420_ (.A(mem_do_wdata),
    .X(_11588_));
 sky130_fd_sc_hd__or2_2 _14421_ (.A(_11551_),
    .B(mem_do_prefetch),
    .X(_11589_));
 sky130_fd_sc_hd__or2_1 _14422_ (.A(_11557_),
    .B(_11589_),
    .X(_11590_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _14423_ (.A(_11553_),
    .X(_11591_));
 sky130_vsdinv _14424_ (.A(_11582_),
    .Y(_11592_));
 sky130_fd_sc_hd__a221o_1 _14425_ (.A1(\mem_state[0] ),
    .A2(_11551_),
    .B1(_11549_),
    .B2(_11547_),
    .C1(_11548_),
    .X(_11593_));
 sky130_fd_sc_hd__o311a_1 _14426_ (.A1(_11588_),
    .A2(_11590_),
    .A3(_11591_),
    .B1(_11592_),
    .C1(_11593_),
    .X(_11594_));
 sky130_fd_sc_hd__o21ai_1 _14427_ (.A1(_11587_),
    .A2(_11594_),
    .B1(_00300_),
    .Y(_11595_));
 sky130_vsdinv _14428_ (.A(_11595_),
    .Y(_11596_));
 sky130_fd_sc_hd__a32o_1 _14429_ (.A1(_14284_),
    .A2(_11584_),
    .A3(_11596_),
    .B1(\mem_state[1] ),
    .B2(_11595_),
    .X(_04068_));
 sky130_fd_sc_hd__a32o_1 _14430_ (.A1(_14283_),
    .A2(_11584_),
    .A3(_11596_),
    .B1(\mem_state[0] ),
    .B2(_11595_),
    .X(_04067_));
 sky130_vsdinv _14431_ (.A(_11551_),
    .Y(_11597_));
 sky130_fd_sc_hd__or2_2 _14432_ (.A(_11597_),
    .B(_11555_),
    .X(_11598_));
 sky130_fd_sc_hd__buf_1 _14433_ (.A(_11598_),
    .X(_11599_));
 sky130_vsdinv _14434_ (.A(_11599_),
    .Y(_11600_));
 sky130_fd_sc_hd__buf_1 _14435_ (.A(_11600_),
    .X(_11601_));
 sky130_fd_sc_hd__clkbuf_2 _14436_ (.A(_11601_),
    .X(_14286_));
 sky130_fd_sc_hd__buf_1 _14437_ (.A(_11599_),
    .X(_11602_));
 sky130_fd_sc_hd__clkbuf_2 _14438_ (.A(_11602_),
    .X(_00337_));
 sky130_vsdinv _14439_ (.A(_00327_),
    .Y(_11603_));
 sky130_fd_sc_hd__or3_1 _14440_ (.A(\mem_rdata_latched[28] ),
    .B(_11603_),
    .C(_00330_),
    .X(_11604_));
 sky130_vsdinv _14441_ (.A(_00325_),
    .Y(_11605_));
 sky130_vsdinv _14442_ (.A(_00324_),
    .Y(_11606_));
 sky130_fd_sc_hd__or3_4 _14443_ (.A(_11605_),
    .B(_11606_),
    .C(_00326_),
    .X(_11607_));
 sky130_fd_sc_hd__or4_4 _14444_ (.A(_00329_),
    .B(_00328_),
    .C(_11604_),
    .D(_11607_),
    .X(_11608_));
 sky130_fd_sc_hd__or2_1 _14445_ (.A(\mem_rdata_latched[27] ),
    .B(_11608_),
    .X(_11609_));
 sky130_fd_sc_hd__or3_1 _14446_ (.A(\mem_rdata_latched[31] ),
    .B(\mem_rdata_latched[30] ),
    .C(\mem_rdata_latched[29] ),
    .X(_11610_));
 sky130_fd_sc_hd__or3_1 _14447_ (.A(\mem_rdata_latched[26] ),
    .B(\mem_rdata_latched[25] ),
    .C(_11610_),
    .X(_11611_));
 sky130_fd_sc_hd__o21ba_1 _14448_ (.A1(_11609_),
    .A2(_11611_),
    .B1_N(\mem_rdata_latched[19] ),
    .X(_11612_));
 sky130_fd_sc_hd__or4b_4 _14449_ (.A(_11609_),
    .B(\mem_rdata_latched[25] ),
    .C(_11610_),
    .D_N(\mem_rdata_latched[26] ),
    .X(_11613_));
 sky130_vsdinv _14450_ (.A(\decoded_rs1[4] ),
    .Y(_00366_));
 sky130_fd_sc_hd__clkbuf_2 _14451_ (.A(_11600_),
    .X(_11614_));
 sky130_fd_sc_hd__o22a_1 _14452_ (.A1(_11602_),
    .A2(_11613_),
    .B1(_00366_),
    .B2(_11614_),
    .X(_11615_));
 sky130_fd_sc_hd__o21ai_1 _14453_ (.A1(_00337_),
    .A2(_11612_),
    .B1(_11615_),
    .Y(_04066_));
 sky130_vsdinv _14454_ (.A(\cpu_state[1] ),
    .Y(_11616_));
 sky130_fd_sc_hd__buf_1 _14455_ (.A(decoder_trigger),
    .X(_11617_));
 sky130_vsdinv _14456_ (.A(_11617_),
    .Y(_11618_));
 sky130_vsdinv _14457_ (.A(\irq_mask[1] ),
    .Y(_11619_));
 sky130_vsdinv _14458_ (.A(\irq_mask[2] ),
    .Y(_11620_));
 sky130_vsdinv _14459_ (.A(\irq_pending[0] ),
    .Y(_11621_));
 sky130_vsdinv _14460_ (.A(\irq_pending[3] ),
    .Y(_11622_));
 sky130_fd_sc_hd__o22ai_1 _14461_ (.A1(\irq_mask[0] ),
    .A2(_11621_),
    .B1(\irq_mask[3] ),
    .B2(_11622_),
    .Y(_11623_));
 sky130_fd_sc_hd__a221o_1 _14462_ (.A1(_11619_),
    .A2(\irq_pending[1] ),
    .B1(_11620_),
    .B2(\irq_pending[2] ),
    .C1(_11623_),
    .X(_11624_));
 sky130_vsdinv _14463_ (.A(\irq_pending[17] ),
    .Y(_11625_));
 sky130_vsdinv _14464_ (.A(\irq_pending[19] ),
    .Y(_11626_));
 sky130_vsdinv _14465_ (.A(\irq_pending[16] ),
    .Y(_11627_));
 sky130_vsdinv _14466_ (.A(\irq_pending[18] ),
    .Y(_11628_));
 sky130_fd_sc_hd__o22a_1 _14467_ (.A1(\irq_mask[16] ),
    .A2(_11627_),
    .B1(\irq_mask[18] ),
    .B2(_11628_),
    .X(_11629_));
 sky130_fd_sc_hd__o221ai_4 _14468_ (.A1(\irq_mask[17] ),
    .A2(_11625_),
    .B1(\irq_mask[19] ),
    .B2(_11626_),
    .C1(_11629_),
    .Y(_11630_));
 sky130_vsdinv _14469_ (.A(\irq_mask[24] ),
    .Y(_11631_));
 sky130_vsdinv _14470_ (.A(\irq_mask[26] ),
    .Y(_11632_));
 sky130_vsdinv _14471_ (.A(\irq_pending[25] ),
    .Y(_11633_));
 sky130_vsdinv _14472_ (.A(\irq_pending[27] ),
    .Y(_11634_));
 sky130_fd_sc_hd__o22ai_1 _14473_ (.A1(\irq_mask[25] ),
    .A2(_11633_),
    .B1(\irq_mask[27] ),
    .B2(_11634_),
    .Y(_11635_));
 sky130_fd_sc_hd__a221o_1 _14474_ (.A1(_11631_),
    .A2(\irq_pending[24] ),
    .B1(_11632_),
    .B2(\irq_pending[26] ),
    .C1(_11635_),
    .X(_11636_));
 sky130_vsdinv _14475_ (.A(\irq_mask[5] ),
    .Y(_11637_));
 sky130_vsdinv _14476_ (.A(\irq_mask[7] ),
    .Y(_11638_));
 sky130_vsdinv _14477_ (.A(\irq_pending[4] ),
    .Y(_11639_));
 sky130_vsdinv _14478_ (.A(\irq_pending[6] ),
    .Y(_11640_));
 sky130_fd_sc_hd__o22ai_1 _14479_ (.A1(\irq_mask[4] ),
    .A2(_11639_),
    .B1(\irq_mask[6] ),
    .B2(_11640_),
    .Y(_11641_));
 sky130_fd_sc_hd__a221o_1 _14480_ (.A1(_11637_),
    .A2(\irq_pending[5] ),
    .B1(_11638_),
    .B2(\irq_pending[7] ),
    .C1(_11641_),
    .X(_11642_));
 sky130_fd_sc_hd__or4_4 _14481_ (.A(_11624_),
    .B(_11630_),
    .C(_11636_),
    .D(_11642_),
    .X(_11643_));
 sky130_vsdinv _14482_ (.A(\irq_mask[13] ),
    .Y(_11644_));
 sky130_vsdinv _14483_ (.A(\irq_mask[15] ),
    .Y(_11645_));
 sky130_vsdinv _14484_ (.A(\irq_pending[12] ),
    .Y(_11646_));
 sky130_vsdinv _14485_ (.A(\irq_pending[14] ),
    .Y(_11647_));
 sky130_fd_sc_hd__o22ai_1 _14486_ (.A1(\irq_mask[12] ),
    .A2(_11646_),
    .B1(\irq_mask[14] ),
    .B2(_11647_),
    .Y(_11648_));
 sky130_fd_sc_hd__a221o_1 _14487_ (.A1(_11644_),
    .A2(\irq_pending[13] ),
    .B1(_11645_),
    .B2(\irq_pending[15] ),
    .C1(_11648_),
    .X(_11649_));
 sky130_vsdinv _14488_ (.A(\irq_mask[28] ),
    .Y(_11650_));
 sky130_vsdinv _14489_ (.A(\irq_mask[30] ),
    .Y(_11651_));
 sky130_vsdinv _14490_ (.A(\irq_pending[29] ),
    .Y(_11652_));
 sky130_vsdinv _14491_ (.A(\irq_pending[31] ),
    .Y(_11653_));
 sky130_fd_sc_hd__o22ai_1 _14492_ (.A1(\irq_mask[29] ),
    .A2(_11652_),
    .B1(\irq_mask[31] ),
    .B2(_11653_),
    .Y(_11654_));
 sky130_fd_sc_hd__a221o_1 _14493_ (.A1(_11650_),
    .A2(\irq_pending[28] ),
    .B1(_11651_),
    .B2(\irq_pending[30] ),
    .C1(_11654_),
    .X(_11655_));
 sky130_vsdinv _14494_ (.A(\irq_mask[9] ),
    .Y(_11656_));
 sky130_vsdinv _14495_ (.A(\irq_mask[11] ),
    .Y(_11657_));
 sky130_vsdinv _14496_ (.A(\irq_pending[8] ),
    .Y(_11658_));
 sky130_vsdinv _14497_ (.A(\irq_pending[10] ),
    .Y(_11659_));
 sky130_fd_sc_hd__o22ai_1 _14498_ (.A1(\irq_mask[8] ),
    .A2(_11658_),
    .B1(\irq_mask[10] ),
    .B2(_11659_),
    .Y(_11660_));
 sky130_fd_sc_hd__a221o_1 _14499_ (.A1(_11656_),
    .A2(\irq_pending[9] ),
    .B1(_11657_),
    .B2(\irq_pending[11] ),
    .C1(_11660_),
    .X(_11661_));
 sky130_vsdinv _14500_ (.A(\irq_mask[20] ),
    .Y(_11662_));
 sky130_vsdinv _14501_ (.A(\irq_mask[22] ),
    .Y(_11663_));
 sky130_vsdinv _14502_ (.A(\irq_pending[21] ),
    .Y(_11664_));
 sky130_vsdinv _14503_ (.A(\irq_pending[23] ),
    .Y(_11665_));
 sky130_fd_sc_hd__o22ai_1 _14504_ (.A1(\irq_mask[21] ),
    .A2(_11664_),
    .B1(\irq_mask[23] ),
    .B2(_11665_),
    .Y(_11666_));
 sky130_fd_sc_hd__a221o_1 _14505_ (.A1(_11662_),
    .A2(\irq_pending[20] ),
    .B1(_11663_),
    .B2(\irq_pending[22] ),
    .C1(_11666_),
    .X(_11667_));
 sky130_fd_sc_hd__or4_4 _14506_ (.A(_11649_),
    .B(_11655_),
    .C(_11661_),
    .D(_11667_),
    .X(_11668_));
 sky130_vsdinv _14507_ (.A(irq_active),
    .Y(_11669_));
 sky130_vsdinv _14508_ (.A(irq_delay),
    .Y(_11670_));
 sky130_fd_sc_hd__o2111a_1 _14509_ (.A1(_11643_),
    .A2(_11668_),
    .B1(_11669_),
    .C1(_11670_),
    .D1(decoder_trigger),
    .X(_11671_));
 sky130_fd_sc_hd__or3_4 _14510_ (.A(\irq_state[1] ),
    .B(\irq_state[0] ),
    .C(_11671_),
    .X(_11672_));
 sky130_fd_sc_hd__o21ai_2 _14511_ (.A1(decoder_trigger),
    .A2(do_waitirq),
    .B1(instr_waitirq),
    .Y(_11673_));
 sky130_vsdinv _14512_ (.A(_11673_),
    .Y(_00309_));
 sky130_fd_sc_hd__or2_1 _14513_ (.A(_11672_),
    .B(_00309_),
    .X(_11674_));
 sky130_fd_sc_hd__or3_4 _14514_ (.A(_11616_),
    .B(_11618_),
    .C(_11674_),
    .X(_11675_));
 sky130_vsdinv _14515_ (.A(_11675_),
    .Y(_11676_));
 sky130_fd_sc_hd__buf_1 _14516_ (.A(irq_active),
    .X(_11677_));
 sky130_fd_sc_hd__clkbuf_2 _14517_ (.A(_11543_),
    .X(_11678_));
 sky130_fd_sc_hd__clkbuf_2 _14518_ (.A(_11678_),
    .X(_11679_));
 sky130_fd_sc_hd__buf_2 _14519_ (.A(_11679_),
    .X(_11680_));
 sky130_fd_sc_hd__buf_2 _14520_ (.A(_11680_),
    .X(_11681_));
 sky130_fd_sc_hd__o221a_1 _14521_ (.A1(irq_delay),
    .A2(_11676_),
    .B1(_11677_),
    .B2(_11675_),
    .C1(_11681_),
    .X(_04065_));
 sky130_fd_sc_hd__buf_1 _14522_ (.A(net330),
    .X(_11682_));
 sky130_vsdinv _14523_ (.A(_11682_),
    .Y(_11683_));
 sky130_fd_sc_hd__buf_2 _14524_ (.A(_11683_),
    .X(_11684_));
 sky130_vsdinv _14525_ (.A(net370),
    .Y(_11685_));
 sky130_fd_sc_hd__or2_4 _14526_ (.A(_11577_),
    .B(_11685_),
    .X(_11686_));
 sky130_fd_sc_hd__or4_4 _14527_ (.A(net298),
    .B(net297),
    .C(net295),
    .D(net294),
    .X(_11687_));
 sky130_fd_sc_hd__or4b_4 _14528_ (.A(net293),
    .B(net292),
    .C(net279),
    .D_N(net291),
    .X(_11688_));
 sky130_fd_sc_hd__or2b_1 _14529_ (.A(net296),
    .B_N(net285),
    .X(_11689_));
 sky130_fd_sc_hd__or4bb_4 _14530_ (.A(net302),
    .B(net299),
    .C_N(net300),
    .D_N(net301),
    .X(_11690_));
 sky130_fd_sc_hd__or4b_4 _14531_ (.A(_11688_),
    .B(_11689_),
    .C(_11690_),
    .D_N(net274),
    .X(_11691_));
 sky130_fd_sc_hd__or3_4 _14532_ (.A(_11686_),
    .B(_11687_),
    .C(_11691_),
    .X(_11692_));
 sky130_fd_sc_hd__or3_4 _14533_ (.A(\pcpi_mul.active[0] ),
    .B(\pcpi_mul.active[1] ),
    .C(_11692_),
    .X(_11693_));
 sky130_fd_sc_hd__buf_1 _14534_ (.A(_11693_),
    .X(_11694_));
 sky130_vsdinv _14535_ (.A(net278),
    .Y(_11695_));
 sky130_fd_sc_hd__or2b_1 _14536_ (.A(_11692_),
    .B_N(net277),
    .X(_11696_));
 sky130_vsdinv _14537_ (.A(_11696_),
    .Y(_11697_));
 sky130_fd_sc_hd__nor3_2 _14538_ (.A(_11695_),
    .B(net277),
    .C(_11692_),
    .Y(_11698_));
 sky130_fd_sc_hd__a21oi_1 _14539_ (.A1(_11695_),
    .A2(_11697_),
    .B1(_11698_),
    .Y(_11699_));
 sky130_vsdinv _14540_ (.A(\pcpi_mul.rs1[32] ),
    .Y(_11700_));
 sky130_fd_sc_hd__buf_1 _14541_ (.A(_11700_),
    .X(_11701_));
 sky130_fd_sc_hd__buf_1 _14542_ (.A(_11701_),
    .X(_11702_));
 sky130_fd_sc_hd__clkbuf_2 _14543_ (.A(_11702_),
    .X(_11703_));
 sky130_fd_sc_hd__clkbuf_2 _14544_ (.A(_11703_),
    .X(_11704_));
 sky130_fd_sc_hd__clkbuf_2 _14545_ (.A(_11704_),
    .X(_11705_));
 sky130_fd_sc_hd__buf_1 _14546_ (.A(_11705_),
    .X(_11706_));
 sky130_fd_sc_hd__clkbuf_2 _14547_ (.A(_11706_),
    .X(_11707_));
 sky130_vsdinv _14548_ (.A(_11693_),
    .Y(_11708_));
 sky130_fd_sc_hd__clkbuf_4 _14549_ (.A(_11708_),
    .X(_11709_));
 sky130_fd_sc_hd__buf_1 _14550_ (.A(_11709_),
    .X(_11710_));
 sky130_fd_sc_hd__o32a_1 _14551_ (.A1(_11684_),
    .A2(_11694_),
    .A3(_11699_),
    .B1(_11707_),
    .B2(_11710_),
    .X(_11711_));
 sky130_vsdinv _14552_ (.A(_11711_),
    .Y(_04064_));
 sky130_fd_sc_hd__buf_2 _14553_ (.A(net362),
    .X(_11712_));
 sky130_vsdinv _14554_ (.A(_11712_),
    .Y(_11713_));
 sky130_fd_sc_hd__buf_2 _14555_ (.A(_11713_),
    .X(_11714_));
 sky130_fd_sc_hd__or2_1 _14556_ (.A(net278),
    .B(_11696_),
    .X(_11715_));
 sky130_vsdinv _14557_ (.A(\pcpi_mul.rs2[32] ),
    .Y(_11716_));
 sky130_fd_sc_hd__buf_1 _14558_ (.A(_11716_),
    .X(_11717_));
 sky130_fd_sc_hd__buf_2 _14559_ (.A(_11717_),
    .X(_11718_));
 sky130_fd_sc_hd__clkbuf_2 _14560_ (.A(_11718_),
    .X(_11719_));
 sky130_fd_sc_hd__buf_1 _14561_ (.A(_11719_),
    .X(_11720_));
 sky130_fd_sc_hd__buf_1 _14562_ (.A(_11720_),
    .X(_11721_));
 sky130_fd_sc_hd__clkbuf_2 _14563_ (.A(_11721_),
    .X(_11722_));
 sky130_fd_sc_hd__buf_2 _14564_ (.A(_11722_),
    .X(_11723_));
 sky130_fd_sc_hd__o32a_1 _14565_ (.A1(_11714_),
    .A2(_11694_),
    .A3(_11715_),
    .B1(_11723_),
    .B2(_11710_),
    .X(_11724_));
 sky130_vsdinv _14566_ (.A(_11724_),
    .Y(_04063_));
 sky130_fd_sc_hd__clkbuf_2 _14567_ (.A(\cpu_state[4] ),
    .X(_11725_));
 sky130_fd_sc_hd__buf_2 _14568_ (.A(_11725_),
    .X(_11726_));
 sky130_vsdinv _14569_ (.A(_00333_),
    .Y(_11727_));
 sky130_vsdinv _14570_ (.A(is_beq_bne_blt_bge_bltu_bgeu),
    .Y(_11728_));
 sky130_fd_sc_hd__buf_1 _14571_ (.A(_11728_),
    .X(_11729_));
 sky130_fd_sc_hd__buf_1 _14572_ (.A(alu_wait),
    .X(_11730_));
 sky130_fd_sc_hd__o21a_1 _14573_ (.A1(_11729_),
    .A2(_11730_),
    .B1(_00333_),
    .X(_11731_));
 sky130_fd_sc_hd__o221a_1 _14574_ (.A1(_11726_),
    .A2(_11727_),
    .B1(latched_stalu),
    .B2(_11731_),
    .C1(_11681_),
    .X(_04062_));
 sky130_vsdinv _14575_ (.A(\cpu_state[4] ),
    .Y(_11732_));
 sky130_fd_sc_hd__buf_1 _14576_ (.A(_11732_),
    .X(_11733_));
 sky130_fd_sc_hd__clkbuf_2 _14577_ (.A(_11733_),
    .X(_11734_));
 sky130_fd_sc_hd__inv_2 _14578_ (.A(alu_wait),
    .Y(_00302_));
 sky130_fd_sc_hd__buf_1 _14579_ (.A(\cpu_state[2] ),
    .X(_11735_));
 sky130_fd_sc_hd__or3_4 _14580_ (.A(_11735_),
    .B(\cpu_state[3] ),
    .C(\cpu_state[1] ),
    .X(_11736_));
 sky130_fd_sc_hd__or2_1 _14581_ (.A(_11725_),
    .B(\cpu_state[6] ),
    .X(_11737_));
 sky130_fd_sc_hd__or2_1 _14582_ (.A(_11736_),
    .B(_11737_),
    .X(_11738_));
 sky130_fd_sc_hd__clkbuf_2 _14583_ (.A(_11735_),
    .X(_11739_));
 sky130_vsdinv _14584_ (.A(instr_rdcycle),
    .Y(_11740_));
 sky130_vsdinv _14585_ (.A(instr_rdinstrh),
    .Y(_11741_));
 sky130_vsdinv _14586_ (.A(instr_rdinstr),
    .Y(_11742_));
 sky130_vsdinv _14587_ (.A(instr_rdcycleh),
    .Y(_11743_));
 sky130_fd_sc_hd__and3_1 _14588_ (.A(_11741_),
    .B(_11742_),
    .C(_11743_),
    .X(_11744_));
 sky130_fd_sc_hd__buf_8 _14589_ (.A(_11744_),
    .X(_01714_));
 sky130_fd_sc_hd__or3_4 _14590_ (.A(instr_setq),
    .B(instr_getq),
    .C(instr_retirq),
    .X(_11745_));
 sky130_fd_sc_hd__nor3_4 _14591_ (.A(instr_maskirq),
    .B(_11745_),
    .C(instr_timer),
    .Y(_01717_));
 sky130_fd_sc_hd__and3_1 _14592_ (.A(_11740_),
    .B(net426),
    .C(net430),
    .X(_11746_));
 sky130_fd_sc_hd__nand2_1 _14593_ (.A(_11739_),
    .B(_11746_),
    .Y(_11747_));
 sky130_vsdinv _14594_ (.A(\pcpi_mul.active[1] ),
    .Y(_11748_));
 sky130_fd_sc_hd__nand2_1 _14595_ (.A(_11740_),
    .B(net426),
    .Y(_11749_));
 sky130_fd_sc_hd__or4_4 _14596_ (.A(instr_and),
    .B(instr_or),
    .C(instr_xor),
    .D(instr_sltu),
    .X(_11750_));
 sky130_fd_sc_hd__or4_4 _14597_ (.A(instr_sltiu),
    .B(instr_slti),
    .C(instr_bgeu),
    .D(instr_bge),
    .X(_11751_));
 sky130_fd_sc_hd__or4_4 _14598_ (.A(instr_maskirq),
    .B(_11745_),
    .C(_11750_),
    .D(_11751_),
    .X(_11752_));
 sky130_fd_sc_hd__or4_4 _14599_ (.A(instr_lw),
    .B(instr_lh),
    .C(instr_lb),
    .D(instr_jalr),
    .X(_11753_));
 sky130_fd_sc_hd__or4_4 _14600_ (.A(instr_sh),
    .B(instr_sb),
    .C(instr_lhu),
    .D(instr_lbu),
    .X(_11754_));
 sky130_fd_sc_hd__or2_2 _14601_ (.A(instr_auipc),
    .B(instr_lui),
    .X(_11755_));
 sky130_fd_sc_hd__or2_2 _14602_ (.A(instr_jal),
    .B(_11755_),
    .X(_00005_));
 sky130_fd_sc_hd__or4_4 _14603_ (.A(instr_sra),
    .B(instr_srai),
    .C(instr_srl),
    .D(instr_srli),
    .X(_11756_));
 sky130_fd_sc_hd__or4_4 _14604_ (.A(_11753_),
    .B(_11754_),
    .C(_00005_),
    .D(_11756_),
    .X(_11757_));
 sky130_fd_sc_hd__or4_4 _14605_ (.A(instr_andi),
    .B(instr_ori),
    .C(instr_xori),
    .D(instr_addi),
    .X(_11758_));
 sky130_fd_sc_hd__or4_4 _14606_ (.A(instr_slt),
    .B(instr_sll),
    .C(instr_sub),
    .D(instr_add),
    .X(_11759_));
 sky130_fd_sc_hd__or4_4 _14607_ (.A(instr_timer),
    .B(instr_waitirq),
    .C(instr_slli),
    .D(instr_sw),
    .X(_11760_));
 sky130_fd_sc_hd__or4_4 _14608_ (.A(instr_bltu),
    .B(instr_blt),
    .C(instr_bne),
    .D(instr_beq),
    .X(_11761_));
 sky130_fd_sc_hd__or4_4 _14609_ (.A(_11758_),
    .B(_11759_),
    .C(_11760_),
    .D(_11761_),
    .X(_11762_));
 sky130_fd_sc_hd__or4_4 _14610_ (.A(_11749_),
    .B(_11752_),
    .C(_11757_),
    .D(_11762_),
    .X(_11763_));
 sky130_fd_sc_hd__o21ai_1 _14611_ (.A1(_11748_),
    .A2(_11763_),
    .B1(\cpu_state[3] ),
    .Y(_11764_));
 sky130_fd_sc_hd__o2111a_1 _14612_ (.A1(_11734_),
    .A2(_00302_),
    .B1(_11738_),
    .C1(_11747_),
    .D1(_11764_),
    .X(_11765_));
 sky130_vsdinv _14613_ (.A(_11765_),
    .Y(_11766_));
 sky130_fd_sc_hd__o221a_1 _14614_ (.A1(_14320_),
    .A2(_11766_),
    .B1(latched_store),
    .B2(_11765_),
    .C1(_11681_),
    .X(_04061_));
 sky130_fd_sc_hd__clkbuf_4 _14615_ (.A(_11581_),
    .X(_11767_));
 sky130_fd_sc_hd__buf_1 _14616_ (.A(_11767_),
    .X(_11768_));
 sky130_fd_sc_hd__buf_2 _14617_ (.A(_11768_),
    .X(_11769_));
 sky130_fd_sc_hd__buf_1 _14618_ (.A(\irq_state[1] ),
    .X(_11770_));
 sky130_fd_sc_hd__buf_1 _14619_ (.A(_11770_),
    .X(_11771_));
 sky130_fd_sc_hd__clkbuf_2 _14620_ (.A(_11616_),
    .X(_11772_));
 sky130_fd_sc_hd__clkbuf_2 _14621_ (.A(_11772_),
    .X(_11773_));
 sky130_fd_sc_hd__clkbuf_2 _14622_ (.A(_11773_),
    .X(_11774_));
 sky130_fd_sc_hd__buf_1 _14623_ (.A(\irq_state[0] ),
    .X(_11775_));
 sky130_vsdinv _14624_ (.A(_11775_),
    .Y(_11776_));
 sky130_fd_sc_hd__clkbuf_2 _14625_ (.A(_11776_),
    .X(_11777_));
 sky130_vsdinv _14626_ (.A(_11770_),
    .Y(_11778_));
 sky130_fd_sc_hd__clkbuf_2 _14627_ (.A(_11778_),
    .X(_11779_));
 sky130_fd_sc_hd__clkbuf_2 _14628_ (.A(_11779_),
    .X(_11780_));
 sky130_fd_sc_hd__clkbuf_2 _14629_ (.A(\cpu_state[1] ),
    .X(_11781_));
 sky130_fd_sc_hd__buf_2 _14630_ (.A(_11781_),
    .X(_11782_));
 sky130_fd_sc_hd__o32a_1 _14631_ (.A1(_11771_),
    .A2(_11774_),
    .A3(_11777_),
    .B1(_11780_),
    .B2(_11782_),
    .X(_11783_));
 sky130_fd_sc_hd__nor2_1 _14632_ (.A(_11769_),
    .B(_11783_),
    .Y(_04060_));
 sky130_fd_sc_hd__clkbuf_4 _14633_ (.A(_11775_),
    .X(_11784_));
 sky130_fd_sc_hd__clkbuf_2 _14634_ (.A(_11784_),
    .X(_11785_));
 sky130_fd_sc_hd__clkbuf_2 _14635_ (.A(_11782_),
    .X(_11786_));
 sky130_fd_sc_hd__buf_1 _14636_ (.A(_11543_),
    .X(_11787_));
 sky130_fd_sc_hd__buf_1 _14637_ (.A(_11787_),
    .X(_11788_));
 sky130_fd_sc_hd__clkbuf_4 _14638_ (.A(_11788_),
    .X(_11789_));
 sky130_fd_sc_hd__clkbuf_2 _14639_ (.A(_11773_),
    .X(_11790_));
 sky130_fd_sc_hd__clkbuf_2 _14640_ (.A(_11790_),
    .X(_11791_));
 sky130_fd_sc_hd__a31o_1 _14641_ (.A1(_11780_),
    .A2(_11777_),
    .A3(_11671_),
    .B1(_11791_),
    .X(_11792_));
 sky130_fd_sc_hd__o211a_1 _14642_ (.A1(_11785_),
    .A2(_11786_),
    .B1(_11789_),
    .C1(_11792_),
    .X(_04059_));
 sky130_vsdinv _14643_ (.A(_00356_),
    .Y(_11793_));
 sky130_fd_sc_hd__or2_1 _14644_ (.A(_11578_),
    .B(_11554_),
    .X(_11794_));
 sky130_fd_sc_hd__buf_1 _14645_ (.A(_11794_),
    .X(_11795_));
 sky130_vsdinv _14646_ (.A(_11795_),
    .Y(_11796_));
 sky130_vsdinv _14647_ (.A(is_lb_lh_lw_lbu_lhu),
    .Y(_11797_));
 sky130_vsdinv _14648_ (.A(_11763_),
    .Y(_11798_));
 sky130_fd_sc_hd__nor2_2 _14649_ (.A(_11797_),
    .B(_11798_),
    .Y(_11799_));
 sky130_vsdinv _14650_ (.A(is_sb_sh_sw),
    .Y(_11800_));
 sky130_fd_sc_hd__clkbuf_2 _14651_ (.A(_11800_),
    .X(_11801_));
 sky130_fd_sc_hd__clkbuf_2 _14652_ (.A(_11798_),
    .X(_00310_));
 sky130_fd_sc_hd__nor2_1 _14653_ (.A(_11801_),
    .B(_00310_),
    .Y(_11802_));
 sky130_fd_sc_hd__a22o_1 _14654_ (.A1(_11725_),
    .A2(_11730_),
    .B1(_11732_),
    .B2(_11736_),
    .X(_11803_));
 sky130_fd_sc_hd__o221a_1 _14655_ (.A1(_11571_),
    .A2(_11799_),
    .B1(_11764_),
    .B2(_11802_),
    .C1(_11803_),
    .X(_11804_));
 sky130_fd_sc_hd__or2_1 _14656_ (.A(_11795_),
    .B(_11804_),
    .X(_11805_));
 sky130_fd_sc_hd__or2_2 _14657_ (.A(\cpu_state[6] ),
    .B(\cpu_state[5] ),
    .X(_11806_));
 sky130_fd_sc_hd__or4_4 _14658_ (.A(_11729_),
    .B(_11730_),
    .C(_11586_),
    .D(_00343_),
    .X(_11807_));
 sky130_fd_sc_hd__nor4_2 _14659_ (.A(\cpu_state[0] ),
    .B(_11736_),
    .C(_11806_),
    .D(_11807_),
    .Y(_11808_));
 sky130_fd_sc_hd__nor2_1 _14660_ (.A(_11597_),
    .B(_11805_),
    .Y(_11809_));
 sky130_fd_sc_hd__a311o_1 _14661_ (.A1(_11793_),
    .A2(_11796_),
    .A3(_11805_),
    .B1(_11808_),
    .C1(_11809_),
    .X(_04058_));
 sky130_fd_sc_hd__or2_2 _14662_ (.A(instr_jal),
    .B(_11675_),
    .X(_11810_));
 sky130_vsdinv _14663_ (.A(_11810_),
    .Y(_11811_));
 sky130_fd_sc_hd__buf_1 _14664_ (.A(instr_jalr),
    .X(_11812_));
 sky130_fd_sc_hd__nor2_1 _14665_ (.A(_11568_),
    .B(_11812_),
    .Y(_11813_));
 sky130_fd_sc_hd__o221a_1 _14666_ (.A1(_11545_),
    .A2(_11811_),
    .B1(_11810_),
    .B2(_11813_),
    .C1(_11796_),
    .X(_04057_));
 sky130_fd_sc_hd__buf_2 _14667_ (.A(\irq_mask[31] ),
    .X(_11814_));
 sky130_vsdinv _14668_ (.A(instr_maskirq),
    .Y(_11815_));
 sky130_fd_sc_hd__or2_1 _14669_ (.A(_11815_),
    .B(_11570_),
    .X(_11816_));
 sky130_fd_sc_hd__clkbuf_2 _14670_ (.A(_11816_),
    .X(_11817_));
 sky130_fd_sc_hd__buf_1 _14671_ (.A(_11817_),
    .X(_11818_));
 sky130_fd_sc_hd__or3b_2 _14672_ (.A(net454),
    .B(_00360_),
    .C_N(net428),
    .X(_11819_));
 sky130_fd_sc_hd__or3_1 _14673_ (.A(net448),
    .B(net439),
    .C(_11819_),
    .X(_11820_));
 sky130_vsdinv _14674_ (.A(_11820_),
    .Y(_11821_));
 sky130_fd_sc_hd__buf_8 _14675_ (.A(_11821_),
    .X(_11822_));
 sky130_fd_sc_hd__clkbuf_8 _14676_ (.A(_11822_),
    .X(_11823_));
 sky130_fd_sc_hd__nor2_8 _14677_ (.A(_01207_),
    .B(_11823_),
    .Y(\cpuregs_rs1[31] ));
 sky130_vsdinv _14678_ (.A(_11816_),
    .Y(_11824_));
 sky130_fd_sc_hd__buf_1 _14679_ (.A(_11824_),
    .X(_11825_));
 sky130_fd_sc_hd__clkbuf_2 _14680_ (.A(_11825_),
    .X(_11826_));
 sky130_fd_sc_hd__buf_2 _14681_ (.A(_11586_),
    .X(_11827_));
 sky130_fd_sc_hd__buf_1 _14682_ (.A(_11827_),
    .X(_11828_));
 sky130_fd_sc_hd__a221o_1 _14683_ (.A1(_11814_),
    .A2(_11818_),
    .B1(\cpuregs_rs1[31] ),
    .B2(_11826_),
    .C1(_11828_),
    .X(_04056_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _14684_ (.A(_11824_),
    .X(_11829_));
 sky130_fd_sc_hd__buf_1 _14685_ (.A(_11829_),
    .X(_11830_));
 sky130_fd_sc_hd__buf_4 _14686_ (.A(_11821_),
    .X(_11831_));
 sky130_fd_sc_hd__clkbuf_8 _14687_ (.A(_11831_),
    .X(_11832_));
 sky130_fd_sc_hd__nor2_8 _14688_ (.A(_01180_),
    .B(_11832_),
    .Y(\cpuregs_rs1[30] ));
 sky130_fd_sc_hd__a221o_1 _14689_ (.A1(\irq_mask[30] ),
    .A2(_11818_),
    .B1(_11830_),
    .B2(\cpuregs_rs1[30] ),
    .C1(_11828_),
    .X(_04055_));
 sky130_fd_sc_hd__clkbuf_2 _14690_ (.A(\irq_mask[29] ),
    .X(_11833_));
 sky130_fd_sc_hd__nor2_8 _14691_ (.A(_01153_),
    .B(_11823_),
    .Y(\cpuregs_rs1[29] ));
 sky130_fd_sc_hd__a221o_1 _14692_ (.A1(_11833_),
    .A2(_11818_),
    .B1(_11830_),
    .B2(\cpuregs_rs1[29] ),
    .C1(_11828_),
    .X(_04054_));
 sky130_fd_sc_hd__nor2_8 _14693_ (.A(_01126_),
    .B(_11832_),
    .Y(\cpuregs_rs1[28] ));
 sky130_fd_sc_hd__a221o_1 _14694_ (.A1(\irq_mask[28] ),
    .A2(_11818_),
    .B1(_11830_),
    .B2(\cpuregs_rs1[28] ),
    .C1(_11828_),
    .X(_04053_));
 sky130_fd_sc_hd__clkbuf_2 _14695_ (.A(\irq_mask[27] ),
    .X(_11834_));
 sky130_fd_sc_hd__buf_1 _14696_ (.A(_11817_),
    .X(_11835_));
 sky130_fd_sc_hd__nor2_8 _14697_ (.A(_01099_),
    .B(_11823_),
    .Y(\cpuregs_rs1[27] ));
 sky130_fd_sc_hd__buf_1 _14698_ (.A(_11827_),
    .X(_11836_));
 sky130_fd_sc_hd__a221o_1 _14699_ (.A1(_11834_),
    .A2(_11835_),
    .B1(_11830_),
    .B2(\cpuregs_rs1[27] ),
    .C1(_11836_),
    .X(_04052_));
 sky130_fd_sc_hd__buf_1 _14700_ (.A(_11829_),
    .X(_11837_));
 sky130_fd_sc_hd__nor2_8 _14701_ (.A(_01072_),
    .B(_11832_),
    .Y(\cpuregs_rs1[26] ));
 sky130_fd_sc_hd__a221o_1 _14702_ (.A1(\irq_mask[26] ),
    .A2(_11835_),
    .B1(_11837_),
    .B2(\cpuregs_rs1[26] ),
    .C1(_11836_),
    .X(_04051_));
 sky130_fd_sc_hd__clkbuf_2 _14703_ (.A(\irq_mask[25] ),
    .X(_11838_));
 sky130_fd_sc_hd__nor2_8 _14704_ (.A(_01045_),
    .B(_11823_),
    .Y(\cpuregs_rs1[25] ));
 sky130_fd_sc_hd__a221o_1 _14705_ (.A1(_11838_),
    .A2(_11835_),
    .B1(_11837_),
    .B2(\cpuregs_rs1[25] ),
    .C1(_11836_),
    .X(_04050_));
 sky130_fd_sc_hd__nor2_8 _14706_ (.A(_01018_),
    .B(_11832_),
    .Y(\cpuregs_rs1[24] ));
 sky130_fd_sc_hd__a221o_1 _14707_ (.A1(\irq_mask[24] ),
    .A2(_11835_),
    .B1(_11837_),
    .B2(\cpuregs_rs1[24] ),
    .C1(_11836_),
    .X(_04049_));
 sky130_fd_sc_hd__clkbuf_2 _14708_ (.A(\irq_mask[23] ),
    .X(_11839_));
 sky130_fd_sc_hd__buf_1 _14709_ (.A(_11817_),
    .X(_11840_));
 sky130_fd_sc_hd__buf_8 _14710_ (.A(_11831_),
    .X(_11841_));
 sky130_fd_sc_hd__nor2_8 _14711_ (.A(_00991_),
    .B(_11841_),
    .Y(\cpuregs_rs1[23] ));
 sky130_fd_sc_hd__buf_1 _14712_ (.A(_11827_),
    .X(_11842_));
 sky130_fd_sc_hd__a221o_1 _14713_ (.A1(_11839_),
    .A2(_11840_),
    .B1(_11837_),
    .B2(\cpuregs_rs1[23] ),
    .C1(_11842_),
    .X(_04048_));
 sky130_fd_sc_hd__buf_1 _14714_ (.A(_11829_),
    .X(_11843_));
 sky130_fd_sc_hd__buf_2 _14715_ (.A(_11821_),
    .X(_11844_));
 sky130_fd_sc_hd__nor2_8 _14716_ (.A(_00964_),
    .B(net413),
    .Y(\cpuregs_rs1[22] ));
 sky130_fd_sc_hd__a221o_1 _14717_ (.A1(\irq_mask[22] ),
    .A2(_11840_),
    .B1(_11843_),
    .B2(\cpuregs_rs1[22] ),
    .C1(_11842_),
    .X(_04047_));
 sky130_fd_sc_hd__clkbuf_2 _14718_ (.A(\irq_mask[21] ),
    .X(_11845_));
 sky130_fd_sc_hd__nor2_8 _14719_ (.A(_00937_),
    .B(_11841_),
    .Y(\cpuregs_rs1[21] ));
 sky130_fd_sc_hd__a221o_1 _14720_ (.A1(_11845_),
    .A2(_11840_),
    .B1(_11843_),
    .B2(\cpuregs_rs1[21] ),
    .C1(_11842_),
    .X(_04046_));
 sky130_fd_sc_hd__nor2_8 _14721_ (.A(_00910_),
    .B(net413),
    .Y(\cpuregs_rs1[20] ));
 sky130_fd_sc_hd__a221o_1 _14722_ (.A1(\irq_mask[20] ),
    .A2(_11840_),
    .B1(_11843_),
    .B2(\cpuregs_rs1[20] ),
    .C1(_11842_),
    .X(_04045_));
 sky130_fd_sc_hd__buf_2 _14723_ (.A(\irq_mask[19] ),
    .X(_11846_));
 sky130_fd_sc_hd__buf_1 _14724_ (.A(_11817_),
    .X(_11847_));
 sky130_fd_sc_hd__nor2_8 _14725_ (.A(_00883_),
    .B(_11841_),
    .Y(\cpuregs_rs1[19] ));
 sky130_fd_sc_hd__clkbuf_2 _14726_ (.A(_11581_),
    .X(_11848_));
 sky130_fd_sc_hd__buf_2 _14727_ (.A(_11848_),
    .X(_11849_));
 sky130_fd_sc_hd__buf_1 _14728_ (.A(_11849_),
    .X(_11850_));
 sky130_fd_sc_hd__a221o_1 _14729_ (.A1(_11846_),
    .A2(_11847_),
    .B1(_11843_),
    .B2(\cpuregs_rs1[19] ),
    .C1(_11850_),
    .X(_04044_));
 sky130_fd_sc_hd__buf_1 _14730_ (.A(_11829_),
    .X(_11851_));
 sky130_fd_sc_hd__nor2_8 _14731_ (.A(_00856_),
    .B(net413),
    .Y(\cpuregs_rs1[18] ));
 sky130_fd_sc_hd__a221o_1 _14732_ (.A1(\irq_mask[18] ),
    .A2(_11847_),
    .B1(_11851_),
    .B2(\cpuregs_rs1[18] ),
    .C1(_11850_),
    .X(_04043_));
 sky130_fd_sc_hd__buf_2 _14733_ (.A(\irq_mask[17] ),
    .X(_11852_));
 sky130_fd_sc_hd__nor2_8 _14734_ (.A(_00829_),
    .B(_11841_),
    .Y(\cpuregs_rs1[17] ));
 sky130_fd_sc_hd__a221o_1 _14735_ (.A1(_11852_),
    .A2(_11847_),
    .B1(_11851_),
    .B2(\cpuregs_rs1[17] ),
    .C1(_11850_),
    .X(_04042_));
 sky130_fd_sc_hd__buf_2 _14736_ (.A(\irq_mask[16] ),
    .X(_11853_));
 sky130_fd_sc_hd__buf_8 _14737_ (.A(_11831_),
    .X(_11854_));
 sky130_fd_sc_hd__nor2_8 _14738_ (.A(_00802_),
    .B(_11854_),
    .Y(\cpuregs_rs1[16] ));
 sky130_fd_sc_hd__a221o_1 _14739_ (.A1(_11853_),
    .A2(_11847_),
    .B1(_11851_),
    .B2(\cpuregs_rs1[16] ),
    .C1(_11850_),
    .X(_04041_));
 sky130_fd_sc_hd__buf_1 _14740_ (.A(_11816_),
    .X(_11855_));
 sky130_fd_sc_hd__buf_1 _14741_ (.A(_11855_),
    .X(_11856_));
 sky130_fd_sc_hd__nor2_8 _14742_ (.A(_00775_),
    .B(_11844_),
    .Y(\cpuregs_rs1[15] ));
 sky130_fd_sc_hd__buf_1 _14743_ (.A(_11849_),
    .X(_11857_));
 sky130_fd_sc_hd__a221o_1 _14744_ (.A1(\irq_mask[15] ),
    .A2(_11856_),
    .B1(_11851_),
    .B2(\cpuregs_rs1[15] ),
    .C1(_11857_),
    .X(_04040_));
 sky130_fd_sc_hd__clkbuf_2 _14745_ (.A(\irq_mask[14] ),
    .X(_11858_));
 sky130_fd_sc_hd__buf_1 _14746_ (.A(_11825_),
    .X(_11859_));
 sky130_fd_sc_hd__nor2_8 _14747_ (.A(_00748_),
    .B(_11854_),
    .Y(\cpuregs_rs1[14] ));
 sky130_fd_sc_hd__a221o_1 _14748_ (.A1(_11858_),
    .A2(_11856_),
    .B1(_11859_),
    .B2(\cpuregs_rs1[14] ),
    .C1(_11857_),
    .X(_04039_));
 sky130_fd_sc_hd__clkbuf_8 _14749_ (.A(_11821_),
    .X(_11860_));
 sky130_fd_sc_hd__nor2_8 _14750_ (.A(_00721_),
    .B(_11860_),
    .Y(\cpuregs_rs1[13] ));
 sky130_fd_sc_hd__a221o_1 _14751_ (.A1(\irq_mask[13] ),
    .A2(_11856_),
    .B1(_11859_),
    .B2(\cpuregs_rs1[13] ),
    .C1(_11857_),
    .X(_04038_));
 sky130_fd_sc_hd__clkbuf_2 _14752_ (.A(\irq_mask[12] ),
    .X(_11861_));
 sky130_fd_sc_hd__nor2_8 _14753_ (.A(_00694_),
    .B(_11854_),
    .Y(\cpuregs_rs1[12] ));
 sky130_fd_sc_hd__a221o_1 _14754_ (.A1(_11861_),
    .A2(_11856_),
    .B1(_11859_),
    .B2(\cpuregs_rs1[12] ),
    .C1(_11857_),
    .X(_04037_));
 sky130_fd_sc_hd__buf_1 _14755_ (.A(_11855_),
    .X(_11862_));
 sky130_fd_sc_hd__nor2_8 _14756_ (.A(_00667_),
    .B(_11860_),
    .Y(\cpuregs_rs1[11] ));
 sky130_fd_sc_hd__buf_1 _14757_ (.A(_11849_),
    .X(_11863_));
 sky130_fd_sc_hd__a221o_1 _14758_ (.A1(\irq_mask[11] ),
    .A2(_11862_),
    .B1(_11859_),
    .B2(\cpuregs_rs1[11] ),
    .C1(_11863_),
    .X(_04036_));
 sky130_fd_sc_hd__clkbuf_2 _14759_ (.A(\irq_mask[10] ),
    .X(_11864_));
 sky130_fd_sc_hd__buf_1 _14760_ (.A(_11825_),
    .X(_11865_));
 sky130_fd_sc_hd__nor2_8 _14761_ (.A(_00640_),
    .B(_11854_),
    .Y(\cpuregs_rs1[10] ));
 sky130_fd_sc_hd__a221o_1 _14762_ (.A1(_11864_),
    .A2(_11862_),
    .B1(_11865_),
    .B2(\cpuregs_rs1[10] ),
    .C1(_11863_),
    .X(_04035_));
 sky130_fd_sc_hd__nor2_8 _14763_ (.A(_00613_),
    .B(_11860_),
    .Y(\cpuregs_rs1[9] ));
 sky130_fd_sc_hd__a221o_1 _14764_ (.A1(\irq_mask[9] ),
    .A2(_11862_),
    .B1(_11865_),
    .B2(\cpuregs_rs1[9] ),
    .C1(_11863_),
    .X(_04034_));
 sky130_fd_sc_hd__buf_2 _14765_ (.A(\irq_mask[8] ),
    .X(_11866_));
 sky130_fd_sc_hd__clkbuf_8 _14766_ (.A(_11831_),
    .X(_11867_));
 sky130_fd_sc_hd__nor2_8 _14767_ (.A(_00586_),
    .B(_11867_),
    .Y(\cpuregs_rs1[8] ));
 sky130_fd_sc_hd__a221o_1 _14768_ (.A1(_11866_),
    .A2(_11862_),
    .B1(_11865_),
    .B2(\cpuregs_rs1[8] ),
    .C1(_11863_),
    .X(_04033_));
 sky130_fd_sc_hd__buf_1 _14769_ (.A(_11855_),
    .X(_11868_));
 sky130_fd_sc_hd__nor2_8 _14770_ (.A(_00559_),
    .B(_11860_),
    .Y(\cpuregs_rs1[7] ));
 sky130_fd_sc_hd__buf_1 _14771_ (.A(_11849_),
    .X(_11869_));
 sky130_fd_sc_hd__a221o_1 _14772_ (.A1(\irq_mask[7] ),
    .A2(_11868_),
    .B1(_11865_),
    .B2(\cpuregs_rs1[7] ),
    .C1(_11869_),
    .X(_04032_));
 sky130_fd_sc_hd__buf_2 _14773_ (.A(\irq_mask[6] ),
    .X(_11870_));
 sky130_fd_sc_hd__buf_1 _14774_ (.A(_11825_),
    .X(_11871_));
 sky130_fd_sc_hd__nor2_8 _14775_ (.A(_00532_),
    .B(_11867_),
    .Y(\cpuregs_rs1[6] ));
 sky130_fd_sc_hd__a221o_1 _14776_ (.A1(_11870_),
    .A2(_11868_),
    .B1(_11871_),
    .B2(\cpuregs_rs1[6] ),
    .C1(_11869_),
    .X(_04031_));
 sky130_fd_sc_hd__nor2_8 _14777_ (.A(_00505_),
    .B(_11822_),
    .Y(\cpuregs_rs1[5] ));
 sky130_fd_sc_hd__a221o_1 _14778_ (.A1(\irq_mask[5] ),
    .A2(_11868_),
    .B1(_11871_),
    .B2(\cpuregs_rs1[5] ),
    .C1(_11869_),
    .X(_04030_));
 sky130_fd_sc_hd__buf_2 _14779_ (.A(\irq_mask[4] ),
    .X(_11872_));
 sky130_fd_sc_hd__nor2_8 _14780_ (.A(_00478_),
    .B(_11867_),
    .Y(\cpuregs_rs1[4] ));
 sky130_fd_sc_hd__a221o_1 _14781_ (.A1(_11872_),
    .A2(_11868_),
    .B1(_11871_),
    .B2(\cpuregs_rs1[4] ),
    .C1(_11869_),
    .X(_04029_));
 sky130_fd_sc_hd__buf_2 _14782_ (.A(\irq_mask[3] ),
    .X(_11873_));
 sky130_fd_sc_hd__buf_1 _14783_ (.A(_11855_),
    .X(_11874_));
 sky130_fd_sc_hd__nor2_8 _14784_ (.A(_00451_),
    .B(_11867_),
    .Y(\cpuregs_rs1[3] ));
 sky130_fd_sc_hd__buf_1 _14785_ (.A(_11587_),
    .X(_11875_));
 sky130_fd_sc_hd__a221o_1 _14786_ (.A1(_11873_),
    .A2(_11874_),
    .B1(_11871_),
    .B2(\cpuregs_rs1[3] ),
    .C1(_11875_),
    .X(_04028_));
 sky130_fd_sc_hd__nor2_8 _14787_ (.A(_00424_),
    .B(_11822_),
    .Y(\cpuregs_rs1[2] ));
 sky130_fd_sc_hd__a221o_1 _14788_ (.A1(\irq_mask[2] ),
    .A2(_11874_),
    .B1(_11826_),
    .B2(\cpuregs_rs1[2] ),
    .C1(_11875_),
    .X(_04027_));
 sky130_fd_sc_hd__nor2_8 _14789_ (.A(_00397_),
    .B(_11822_),
    .Y(\cpuregs_rs1[1] ));
 sky130_fd_sc_hd__a221o_1 _14790_ (.A1(\irq_mask[1] ),
    .A2(_11874_),
    .B1(_11826_),
    .B2(\cpuregs_rs1[1] ),
    .C1(_11875_),
    .X(_04026_));
 sky130_fd_sc_hd__and2_1 _14791_ (.A(_00370_),
    .B(_11820_),
    .X(_11876_));
 sky130_fd_sc_hd__buf_4 _14792_ (.A(_11876_),
    .X(\cpuregs_rs1[0] ));
 sky130_fd_sc_hd__a221o_1 _14793_ (.A1(\irq_mask[0] ),
    .A2(_11874_),
    .B1(_11826_),
    .B2(\cpuregs_rs1[0] ),
    .C1(_11875_),
    .X(_04025_));
 sky130_vsdinv _14794_ (.A(_11588_),
    .Y(_11877_));
 sky130_fd_sc_hd__clkbuf_2 _14795_ (.A(_11877_),
    .X(_11878_));
 sky130_fd_sc_hd__clkbuf_2 _14796_ (.A(_11878_),
    .X(_00291_));
 sky130_vsdinv _14797_ (.A(_11589_),
    .Y(_11879_));
 sky130_fd_sc_hd__a311o_4 _14798_ (.A1(_11558_),
    .A2(_11879_),
    .A3(_11877_),
    .B1(_11591_),
    .C1(_11578_),
    .X(_00316_));
 sky130_fd_sc_hd__or2_4 _14799_ (.A(net408),
    .B(_00316_),
    .X(_11880_));
 sky130_vsdinv _14800_ (.A(_11880_),
    .Y(_11881_));
 sky130_fd_sc_hd__buf_4 _14801_ (.A(_11881_),
    .X(_11882_));
 sky130_fd_sc_hd__clkbuf_2 _14802_ (.A(_11880_),
    .X(_11883_));
 sky130_fd_sc_hd__buf_6 _14803_ (.A(_11883_),
    .X(_11884_));
 sky130_fd_sc_hd__a32o_1 _14804_ (.A1(_00291_),
    .A2(_11589_),
    .A3(_11882_),
    .B1(net166),
    .B2(_11884_),
    .X(_04024_));
 sky130_fd_sc_hd__buf_1 _14805_ (.A(_11599_),
    .X(_11885_));
 sky130_fd_sc_hd__buf_2 _14806_ (.A(_11885_),
    .X(_11886_));
 sky130_fd_sc_hd__clkbuf_2 _14807_ (.A(_00329_),
    .X(_11887_));
 sky130_vsdinv _14808_ (.A(_11887_),
    .Y(_11888_));
 sky130_fd_sc_hd__or3b_4 _14809_ (.A(_11888_),
    .B(_00328_),
    .C_N(_00330_),
    .X(_11889_));
 sky130_fd_sc_hd__nor3_4 _14810_ (.A(_00327_),
    .B(_11607_),
    .C(_11889_),
    .Y(_11890_));
 sky130_fd_sc_hd__buf_2 _14811_ (.A(is_beq_bne_blt_bge_bltu_bgeu),
    .X(_11891_));
 sky130_fd_sc_hd__o221a_1 _14812_ (.A1(_11886_),
    .A2(_11890_),
    .B1(_11891_),
    .B2(_11614_),
    .C1(_11681_),
    .X(_04023_));
 sky130_fd_sc_hd__buf_1 _14813_ (.A(_11600_),
    .X(_11892_));
 sky130_fd_sc_hd__buf_1 _14814_ (.A(_11892_),
    .X(_11893_));
 sky130_fd_sc_hd__clkbuf_2 _14815_ (.A(_11613_),
    .X(_11894_));
 sky130_fd_sc_hd__buf_1 _14816_ (.A(_11599_),
    .X(_11895_));
 sky130_fd_sc_hd__clkbuf_2 _14817_ (.A(_11895_),
    .X(_11896_));
 sky130_fd_sc_hd__a32o_1 _14818_ (.A1(\mem_rdata_latched[18] ),
    .A2(_11893_),
    .A3(_11894_),
    .B1(\decoded_rs1[3] ),
    .B2(_11896_),
    .X(_04022_));
 sky130_fd_sc_hd__a32o_1 _14819_ (.A1(\mem_rdata_latched[17] ),
    .A2(_11893_),
    .A3(_11894_),
    .B1(\decoded_rs1[2] ),
    .B2(_11896_),
    .X(_04021_));
 sky130_fd_sc_hd__clkbuf_2 _14820_ (.A(_11602_),
    .X(_11897_));
 sky130_fd_sc_hd__a32o_1 _14821_ (.A1(\mem_rdata_latched[16] ),
    .A2(_11893_),
    .A3(_11894_),
    .B1(\decoded_rs1[1] ),
    .B2(_11897_),
    .X(_04020_));
 sky130_fd_sc_hd__a32o_1 _14822_ (.A1(\mem_rdata_latched[15] ),
    .A2(_11893_),
    .A3(_11613_),
    .B1(\decoded_rs1[0] ),
    .B2(_11897_),
    .X(_04019_));
 sky130_fd_sc_hd__or2_2 _14823_ (.A(_11618_),
    .B(decoder_pseudo_trigger),
    .X(_11898_));
 sky130_fd_sc_hd__buf_1 _14824_ (.A(_11898_),
    .X(_11899_));
 sky130_fd_sc_hd__clkbuf_2 _14825_ (.A(_11899_),
    .X(_11900_));
 sky130_fd_sc_hd__buf_1 _14826_ (.A(_11900_),
    .X(_11901_));
 sky130_vsdinv _14827_ (.A(\mem_rdata_q[13] ),
    .Y(_11902_));
 sky130_fd_sc_hd__clkbuf_4 _14828_ (.A(_11902_),
    .X(_11903_));
 sky130_vsdinv _14829_ (.A(\mem_rdata_q[12] ),
    .Y(_11904_));
 sky130_fd_sc_hd__buf_2 _14830_ (.A(_11904_),
    .X(_11905_));
 sky130_vsdinv _14831_ (.A(\mem_rdata_q[14] ),
    .Y(_11906_));
 sky130_fd_sc_hd__clkbuf_4 _14832_ (.A(_11906_),
    .X(_00334_));
 sky130_fd_sc_hd__or3_4 _14833_ (.A(_11903_),
    .B(_11905_),
    .C(_00334_),
    .X(_11907_));
 sky130_vsdinv _14834_ (.A(is_alu_reg_reg),
    .Y(_11908_));
 sky130_fd_sc_hd__or4_4 _14835_ (.A(\mem_rdata_q[28] ),
    .B(\mem_rdata_q[26] ),
    .C(\mem_rdata_q[27] ),
    .D(\mem_rdata_q[25] ),
    .X(_11909_));
 sky130_fd_sc_hd__or4_4 _14836_ (.A(\mem_rdata_q[31] ),
    .B(\mem_rdata_q[30] ),
    .C(\mem_rdata_q[29] ),
    .D(_11909_),
    .X(_11910_));
 sky130_fd_sc_hd__or2_2 _14837_ (.A(_11898_),
    .B(_11910_),
    .X(_11911_));
 sky130_fd_sc_hd__or2_1 _14838_ (.A(_11908_),
    .B(_11911_),
    .X(_11912_));
 sky130_fd_sc_hd__o2bb2a_1 _14839_ (.A1_N(instr_and),
    .A2_N(_11901_),
    .B1(_11907_),
    .B2(_11912_),
    .X(_11913_));
 sky130_fd_sc_hd__nor2_1 _14840_ (.A(_11769_),
    .B(_11913_),
    .Y(_04018_));
 sky130_fd_sc_hd__buf_1 _14841_ (.A(_11912_),
    .X(_11914_));
 sky130_fd_sc_hd__buf_1 _14842_ (.A(\mem_rdata_q[12] ),
    .X(_11915_));
 sky130_fd_sc_hd__or3_4 _14843_ (.A(_11903_),
    .B(_11915_),
    .C(_11906_),
    .X(_11916_));
 sky130_fd_sc_hd__o2bb2a_1 _14844_ (.A1_N(instr_or),
    .A2_N(_11901_),
    .B1(_11914_),
    .B2(_11916_),
    .X(_11917_));
 sky130_fd_sc_hd__nor2_1 _14845_ (.A(_11769_),
    .B(_11917_),
    .Y(_04017_));
 sky130_fd_sc_hd__buf_1 _14846_ (.A(_11908_),
    .X(_11918_));
 sky130_fd_sc_hd__buf_1 _14847_ (.A(\mem_rdata_q[13] ),
    .X(_11919_));
 sky130_fd_sc_hd__or3_4 _14848_ (.A(_11919_),
    .B(_11904_),
    .C(_11906_),
    .X(_11920_));
 sky130_fd_sc_hd__buf_1 _14849_ (.A(\mem_rdata_q[29] ),
    .X(_11921_));
 sky130_fd_sc_hd__buf_1 _14850_ (.A(_11898_),
    .X(_11922_));
 sky130_fd_sc_hd__buf_1 _14851_ (.A(\mem_rdata_q[31] ),
    .X(_11923_));
 sky130_fd_sc_hd__clkbuf_2 _14852_ (.A(\mem_rdata_q[30] ),
    .X(_11924_));
 sky130_vsdinv _14853_ (.A(_11924_),
    .Y(_11925_));
 sky130_fd_sc_hd__clkbuf_2 _14854_ (.A(_11925_),
    .X(_11926_));
 sky130_fd_sc_hd__or3_1 _14855_ (.A(_11923_),
    .B(_11926_),
    .C(_11909_),
    .X(_11927_));
 sky130_fd_sc_hd__or3_4 _14856_ (.A(_11921_),
    .B(_11922_),
    .C(_11927_),
    .X(_11928_));
 sky130_vsdinv _14857_ (.A(instr_sra),
    .Y(_11929_));
 sky130_vsdinv _14858_ (.A(_11898_),
    .Y(_11930_));
 sky130_fd_sc_hd__buf_1 _14859_ (.A(_11930_),
    .X(_11931_));
 sky130_fd_sc_hd__buf_2 _14860_ (.A(_11931_),
    .X(_11932_));
 sky130_fd_sc_hd__o32a_1 _14861_ (.A1(_11918_),
    .A2(_11920_),
    .A3(_11928_),
    .B1(_11929_),
    .B2(_11932_),
    .X(_11933_));
 sky130_fd_sc_hd__nor2_1 _14862_ (.A(_11769_),
    .B(_11933_),
    .Y(_04016_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _14863_ (.A(_11768_),
    .X(_11934_));
 sky130_vsdinv _14864_ (.A(instr_srl),
    .Y(_11935_));
 sky130_fd_sc_hd__o32a_1 _14865_ (.A1(_11918_),
    .A2(_11920_),
    .A3(_11911_),
    .B1(_11935_),
    .B2(_11932_),
    .X(_11936_));
 sky130_fd_sc_hd__nor2_1 _14866_ (.A(_11934_),
    .B(_11936_),
    .Y(_04015_));
 sky130_fd_sc_hd__or3_4 _14867_ (.A(_11919_),
    .B(_11915_),
    .C(_11906_),
    .X(_11937_));
 sky130_fd_sc_hd__o2bb2a_1 _14868_ (.A1_N(instr_xor),
    .A2_N(_11901_),
    .B1(_11914_),
    .B2(_11937_),
    .X(_11938_));
 sky130_fd_sc_hd__nor2_1 _14869_ (.A(_11934_),
    .B(_11938_),
    .Y(_04014_));
 sky130_fd_sc_hd__buf_1 _14870_ (.A(\mem_rdata_q[14] ),
    .X(_11939_));
 sky130_fd_sc_hd__or3_4 _14871_ (.A(_11903_),
    .B(_11904_),
    .C(_11939_),
    .X(_11940_));
 sky130_fd_sc_hd__o2bb2a_1 _14872_ (.A1_N(instr_sltu),
    .A2_N(_11901_),
    .B1(_11914_),
    .B2(_11940_),
    .X(_11941_));
 sky130_fd_sc_hd__nor2_1 _14873_ (.A(_11934_),
    .B(_11941_),
    .Y(_04013_));
 sky130_fd_sc_hd__buf_1 _14874_ (.A(_11900_),
    .X(_11942_));
 sky130_fd_sc_hd__or3_4 _14875_ (.A(_11902_),
    .B(\mem_rdata_q[12] ),
    .C(\mem_rdata_q[14] ),
    .X(_11943_));
 sky130_fd_sc_hd__clkbuf_2 _14876_ (.A(_11943_),
    .X(_11944_));
 sky130_fd_sc_hd__o2bb2a_1 _14877_ (.A1_N(instr_slt),
    .A2_N(_11942_),
    .B1(_11914_),
    .B2(_11944_),
    .X(_11945_));
 sky130_fd_sc_hd__nor2_1 _14878_ (.A(_11934_),
    .B(_11945_),
    .Y(_04012_));
 sky130_fd_sc_hd__buf_1 _14879_ (.A(_11768_),
    .X(_11946_));
 sky130_fd_sc_hd__clkbuf_2 _14880_ (.A(_11919_),
    .X(_11947_));
 sky130_fd_sc_hd__or3_4 _14881_ (.A(_11947_),
    .B(_11905_),
    .C(_11939_),
    .X(_11948_));
 sky130_fd_sc_hd__o2bb2a_1 _14882_ (.A1_N(instr_sll),
    .A2_N(_11942_),
    .B1(_11912_),
    .B2(_11948_),
    .X(_11949_));
 sky130_fd_sc_hd__nor2_1 _14883_ (.A(_11946_),
    .B(_11949_),
    .Y(_04011_));
 sky130_fd_sc_hd__or3_4 _14884_ (.A(_11919_),
    .B(\mem_rdata_q[12] ),
    .C(\mem_rdata_q[14] ),
    .X(_11950_));
 sky130_fd_sc_hd__clkbuf_2 _14885_ (.A(_11950_),
    .X(_11951_));
 sky130_vsdinv _14886_ (.A(instr_sub),
    .Y(_11952_));
 sky130_fd_sc_hd__o32a_1 _14887_ (.A1(_11918_),
    .A2(_11951_),
    .A3(_11928_),
    .B1(_11952_),
    .B2(_11932_),
    .X(_11953_));
 sky130_fd_sc_hd__nor2_1 _14888_ (.A(_11946_),
    .B(_11953_),
    .Y(_04010_));
 sky130_vsdinv _14889_ (.A(instr_add),
    .Y(_11954_));
 sky130_fd_sc_hd__buf_1 _14890_ (.A(_11930_),
    .X(_11955_));
 sky130_fd_sc_hd__clkbuf_2 _14891_ (.A(_11955_),
    .X(_11956_));
 sky130_fd_sc_hd__buf_1 _14892_ (.A(_11956_),
    .X(_11957_));
 sky130_fd_sc_hd__o32a_1 _14893_ (.A1(_11908_),
    .A2(_11950_),
    .A3(_11911_),
    .B1(_11954_),
    .B2(_11957_),
    .X(_11958_));
 sky130_fd_sc_hd__nor2_1 _14894_ (.A(_11946_),
    .B(_11958_),
    .Y(_04009_));
 sky130_fd_sc_hd__buf_1 _14895_ (.A(is_alu_reg_imm),
    .X(_11959_));
 sky130_vsdinv _14896_ (.A(_11959_),
    .Y(_11960_));
 sky130_fd_sc_hd__clkbuf_2 _14897_ (.A(_11960_),
    .X(_11961_));
 sky130_fd_sc_hd__clkbuf_2 _14898_ (.A(_11899_),
    .X(_11962_));
 sky130_fd_sc_hd__buf_1 _14899_ (.A(_11962_),
    .X(_11963_));
 sky130_vsdinv _14900_ (.A(instr_andi),
    .Y(_11964_));
 sky130_fd_sc_hd__o32a_1 _14901_ (.A1(_11961_),
    .A2(_11963_),
    .A3(_11907_),
    .B1(_11964_),
    .B2(_11957_),
    .X(_11965_));
 sky130_fd_sc_hd__nor2_1 _14902_ (.A(_11946_),
    .B(_11965_),
    .Y(_04008_));
 sky130_fd_sc_hd__buf_1 _14903_ (.A(_11768_),
    .X(_11966_));
 sky130_vsdinv _14904_ (.A(instr_ori),
    .Y(_11967_));
 sky130_fd_sc_hd__o32a_1 _14905_ (.A1(_11961_),
    .A2(_11963_),
    .A3(_11916_),
    .B1(_11967_),
    .B2(_11957_),
    .X(_11968_));
 sky130_fd_sc_hd__nor2_1 _14906_ (.A(_11966_),
    .B(_11968_),
    .Y(_04007_));
 sky130_fd_sc_hd__buf_1 _14907_ (.A(_11960_),
    .X(_11969_));
 sky130_vsdinv _14908_ (.A(instr_xori),
    .Y(_11970_));
 sky130_fd_sc_hd__o32a_1 _14909_ (.A1(_11969_),
    .A2(_11963_),
    .A3(_11937_),
    .B1(_11970_),
    .B2(_11957_),
    .X(_11971_));
 sky130_fd_sc_hd__nor2_1 _14910_ (.A(_11966_),
    .B(_11971_),
    .Y(_04006_));
 sky130_fd_sc_hd__buf_1 _14911_ (.A(_11962_),
    .X(_11972_));
 sky130_vsdinv _14912_ (.A(instr_sltiu),
    .Y(_11973_));
 sky130_fd_sc_hd__buf_1 _14913_ (.A(_11956_),
    .X(_11974_));
 sky130_fd_sc_hd__o32a_1 _14914_ (.A1(_11969_),
    .A2(_11972_),
    .A3(_11940_),
    .B1(_11973_),
    .B2(_11974_),
    .X(_11975_));
 sky130_fd_sc_hd__nor2_1 _14915_ (.A(_11966_),
    .B(_11975_),
    .Y(_04005_));
 sky130_vsdinv _14916_ (.A(instr_slti),
    .Y(_11976_));
 sky130_fd_sc_hd__o32a_1 _14917_ (.A1(_11969_),
    .A2(_11972_),
    .A3(_11944_),
    .B1(_11976_),
    .B2(_11974_),
    .X(_11977_));
 sky130_fd_sc_hd__nor2_1 _14918_ (.A(_11966_),
    .B(_11977_),
    .Y(_04004_));
 sky130_fd_sc_hd__clkbuf_2 _14919_ (.A(_11767_),
    .X(_11978_));
 sky130_fd_sc_hd__buf_1 _14920_ (.A(_11978_),
    .X(_11979_));
 sky130_vsdinv _14921_ (.A(instr_addi),
    .Y(_11980_));
 sky130_fd_sc_hd__o32a_1 _14922_ (.A1(_11969_),
    .A2(_11972_),
    .A3(_11951_),
    .B1(_11980_),
    .B2(_11974_),
    .X(_11981_));
 sky130_fd_sc_hd__nor2_1 _14923_ (.A(_11979_),
    .B(_11981_),
    .Y(_04003_));
 sky130_fd_sc_hd__buf_2 _14924_ (.A(_11729_),
    .X(_11982_));
 sky130_vsdinv _14925_ (.A(instr_bgeu),
    .Y(_11983_));
 sky130_fd_sc_hd__o32a_1 _14926_ (.A1(_11982_),
    .A2(_11972_),
    .A3(_11907_),
    .B1(_11983_),
    .B2(_11974_),
    .X(_11984_));
 sky130_fd_sc_hd__nor2_1 _14927_ (.A(_11979_),
    .B(_11984_),
    .Y(_04002_));
 sky130_fd_sc_hd__buf_1 _14928_ (.A(_11962_),
    .X(_11985_));
 sky130_vsdinv _14929_ (.A(instr_bltu),
    .Y(_11986_));
 sky130_fd_sc_hd__buf_1 _14930_ (.A(_11956_),
    .X(_11987_));
 sky130_fd_sc_hd__o32a_1 _14931_ (.A1(_11982_),
    .A2(_11985_),
    .A3(_11916_),
    .B1(_11986_),
    .B2(_11987_),
    .X(_11988_));
 sky130_fd_sc_hd__nor2_1 _14932_ (.A(_11979_),
    .B(_11988_),
    .Y(_04001_));
 sky130_vsdinv _14933_ (.A(instr_bge),
    .Y(_11989_));
 sky130_fd_sc_hd__o32a_1 _14934_ (.A1(_11982_),
    .A2(_11985_),
    .A3(_11920_),
    .B1(_11989_),
    .B2(_11987_),
    .X(_11990_));
 sky130_fd_sc_hd__nor2_1 _14935_ (.A(_11979_),
    .B(_11990_),
    .Y(_04000_));
 sky130_fd_sc_hd__buf_1 _14936_ (.A(_11978_),
    .X(_11991_));
 sky130_fd_sc_hd__buf_2 _14937_ (.A(_11729_),
    .X(_11992_));
 sky130_vsdinv _14938_ (.A(instr_blt),
    .Y(_11993_));
 sky130_fd_sc_hd__o32a_1 _14939_ (.A1(_11992_),
    .A2(_11985_),
    .A3(_11937_),
    .B1(_11993_),
    .B2(_11987_),
    .X(_11994_));
 sky130_fd_sc_hd__nor2_1 _14940_ (.A(_11991_),
    .B(_11994_),
    .Y(_03999_));
 sky130_vsdinv _14941_ (.A(instr_bne),
    .Y(_11995_));
 sky130_fd_sc_hd__o32a_1 _14942_ (.A1(_11992_),
    .A2(_11985_),
    .A3(_11948_),
    .B1(_11995_),
    .B2(_11987_),
    .X(_11996_));
 sky130_fd_sc_hd__nor2_1 _14943_ (.A(_11991_),
    .B(_11996_),
    .Y(_03998_));
 sky130_fd_sc_hd__clkbuf_2 _14944_ (.A(_11962_),
    .X(_11997_));
 sky130_vsdinv _14945_ (.A(instr_beq),
    .Y(_11998_));
 sky130_fd_sc_hd__clkbuf_4 _14946_ (.A(_11956_),
    .X(_11999_));
 sky130_fd_sc_hd__o32a_1 _14947_ (.A1(_11992_),
    .A2(_11997_),
    .A3(_11951_),
    .B1(_11998_),
    .B2(_11999_),
    .X(_12000_));
 sky130_fd_sc_hd__nor2_1 _14948_ (.A(_11991_),
    .B(_12000_),
    .Y(_03997_));
 sky130_fd_sc_hd__or2_1 _14949_ (.A(\pcpi_timeout_counter[1] ),
    .B(\pcpi_timeout_counter[0] ),
    .X(_12001_));
 sky130_fd_sc_hd__or2_1 _14950_ (.A(\pcpi_timeout_counter[2] ),
    .B(_12001_),
    .X(_12002_));
 sky130_fd_sc_hd__buf_1 _14951_ (.A(_11686_),
    .X(_12003_));
 sky130_fd_sc_hd__a21o_1 _14952_ (.A1(\pcpi_timeout_counter[3] ),
    .A2(_12002_),
    .B1(_12003_),
    .X(_03996_));
 sky130_vsdinv _14953_ (.A(_12002_),
    .Y(_12004_));
 sky130_fd_sc_hd__a221o_1 _14954_ (.A1(\pcpi_timeout_counter[2] ),
    .A2(_12001_),
    .B1(\pcpi_timeout_counter[3] ),
    .B2(_12004_),
    .C1(_12003_),
    .X(_03995_));
 sky130_vsdinv _14955_ (.A(_12001_),
    .Y(_12005_));
 sky130_fd_sc_hd__or2_1 _14956_ (.A(\pcpi_timeout_counter[3] ),
    .B(_12002_),
    .X(_12006_));
 sky130_fd_sc_hd__a221o_1 _14957_ (.A1(\pcpi_timeout_counter[1] ),
    .A2(\pcpi_timeout_counter[0] ),
    .B1(_12005_),
    .B2(_12006_),
    .C1(_12003_),
    .X(_03994_));
 sky130_vsdinv _14958_ (.A(\pcpi_timeout_counter[0] ),
    .Y(_12007_));
 sky130_fd_sc_hd__a21o_1 _14959_ (.A1(_12007_),
    .A2(_12006_),
    .B1(_12003_),
    .X(_03993_));
 sky130_vsdinv _14960_ (.A(_11556_),
    .Y(_12008_));
 sky130_fd_sc_hd__buf_1 _14961_ (.A(_12008_),
    .X(_12009_));
 sky130_fd_sc_hd__buf_2 _14962_ (.A(_12009_),
    .X(_00296_));
 sky130_fd_sc_hd__or2_2 _14963_ (.A(_11585_),
    .B(_11588_),
    .X(_12010_));
 sky130_fd_sc_hd__or4_4 _14964_ (.A(\cpu_state[0] ),
    .B(_11736_),
    .C(_11737_),
    .D(_12010_),
    .X(_12011_));
 sky130_fd_sc_hd__o22ai_1 _14965_ (.A1(_00291_),
    .A2(_11795_),
    .B1(_00296_),
    .B2(_12011_),
    .Y(_03992_));
 sky130_fd_sc_hd__buf_1 _14966_ (.A(_11558_),
    .X(_12012_));
 sky130_fd_sc_hd__buf_1 _14967_ (.A(_12012_),
    .X(_12013_));
 sky130_fd_sc_hd__or3_4 _14968_ (.A(_11585_),
    .B(_11557_),
    .C(_11560_),
    .X(_12014_));
 sky130_fd_sc_hd__o22ai_1 _14969_ (.A1(_12013_),
    .A2(_11795_),
    .B1(_00296_),
    .B2(_12014_),
    .Y(_03991_));
 sky130_fd_sc_hd__clkbuf_2 _14970_ (.A(_11781_),
    .X(_12015_));
 sky130_fd_sc_hd__clkbuf_2 _14971_ (.A(_12015_),
    .X(_12016_));
 sky130_fd_sc_hd__buf_1 _14972_ (.A(_11680_),
    .X(_12017_));
 sky130_fd_sc_hd__o221a_1 _14973_ (.A1(\reg_next_pc[31] ),
    .A2(_12016_),
    .B1(_02530_),
    .B2(_11791_),
    .C1(_12017_),
    .X(_03990_));
 sky130_fd_sc_hd__buf_1 _14974_ (.A(_11774_),
    .X(_12018_));
 sky130_fd_sc_hd__o221a_1 _14975_ (.A1(_11786_),
    .A2(\reg_next_pc[30] ),
    .B1(_12018_),
    .B2(_02529_),
    .C1(_12017_),
    .X(_03989_));
 sky130_fd_sc_hd__o221a_1 _14976_ (.A1(_11786_),
    .A2(\reg_next_pc[29] ),
    .B1(_12018_),
    .B2(_02527_),
    .C1(_12017_),
    .X(_03988_));
 sky130_fd_sc_hd__o221a_1 _14977_ (.A1(_11786_),
    .A2(\reg_next_pc[28] ),
    .B1(_12018_),
    .B2(_02526_),
    .C1(_12017_),
    .X(_03987_));
 sky130_fd_sc_hd__buf_1 _14978_ (.A(_11782_),
    .X(_12019_));
 sky130_fd_sc_hd__buf_1 _14979_ (.A(_11680_),
    .X(_12020_));
 sky130_fd_sc_hd__o221a_1 _14980_ (.A1(_12019_),
    .A2(\reg_next_pc[27] ),
    .B1(_12018_),
    .B2(_02525_),
    .C1(_12020_),
    .X(_03986_));
 sky130_fd_sc_hd__buf_1 _14981_ (.A(_11774_),
    .X(_12021_));
 sky130_fd_sc_hd__o221a_1 _14982_ (.A1(_12019_),
    .A2(\reg_next_pc[26] ),
    .B1(_12021_),
    .B2(_02524_),
    .C1(_12020_),
    .X(_03985_));
 sky130_fd_sc_hd__o221a_1 _14983_ (.A1(_12019_),
    .A2(\reg_next_pc[25] ),
    .B1(_12021_),
    .B2(_02523_),
    .C1(_12020_),
    .X(_03984_));
 sky130_fd_sc_hd__o221a_1 _14984_ (.A1(_12019_),
    .A2(\reg_next_pc[24] ),
    .B1(_12021_),
    .B2(_02522_),
    .C1(_12020_),
    .X(_03983_));
 sky130_fd_sc_hd__buf_1 _14985_ (.A(_11782_),
    .X(_12022_));
 sky130_fd_sc_hd__buf_2 _14986_ (.A(_11679_),
    .X(_12023_));
 sky130_fd_sc_hd__buf_1 _14987_ (.A(_12023_),
    .X(_12024_));
 sky130_fd_sc_hd__o221a_1 _14988_ (.A1(_12022_),
    .A2(\reg_next_pc[23] ),
    .B1(_12021_),
    .B2(_02521_),
    .C1(_12024_),
    .X(_03982_));
 sky130_fd_sc_hd__clkbuf_2 _14989_ (.A(_11774_),
    .X(_12025_));
 sky130_fd_sc_hd__o221a_1 _14990_ (.A1(_12022_),
    .A2(\reg_next_pc[22] ),
    .B1(_12025_),
    .B2(_02520_),
    .C1(_12024_),
    .X(_03981_));
 sky130_fd_sc_hd__o221a_1 _14991_ (.A1(_12022_),
    .A2(\reg_next_pc[21] ),
    .B1(_12025_),
    .B2(_02519_),
    .C1(_12024_),
    .X(_03980_));
 sky130_fd_sc_hd__o221a_1 _14992_ (.A1(_12022_),
    .A2(\reg_next_pc[20] ),
    .B1(_12025_),
    .B2(_02518_),
    .C1(_12024_),
    .X(_03979_));
 sky130_fd_sc_hd__clkbuf_2 _14993_ (.A(_12015_),
    .X(_12026_));
 sky130_fd_sc_hd__buf_1 _14994_ (.A(_12026_),
    .X(_12027_));
 sky130_fd_sc_hd__buf_1 _14995_ (.A(_12023_),
    .X(_12028_));
 sky130_fd_sc_hd__o221a_1 _14996_ (.A1(_12027_),
    .A2(\reg_next_pc[19] ),
    .B1(_12025_),
    .B2(_02516_),
    .C1(_12028_),
    .X(_03978_));
 sky130_fd_sc_hd__buf_2 _14997_ (.A(_11790_),
    .X(_12029_));
 sky130_fd_sc_hd__buf_1 _14998_ (.A(_12029_),
    .X(_12030_));
 sky130_fd_sc_hd__o221a_1 _14999_ (.A1(_12027_),
    .A2(\reg_next_pc[18] ),
    .B1(_12030_),
    .B2(_02515_),
    .C1(_12028_),
    .X(_03977_));
 sky130_fd_sc_hd__o221a_1 _15000_ (.A1(_12027_),
    .A2(\reg_next_pc[17] ),
    .B1(_12030_),
    .B2(_02514_),
    .C1(_12028_),
    .X(_03976_));
 sky130_fd_sc_hd__o221a_1 _15001_ (.A1(_12027_),
    .A2(\reg_next_pc[16] ),
    .B1(_12030_),
    .B2(_02513_),
    .C1(_12028_),
    .X(_03975_));
 sky130_fd_sc_hd__buf_1 _15002_ (.A(_12026_),
    .X(_12031_));
 sky130_fd_sc_hd__buf_1 _15003_ (.A(_12023_),
    .X(_12032_));
 sky130_fd_sc_hd__o221a_1 _15004_ (.A1(_12031_),
    .A2(\reg_next_pc[15] ),
    .B1(_12030_),
    .B2(_02512_),
    .C1(_12032_),
    .X(_03974_));
 sky130_fd_sc_hd__buf_1 _15005_ (.A(_12029_),
    .X(_12033_));
 sky130_fd_sc_hd__o221a_1 _15006_ (.A1(_12031_),
    .A2(\reg_next_pc[14] ),
    .B1(_12033_),
    .B2(_02511_),
    .C1(_12032_),
    .X(_03973_));
 sky130_fd_sc_hd__o221a_1 _15007_ (.A1(_12031_),
    .A2(\reg_next_pc[13] ),
    .B1(_12033_),
    .B2(_02510_),
    .C1(_12032_),
    .X(_03972_));
 sky130_fd_sc_hd__o221a_1 _15008_ (.A1(_12031_),
    .A2(\reg_next_pc[12] ),
    .B1(_12033_),
    .B2(_02509_),
    .C1(_12032_),
    .X(_03971_));
 sky130_fd_sc_hd__buf_1 _15009_ (.A(_12026_),
    .X(_12034_));
 sky130_fd_sc_hd__buf_1 _15010_ (.A(_12023_),
    .X(_12035_));
 sky130_fd_sc_hd__o221a_1 _15011_ (.A1(_12034_),
    .A2(\reg_next_pc[11] ),
    .B1(_12033_),
    .B2(_02508_),
    .C1(_12035_),
    .X(_03970_));
 sky130_fd_sc_hd__buf_1 _15012_ (.A(_12029_),
    .X(_12036_));
 sky130_fd_sc_hd__o221a_1 _15013_ (.A1(_12034_),
    .A2(\reg_next_pc[10] ),
    .B1(_12036_),
    .B2(_02507_),
    .C1(_12035_),
    .X(_03969_));
 sky130_fd_sc_hd__o221a_1 _15014_ (.A1(_12034_),
    .A2(\reg_next_pc[9] ),
    .B1(_12036_),
    .B2(_02537_),
    .C1(_12035_),
    .X(_03968_));
 sky130_fd_sc_hd__o221a_1 _15015_ (.A1(_12034_),
    .A2(\reg_next_pc[8] ),
    .B1(_12036_),
    .B2(_02536_),
    .C1(_12035_),
    .X(_03967_));
 sky130_fd_sc_hd__buf_1 _15016_ (.A(_12026_),
    .X(_12037_));
 sky130_fd_sc_hd__clkbuf_2 _15017_ (.A(_11679_),
    .X(_12038_));
 sky130_fd_sc_hd__buf_1 _15018_ (.A(_12038_),
    .X(_12039_));
 sky130_fd_sc_hd__o221a_1 _15019_ (.A1(_12037_),
    .A2(\reg_next_pc[7] ),
    .B1(_12036_),
    .B2(_02535_),
    .C1(_12039_),
    .X(_03966_));
 sky130_fd_sc_hd__clkbuf_2 _15020_ (.A(_12029_),
    .X(_12040_));
 sky130_fd_sc_hd__o221a_1 _15021_ (.A1(_12037_),
    .A2(\reg_next_pc[6] ),
    .B1(_12040_),
    .B2(_02534_),
    .C1(_12039_),
    .X(_03965_));
 sky130_fd_sc_hd__o221a_1 _15022_ (.A1(_12037_),
    .A2(\reg_next_pc[5] ),
    .B1(_12040_),
    .B2(_02533_),
    .C1(_12039_),
    .X(_03964_));
 sky130_fd_sc_hd__o221a_1 _15023_ (.A1(_12037_),
    .A2(\reg_next_pc[4] ),
    .B1(_12040_),
    .B2(_02532_),
    .C1(_12039_),
    .X(_03963_));
 sky130_fd_sc_hd__clkbuf_2 _15024_ (.A(_12015_),
    .X(_12041_));
 sky130_fd_sc_hd__clkbuf_2 _15025_ (.A(_12041_),
    .X(_12042_));
 sky130_fd_sc_hd__buf_1 _15026_ (.A(_12038_),
    .X(_12043_));
 sky130_fd_sc_hd__o221a_1 _15027_ (.A1(_12042_),
    .A2(\reg_next_pc[3] ),
    .B1(_12040_),
    .B2(_02531_),
    .C1(_12043_),
    .X(_03962_));
 sky130_fd_sc_hd__clkbuf_2 _15028_ (.A(_11790_),
    .X(_12044_));
 sky130_fd_sc_hd__clkbuf_2 _15029_ (.A(_12044_),
    .X(_12045_));
 sky130_fd_sc_hd__o221a_1 _15030_ (.A1(_12042_),
    .A2(\reg_next_pc[2] ),
    .B1(_12045_),
    .B2(_02528_),
    .C1(_12043_),
    .X(_03961_));
 sky130_fd_sc_hd__o221a_1 _15031_ (.A1(_12042_),
    .A2(\reg_next_pc[1] ),
    .B1(_12045_),
    .B2(_02517_),
    .C1(_12043_),
    .X(_03960_));
 sky130_fd_sc_hd__buf_1 _15032_ (.A(\reg_pc[31] ),
    .X(_12046_));
 sky130_fd_sc_hd__o221a_1 _15033_ (.A1(_12042_),
    .A2(_12046_),
    .B1(_12045_),
    .B2(_02581_),
    .C1(_12043_),
    .X(_03959_));
 sky130_fd_sc_hd__buf_1 _15034_ (.A(_12041_),
    .X(_12047_));
 sky130_fd_sc_hd__buf_1 _15035_ (.A(\reg_pc[30] ),
    .X(_12048_));
 sky130_fd_sc_hd__clkbuf_2 _15036_ (.A(_02580_),
    .X(_12049_));
 sky130_fd_sc_hd__buf_1 _15037_ (.A(_12038_),
    .X(_12050_));
 sky130_fd_sc_hd__o221a_1 _15038_ (.A1(_12047_),
    .A2(_12048_),
    .B1(_12045_),
    .B2(_12049_),
    .C1(_12050_),
    .X(_03958_));
 sky130_fd_sc_hd__buf_1 _15039_ (.A(_12044_),
    .X(_12051_));
 sky130_fd_sc_hd__o221a_1 _15040_ (.A1(_12047_),
    .A2(\reg_pc[29] ),
    .B1(_12051_),
    .B2(_02579_),
    .C1(_12050_),
    .X(_03957_));
 sky130_fd_sc_hd__clkbuf_2 _15041_ (.A(\reg_pc[28] ),
    .X(_12052_));
 sky130_fd_sc_hd__o221a_1 _15042_ (.A1(_12047_),
    .A2(_12052_),
    .B1(_12051_),
    .B2(_02578_),
    .C1(_12050_),
    .X(_03956_));
 sky130_fd_sc_hd__o221a_1 _15043_ (.A1(_12047_),
    .A2(\reg_pc[27] ),
    .B1(_12051_),
    .B2(_02577_),
    .C1(_12050_),
    .X(_03955_));
 sky130_fd_sc_hd__buf_1 _15044_ (.A(_12041_),
    .X(_12053_));
 sky130_fd_sc_hd__buf_1 _15045_ (.A(_12038_),
    .X(_12054_));
 sky130_fd_sc_hd__o221a_1 _15046_ (.A1(_12053_),
    .A2(\reg_pc[26] ),
    .B1(_12051_),
    .B2(_02576_),
    .C1(_12054_),
    .X(_03954_));
 sky130_fd_sc_hd__buf_1 _15047_ (.A(_12044_),
    .X(_12055_));
 sky130_fd_sc_hd__o221a_1 _15048_ (.A1(_12053_),
    .A2(\reg_pc[25] ),
    .B1(_12055_),
    .B2(_02575_),
    .C1(_12054_),
    .X(_03953_));
 sky130_fd_sc_hd__o221a_1 _15049_ (.A1(_12053_),
    .A2(\reg_pc[24] ),
    .B1(_12055_),
    .B2(_02574_),
    .C1(_12054_),
    .X(_03952_));
 sky130_fd_sc_hd__o221a_1 _15050_ (.A1(_12053_),
    .A2(\reg_pc[23] ),
    .B1(_12055_),
    .B2(_02573_),
    .C1(_12054_),
    .X(_03951_));
 sky130_fd_sc_hd__buf_1 _15051_ (.A(_12041_),
    .X(_12056_));
 sky130_fd_sc_hd__buf_2 _15052_ (.A(_11679_),
    .X(_12057_));
 sky130_fd_sc_hd__buf_1 _15053_ (.A(_12057_),
    .X(_12058_));
 sky130_fd_sc_hd__o221a_1 _15054_ (.A1(_12056_),
    .A2(\reg_pc[22] ),
    .B1(_12055_),
    .B2(_02572_),
    .C1(_12058_),
    .X(_03950_));
 sky130_fd_sc_hd__clkbuf_2 _15055_ (.A(_12044_),
    .X(_12059_));
 sky130_fd_sc_hd__o221a_1 _15056_ (.A1(_12056_),
    .A2(\reg_pc[21] ),
    .B1(_12059_),
    .B2(_02570_),
    .C1(_12058_),
    .X(_03949_));
 sky130_fd_sc_hd__buf_1 _15057_ (.A(_02569_),
    .X(_12060_));
 sky130_fd_sc_hd__o221a_1 _15058_ (.A1(_12056_),
    .A2(\reg_pc[20] ),
    .B1(_12059_),
    .B2(_12060_),
    .C1(_12058_),
    .X(_03948_));
 sky130_fd_sc_hd__o221a_1 _15059_ (.A1(_12056_),
    .A2(\reg_pc[19] ),
    .B1(_12059_),
    .B2(_02568_),
    .C1(_12058_),
    .X(_03947_));
 sky130_fd_sc_hd__clkbuf_2 _15060_ (.A(_12015_),
    .X(_12061_));
 sky130_fd_sc_hd__buf_1 _15061_ (.A(_12061_),
    .X(_12062_));
 sky130_fd_sc_hd__buf_1 _15062_ (.A(_02567_),
    .X(_12063_));
 sky130_fd_sc_hd__buf_1 _15063_ (.A(_12057_),
    .X(_12064_));
 sky130_fd_sc_hd__o221a_1 _15064_ (.A1(_12062_),
    .A2(\reg_pc[18] ),
    .B1(_12059_),
    .B2(_12063_),
    .C1(_12064_),
    .X(_03946_));
 sky130_fd_sc_hd__buf_2 _15065_ (.A(_11773_),
    .X(_12065_));
 sky130_fd_sc_hd__buf_1 _15066_ (.A(_12065_),
    .X(_12066_));
 sky130_fd_sc_hd__o221a_1 _15067_ (.A1(_12062_),
    .A2(\reg_pc[17] ),
    .B1(_12066_),
    .B2(_02566_),
    .C1(_12064_),
    .X(_03945_));
 sky130_fd_sc_hd__o221a_1 _15068_ (.A1(_12062_),
    .A2(\reg_pc[16] ),
    .B1(_12066_),
    .B2(_02565_),
    .C1(_12064_),
    .X(_03944_));
 sky130_fd_sc_hd__o221a_1 _15069_ (.A1(_12062_),
    .A2(\reg_pc[15] ),
    .B1(_12066_),
    .B2(_02564_),
    .C1(_12064_),
    .X(_03943_));
 sky130_fd_sc_hd__buf_1 _15070_ (.A(_12061_),
    .X(_12067_));
 sky130_fd_sc_hd__buf_1 _15071_ (.A(_12057_),
    .X(_12068_));
 sky130_fd_sc_hd__o221a_1 _15072_ (.A1(_12067_),
    .A2(\reg_pc[14] ),
    .B1(_12066_),
    .B2(_02563_),
    .C1(_12068_),
    .X(_03942_));
 sky130_fd_sc_hd__buf_1 _15073_ (.A(_12065_),
    .X(_12069_));
 sky130_fd_sc_hd__o221a_1 _15074_ (.A1(_12067_),
    .A2(\reg_pc[13] ),
    .B1(_12069_),
    .B2(_02562_),
    .C1(_12068_),
    .X(_03941_));
 sky130_fd_sc_hd__o221a_1 _15075_ (.A1(_12067_),
    .A2(\reg_pc[12] ),
    .B1(_12069_),
    .B2(_02561_),
    .C1(_12068_),
    .X(_03940_));
 sky130_fd_sc_hd__o221a_1 _15076_ (.A1(_12067_),
    .A2(\reg_pc[11] ),
    .B1(_12069_),
    .B2(_02589_),
    .C1(_12068_),
    .X(_03939_));
 sky130_fd_sc_hd__buf_1 _15077_ (.A(_12061_),
    .X(_12070_));
 sky130_fd_sc_hd__buf_1 _15078_ (.A(_02588_),
    .X(_12071_));
 sky130_fd_sc_hd__buf_1 _15079_ (.A(_12057_),
    .X(_12072_));
 sky130_fd_sc_hd__o221a_1 _15080_ (.A1(_12070_),
    .A2(\reg_pc[10] ),
    .B1(_12069_),
    .B2(_12071_),
    .C1(_12072_),
    .X(_03938_));
 sky130_fd_sc_hd__buf_1 _15081_ (.A(_12065_),
    .X(_12073_));
 sky130_fd_sc_hd__o221a_1 _15082_ (.A1(_12070_),
    .A2(\reg_pc[9] ),
    .B1(_12073_),
    .B2(_02587_),
    .C1(_12072_),
    .X(_03937_));
 sky130_fd_sc_hd__buf_1 _15083_ (.A(_02586_),
    .X(_12074_));
 sky130_fd_sc_hd__o221a_1 _15084_ (.A1(_12070_),
    .A2(\reg_pc[8] ),
    .B1(_12073_),
    .B2(_12074_),
    .C1(_12072_),
    .X(_03936_));
 sky130_fd_sc_hd__o221a_1 _15085_ (.A1(_12070_),
    .A2(\reg_pc[7] ),
    .B1(_12073_),
    .B2(_02585_),
    .C1(_12072_),
    .X(_03935_));
 sky130_fd_sc_hd__buf_1 _15086_ (.A(_12061_),
    .X(_12075_));
 sky130_fd_sc_hd__clkbuf_2 _15087_ (.A(\reg_pc[6] ),
    .X(_12076_));
 sky130_fd_sc_hd__buf_1 _15088_ (.A(_02584_),
    .X(_12077_));
 sky130_fd_sc_hd__clkbuf_2 _15089_ (.A(_11544_),
    .X(_12078_));
 sky130_fd_sc_hd__buf_2 _15090_ (.A(_12078_),
    .X(_12079_));
 sky130_fd_sc_hd__o221a_1 _15091_ (.A1(_12075_),
    .A2(_12076_),
    .B1(_12073_),
    .B2(_12077_),
    .C1(_12079_),
    .X(_03934_));
 sky130_fd_sc_hd__clkbuf_2 _15092_ (.A(_12065_),
    .X(_12080_));
 sky130_fd_sc_hd__o221a_1 _15093_ (.A1(_12075_),
    .A2(\reg_pc[5] ),
    .B1(_12080_),
    .B2(_02583_),
    .C1(_12079_),
    .X(_03933_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _15094_ (.A(\reg_pc[4] ),
    .X(_12081_));
 sky130_vsdinv _15095_ (.A(_01475_),
    .Y(_12082_));
 sky130_fd_sc_hd__clkbuf_2 _15096_ (.A(_12082_),
    .X(_02582_));
 sky130_fd_sc_hd__o221a_1 _15097_ (.A1(_12075_),
    .A2(_12081_),
    .B1(_12080_),
    .B2(_02582_),
    .C1(_12079_),
    .X(_03932_));
 sky130_fd_sc_hd__o221a_1 _15098_ (.A1(_12075_),
    .A2(\reg_pc[3] ),
    .B1(_12080_),
    .B2(_02571_),
    .C1(_12079_),
    .X(_03931_));
 sky130_fd_sc_hd__buf_1 _15099_ (.A(_02560_),
    .X(_12083_));
 sky130_fd_sc_hd__clkbuf_4 _15100_ (.A(_12078_),
    .X(_12084_));
 sky130_fd_sc_hd__o221a_1 _15101_ (.A1(_12016_),
    .A2(\reg_pc[2] ),
    .B1(_12080_),
    .B2(_12083_),
    .C1(_12084_),
    .X(_03930_));
 sky130_fd_sc_hd__o221a_1 _15102_ (.A1(_12016_),
    .A2(\reg_pc[1] ),
    .B1(_11791_),
    .B2(_02590_),
    .C1(_12084_),
    .X(_03929_));
 sky130_vsdinv _15103_ (.A(\count_instr[62] ),
    .Y(_12085_));
 sky130_vsdinv _15104_ (.A(\count_instr[61] ),
    .Y(_12086_));
 sky130_vsdinv _15105_ (.A(\count_instr[60] ),
    .Y(_12087_));
 sky130_vsdinv _15106_ (.A(\count_instr[59] ),
    .Y(_12088_));
 sky130_vsdinv _15107_ (.A(\count_instr[58] ),
    .Y(_12089_));
 sky130_vsdinv _15108_ (.A(\count_instr[57] ),
    .Y(_12090_));
 sky130_vsdinv _15109_ (.A(\count_instr[56] ),
    .Y(_12091_));
 sky130_vsdinv _15110_ (.A(\count_instr[55] ),
    .Y(_12092_));
 sky130_vsdinv _15111_ (.A(\count_instr[54] ),
    .Y(_12093_));
 sky130_vsdinv _15112_ (.A(\count_instr[53] ),
    .Y(_12094_));
 sky130_vsdinv _15113_ (.A(\count_instr[52] ),
    .Y(_12095_));
 sky130_vsdinv _15114_ (.A(\count_instr[51] ),
    .Y(_12096_));
 sky130_vsdinv _15115_ (.A(\count_instr[50] ),
    .Y(_12097_));
 sky130_vsdinv _15116_ (.A(\count_instr[49] ),
    .Y(_12098_));
 sky130_vsdinv _15117_ (.A(\count_instr[48] ),
    .Y(_12099_));
 sky130_vsdinv _15118_ (.A(\count_instr[47] ),
    .Y(_12100_));
 sky130_vsdinv _15119_ (.A(\count_instr[46] ),
    .Y(_12101_));
 sky130_vsdinv _15120_ (.A(\count_instr[45] ),
    .Y(_12102_));
 sky130_vsdinv _15121_ (.A(\count_instr[44] ),
    .Y(_12103_));
 sky130_vsdinv _15122_ (.A(\count_instr[43] ),
    .Y(_12104_));
 sky130_vsdinv _15123_ (.A(\count_instr[42] ),
    .Y(_12105_));
 sky130_vsdinv _15124_ (.A(\count_instr[41] ),
    .Y(_12106_));
 sky130_vsdinv _15125_ (.A(\count_instr[40] ),
    .Y(_12107_));
 sky130_vsdinv _15126_ (.A(\count_instr[39] ),
    .Y(_12108_));
 sky130_vsdinv _15127_ (.A(\count_instr[38] ),
    .Y(_12109_));
 sky130_vsdinv _15128_ (.A(\count_instr[37] ),
    .Y(_12110_));
 sky130_vsdinv _15129_ (.A(\count_instr[36] ),
    .Y(_12111_));
 sky130_vsdinv _15130_ (.A(\count_instr[35] ),
    .Y(_12112_));
 sky130_vsdinv _15131_ (.A(\count_instr[34] ),
    .Y(_12113_));
 sky130_vsdinv _15132_ (.A(\count_instr[33] ),
    .Y(_12114_));
 sky130_vsdinv _15133_ (.A(\count_instr[32] ),
    .Y(_12115_));
 sky130_vsdinv _15134_ (.A(\count_instr[31] ),
    .Y(_12116_));
 sky130_vsdinv _15135_ (.A(\count_instr[30] ),
    .Y(_12117_));
 sky130_vsdinv _15136_ (.A(\count_instr[29] ),
    .Y(_12118_));
 sky130_vsdinv _15137_ (.A(\count_instr[28] ),
    .Y(_12119_));
 sky130_vsdinv _15138_ (.A(\count_instr[27] ),
    .Y(_12120_));
 sky130_vsdinv _15139_ (.A(\count_instr[26] ),
    .Y(_12121_));
 sky130_vsdinv _15140_ (.A(\count_instr[25] ),
    .Y(_12122_));
 sky130_vsdinv _15141_ (.A(\count_instr[24] ),
    .Y(_12123_));
 sky130_vsdinv _15142_ (.A(\count_instr[23] ),
    .Y(_12124_));
 sky130_vsdinv _15143_ (.A(\count_instr[22] ),
    .Y(_12125_));
 sky130_vsdinv _15144_ (.A(\count_instr[21] ),
    .Y(_12126_));
 sky130_vsdinv _15145_ (.A(\count_instr[20] ),
    .Y(_12127_));
 sky130_vsdinv _15146_ (.A(\count_instr[19] ),
    .Y(_12128_));
 sky130_vsdinv _15147_ (.A(\count_instr[18] ),
    .Y(_12129_));
 sky130_vsdinv _15148_ (.A(\count_instr[17] ),
    .Y(_12130_));
 sky130_vsdinv _15149_ (.A(\count_instr[16] ),
    .Y(_12131_));
 sky130_vsdinv _15150_ (.A(\count_instr[15] ),
    .Y(_12132_));
 sky130_vsdinv _15151_ (.A(\count_instr[14] ),
    .Y(_12133_));
 sky130_vsdinv _15152_ (.A(\count_instr[13] ),
    .Y(_12134_));
 sky130_vsdinv _15153_ (.A(\count_instr[12] ),
    .Y(_12135_));
 sky130_vsdinv _15154_ (.A(\count_instr[11] ),
    .Y(_12136_));
 sky130_vsdinv _15155_ (.A(\count_instr[10] ),
    .Y(_12137_));
 sky130_vsdinv _15156_ (.A(\count_instr[9] ),
    .Y(_12138_));
 sky130_vsdinv _15157_ (.A(\count_instr[8] ),
    .Y(_12139_));
 sky130_vsdinv _15158_ (.A(\count_instr[7] ),
    .Y(_12140_));
 sky130_vsdinv _15159_ (.A(\count_instr[6] ),
    .Y(_12141_));
 sky130_vsdinv _15160_ (.A(\count_instr[5] ),
    .Y(_12142_));
 sky130_vsdinv _15161_ (.A(\count_instr[4] ),
    .Y(_12143_));
 sky130_vsdinv _15162_ (.A(\count_instr[3] ),
    .Y(_12144_));
 sky130_vsdinv _15163_ (.A(\count_instr[2] ),
    .Y(_12145_));
 sky130_vsdinv _15164_ (.A(\count_instr[1] ),
    .Y(_12146_));
 sky130_vsdinv _15165_ (.A(\count_instr[0] ),
    .Y(_12147_));
 sky130_fd_sc_hd__or2_1 _15166_ (.A(_12147_),
    .B(_11675_),
    .X(_12148_));
 sky130_fd_sc_hd__or3_1 _15167_ (.A(_12145_),
    .B(_12146_),
    .C(_12148_),
    .X(_12149_));
 sky130_fd_sc_hd__or2_2 _15168_ (.A(_12144_),
    .B(_12149_),
    .X(_12150_));
 sky130_fd_sc_hd__or2_1 _15169_ (.A(_12143_),
    .B(_12150_),
    .X(_12151_));
 sky130_fd_sc_hd__or2_2 _15170_ (.A(_12142_),
    .B(_12151_),
    .X(_12152_));
 sky130_fd_sc_hd__or2_1 _15171_ (.A(_12141_),
    .B(_12152_),
    .X(_12153_));
 sky130_fd_sc_hd__or2_2 _15172_ (.A(_12140_),
    .B(_12153_),
    .X(_12154_));
 sky130_fd_sc_hd__or2_1 _15173_ (.A(_12139_),
    .B(_12154_),
    .X(_12155_));
 sky130_fd_sc_hd__or2_1 _15174_ (.A(_12138_),
    .B(_12155_),
    .X(_12156_));
 sky130_fd_sc_hd__or2_1 _15175_ (.A(_12137_),
    .B(_12156_),
    .X(_12157_));
 sky130_fd_sc_hd__or2_1 _15176_ (.A(_12136_),
    .B(_12157_),
    .X(_12158_));
 sky130_fd_sc_hd__or2_1 _15177_ (.A(_12135_),
    .B(_12158_),
    .X(_12159_));
 sky130_fd_sc_hd__or2_2 _15178_ (.A(_12134_),
    .B(_12159_),
    .X(_12160_));
 sky130_fd_sc_hd__or2_1 _15179_ (.A(_12133_),
    .B(_12160_),
    .X(_12161_));
 sky130_fd_sc_hd__or2_2 _15180_ (.A(_12132_),
    .B(_12161_),
    .X(_12162_));
 sky130_fd_sc_hd__or2_1 _15181_ (.A(_12131_),
    .B(_12162_),
    .X(_12163_));
 sky130_fd_sc_hd__or2_1 _15182_ (.A(_12130_),
    .B(_12163_),
    .X(_12164_));
 sky130_fd_sc_hd__or2_1 _15183_ (.A(_12129_),
    .B(_12164_),
    .X(_12165_));
 sky130_fd_sc_hd__or2_2 _15184_ (.A(_12128_),
    .B(_12165_),
    .X(_12166_));
 sky130_fd_sc_hd__or2_1 _15185_ (.A(_12127_),
    .B(_12166_),
    .X(_12167_));
 sky130_fd_sc_hd__or2_2 _15186_ (.A(_12126_),
    .B(_12167_),
    .X(_12168_));
 sky130_fd_sc_hd__or2_1 _15187_ (.A(_12125_),
    .B(_12168_),
    .X(_12169_));
 sky130_fd_sc_hd__or2_2 _15188_ (.A(_12124_),
    .B(_12169_),
    .X(_12170_));
 sky130_fd_sc_hd__or2_1 _15189_ (.A(_12123_),
    .B(_12170_),
    .X(_12171_));
 sky130_fd_sc_hd__or2_1 _15190_ (.A(_12122_),
    .B(_12171_),
    .X(_12172_));
 sky130_fd_sc_hd__or2_1 _15191_ (.A(_12121_),
    .B(_12172_),
    .X(_12173_));
 sky130_fd_sc_hd__or2_2 _15192_ (.A(_12120_),
    .B(_12173_),
    .X(_12174_));
 sky130_fd_sc_hd__or2_1 _15193_ (.A(_12119_),
    .B(_12174_),
    .X(_12175_));
 sky130_fd_sc_hd__or2_1 _15194_ (.A(_12118_),
    .B(_12175_),
    .X(_12176_));
 sky130_fd_sc_hd__or2_1 _15195_ (.A(_12117_),
    .B(_12176_),
    .X(_12177_));
 sky130_fd_sc_hd__or2_2 _15196_ (.A(_12116_),
    .B(_12177_),
    .X(_12178_));
 sky130_fd_sc_hd__or2_1 _15197_ (.A(_12115_),
    .B(_12178_),
    .X(_12179_));
 sky130_fd_sc_hd__or2_2 _15198_ (.A(_12114_),
    .B(_12179_),
    .X(_12180_));
 sky130_fd_sc_hd__or2_1 _15199_ (.A(_12113_),
    .B(_12180_),
    .X(_12181_));
 sky130_fd_sc_hd__or2_2 _15200_ (.A(_12112_),
    .B(_12181_),
    .X(_12182_));
 sky130_fd_sc_hd__or2_1 _15201_ (.A(_12111_),
    .B(_12182_),
    .X(_12183_));
 sky130_fd_sc_hd__or2_2 _15202_ (.A(_12110_),
    .B(_12183_),
    .X(_12184_));
 sky130_fd_sc_hd__or2_1 _15203_ (.A(_12109_),
    .B(_12184_),
    .X(_12185_));
 sky130_fd_sc_hd__or2_1 _15204_ (.A(_12108_),
    .B(_12185_),
    .X(_12186_));
 sky130_fd_sc_hd__or2_1 _15205_ (.A(_12107_),
    .B(_12186_),
    .X(_12187_));
 sky130_fd_sc_hd__or2_1 _15206_ (.A(_12106_),
    .B(_12187_),
    .X(_12188_));
 sky130_fd_sc_hd__or2_1 _15207_ (.A(_12105_),
    .B(_12188_),
    .X(_12189_));
 sky130_fd_sc_hd__or2_2 _15208_ (.A(_12104_),
    .B(_12189_),
    .X(_12190_));
 sky130_fd_sc_hd__or2_1 _15209_ (.A(_12103_),
    .B(_12190_),
    .X(_12191_));
 sky130_fd_sc_hd__or2_2 _15210_ (.A(_12102_),
    .B(_12191_),
    .X(_12192_));
 sky130_fd_sc_hd__or2_1 _15211_ (.A(_12101_),
    .B(_12192_),
    .X(_12193_));
 sky130_fd_sc_hd__or2_1 _15212_ (.A(_12100_),
    .B(_12193_),
    .X(_12194_));
 sky130_fd_sc_hd__or2_1 _15213_ (.A(_12099_),
    .B(_12194_),
    .X(_12195_));
 sky130_fd_sc_hd__or2_1 _15214_ (.A(_12098_),
    .B(_12195_),
    .X(_12196_));
 sky130_fd_sc_hd__or2_1 _15215_ (.A(_12097_),
    .B(_12196_),
    .X(_12197_));
 sky130_fd_sc_hd__or2_2 _15216_ (.A(_12096_),
    .B(_12197_),
    .X(_12198_));
 sky130_fd_sc_hd__or2_1 _15217_ (.A(_12095_),
    .B(_12198_),
    .X(_12199_));
 sky130_fd_sc_hd__or2_1 _15218_ (.A(_12094_),
    .B(_12199_),
    .X(_12200_));
 sky130_fd_sc_hd__or2_1 _15219_ (.A(_12093_),
    .B(_12200_),
    .X(_12201_));
 sky130_fd_sc_hd__or2_2 _15220_ (.A(_12092_),
    .B(_12201_),
    .X(_12202_));
 sky130_fd_sc_hd__or2_1 _15221_ (.A(_12091_),
    .B(_12202_),
    .X(_12203_));
 sky130_fd_sc_hd__or2_2 _15222_ (.A(_12090_),
    .B(_12203_),
    .X(_12204_));
 sky130_fd_sc_hd__or2_1 _15223_ (.A(_12089_),
    .B(_12204_),
    .X(_12205_));
 sky130_fd_sc_hd__or2_2 _15224_ (.A(_12088_),
    .B(_12205_),
    .X(_12206_));
 sky130_fd_sc_hd__or2_1 _15225_ (.A(_12087_),
    .B(_12206_),
    .X(_12207_));
 sky130_fd_sc_hd__or2_2 _15226_ (.A(_12086_),
    .B(_12207_),
    .X(_12208_));
 sky130_fd_sc_hd__or2_1 _15227_ (.A(_12085_),
    .B(_12208_),
    .X(_12209_));
 sky130_vsdinv _15228_ (.A(_12209_),
    .Y(_12210_));
 sky130_vsdinv _15229_ (.A(\count_instr[63] ),
    .Y(_12211_));
 sky130_fd_sc_hd__o221a_1 _15230_ (.A1(\count_instr[63] ),
    .A2(_12210_),
    .B1(_12211_),
    .B2(_12209_),
    .C1(_12084_),
    .X(_03928_));
 sky130_fd_sc_hd__clkbuf_2 _15231_ (.A(_11848_),
    .X(_12212_));
 sky130_fd_sc_hd__buf_2 _15232_ (.A(_12212_),
    .X(_12213_));
 sky130_fd_sc_hd__a211oi_2 _15233_ (.A1(_12085_),
    .A2(_12208_),
    .B1(_12213_),
    .C1(_12210_),
    .Y(_03927_));
 sky130_vsdinv _15234_ (.A(_12207_),
    .Y(_12214_));
 sky130_fd_sc_hd__o211a_1 _15235_ (.A1(\count_instr[61] ),
    .A2(_12214_),
    .B1(_11789_),
    .C1(_12208_),
    .X(_03926_));
 sky130_fd_sc_hd__buf_2 _15236_ (.A(_11978_),
    .X(_12215_));
 sky130_fd_sc_hd__a211oi_2 _15237_ (.A1(_12087_),
    .A2(_12206_),
    .B1(_12215_),
    .C1(_12214_),
    .Y(_03925_));
 sky130_vsdinv _15238_ (.A(_12205_),
    .Y(_12216_));
 sky130_fd_sc_hd__clkbuf_2 _15239_ (.A(_11787_),
    .X(_12217_));
 sky130_fd_sc_hd__buf_1 _15240_ (.A(_12217_),
    .X(_12218_));
 sky130_fd_sc_hd__o211a_1 _15241_ (.A1(\count_instr[59] ),
    .A2(_12216_),
    .B1(_12218_),
    .C1(_12206_),
    .X(_03924_));
 sky130_fd_sc_hd__a211oi_2 _15242_ (.A1(_12089_),
    .A2(_12204_),
    .B1(_12215_),
    .C1(_12216_),
    .Y(_03923_));
 sky130_vsdinv _15243_ (.A(_12203_),
    .Y(_12219_));
 sky130_fd_sc_hd__o211a_1 _15244_ (.A1(\count_instr[57] ),
    .A2(_12219_),
    .B1(_12218_),
    .C1(_12204_),
    .X(_03922_));
 sky130_fd_sc_hd__a211oi_2 _15245_ (.A1(_12091_),
    .A2(_12202_),
    .B1(_12215_),
    .C1(_12219_),
    .Y(_03921_));
 sky130_vsdinv _15246_ (.A(_12201_),
    .Y(_12220_));
 sky130_fd_sc_hd__o211a_1 _15247_ (.A1(\count_instr[55] ),
    .A2(_12220_),
    .B1(_12218_),
    .C1(_12202_),
    .X(_03920_));
 sky130_fd_sc_hd__a211oi_2 _15248_ (.A1(_12093_),
    .A2(_12200_),
    .B1(_12215_),
    .C1(_12220_),
    .Y(_03919_));
 sky130_vsdinv _15249_ (.A(_12199_),
    .Y(_12221_));
 sky130_fd_sc_hd__o211a_1 _15250_ (.A1(\count_instr[53] ),
    .A2(_12221_),
    .B1(_12218_),
    .C1(_12200_),
    .X(_03918_));
 sky130_fd_sc_hd__clkbuf_2 _15251_ (.A(_11767_),
    .X(_12222_));
 sky130_fd_sc_hd__clkbuf_2 _15252_ (.A(_12222_),
    .X(_12223_));
 sky130_fd_sc_hd__a211oi_2 _15253_ (.A1(_12095_),
    .A2(_12198_),
    .B1(_12223_),
    .C1(_12221_),
    .Y(_03917_));
 sky130_vsdinv _15254_ (.A(_12197_),
    .Y(_12224_));
 sky130_fd_sc_hd__clkbuf_2 _15255_ (.A(_12217_),
    .X(_12225_));
 sky130_fd_sc_hd__o211a_1 _15256_ (.A1(\count_instr[51] ),
    .A2(_12224_),
    .B1(_12225_),
    .C1(_12198_),
    .X(_03916_));
 sky130_fd_sc_hd__a211oi_2 _15257_ (.A1(_12097_),
    .A2(_12196_),
    .B1(_12223_),
    .C1(_12224_),
    .Y(_03915_));
 sky130_vsdinv _15258_ (.A(_12195_),
    .Y(_12226_));
 sky130_fd_sc_hd__o211a_1 _15259_ (.A1(\count_instr[49] ),
    .A2(_12226_),
    .B1(_12225_),
    .C1(_12196_),
    .X(_03914_));
 sky130_fd_sc_hd__a211oi_1 _15260_ (.A1(_12099_),
    .A2(_12194_),
    .B1(_12223_),
    .C1(_12226_),
    .Y(_03913_));
 sky130_vsdinv _15261_ (.A(_12193_),
    .Y(_12227_));
 sky130_fd_sc_hd__o211a_1 _15262_ (.A1(\count_instr[47] ),
    .A2(_12227_),
    .B1(_12225_),
    .C1(_12194_),
    .X(_03912_));
 sky130_fd_sc_hd__a211oi_2 _15263_ (.A1(_12101_),
    .A2(_12192_),
    .B1(_12223_),
    .C1(_12227_),
    .Y(_03911_));
 sky130_vsdinv _15264_ (.A(_12191_),
    .Y(_12228_));
 sky130_fd_sc_hd__o211a_1 _15265_ (.A1(\count_instr[45] ),
    .A2(_12228_),
    .B1(_12225_),
    .C1(_12192_),
    .X(_03910_));
 sky130_fd_sc_hd__buf_2 _15266_ (.A(_12222_),
    .X(_12229_));
 sky130_fd_sc_hd__a211oi_2 _15267_ (.A1(_12103_),
    .A2(_12190_),
    .B1(_12229_),
    .C1(_12228_),
    .Y(_03909_));
 sky130_vsdinv _15268_ (.A(_12189_),
    .Y(_12230_));
 sky130_fd_sc_hd__clkbuf_2 _15269_ (.A(_12217_),
    .X(_12231_));
 sky130_fd_sc_hd__o211a_1 _15270_ (.A1(\count_instr[43] ),
    .A2(_12230_),
    .B1(_12231_),
    .C1(_12190_),
    .X(_03908_));
 sky130_fd_sc_hd__a211oi_2 _15271_ (.A1(_12105_),
    .A2(_12188_),
    .B1(_12229_),
    .C1(_12230_),
    .Y(_03907_));
 sky130_vsdinv _15272_ (.A(_12187_),
    .Y(_12232_));
 sky130_fd_sc_hd__o211a_1 _15273_ (.A1(\count_instr[41] ),
    .A2(_12232_),
    .B1(_12231_),
    .C1(_12188_),
    .X(_03906_));
 sky130_fd_sc_hd__a211oi_1 _15274_ (.A1(_12107_),
    .A2(_12186_),
    .B1(_12229_),
    .C1(_12232_),
    .Y(_03905_));
 sky130_vsdinv _15275_ (.A(_12185_),
    .Y(_12233_));
 sky130_fd_sc_hd__o211a_1 _15276_ (.A1(\count_instr[39] ),
    .A2(_12233_),
    .B1(_12231_),
    .C1(_12186_),
    .X(_03904_));
 sky130_fd_sc_hd__a211oi_2 _15277_ (.A1(_12109_),
    .A2(_12184_),
    .B1(_12229_),
    .C1(_12233_),
    .Y(_03903_));
 sky130_vsdinv _15278_ (.A(_12183_),
    .Y(_12234_));
 sky130_fd_sc_hd__o211a_1 _15279_ (.A1(\count_instr[37] ),
    .A2(_12234_),
    .B1(_12231_),
    .C1(_12184_),
    .X(_03902_));
 sky130_fd_sc_hd__buf_2 _15280_ (.A(_12222_),
    .X(_12235_));
 sky130_fd_sc_hd__a211oi_2 _15281_ (.A1(_12111_),
    .A2(_12182_),
    .B1(_12235_),
    .C1(_12234_),
    .Y(_03901_));
 sky130_vsdinv _15282_ (.A(_12181_),
    .Y(_12236_));
 sky130_fd_sc_hd__buf_1 _15283_ (.A(_12217_),
    .X(_12237_));
 sky130_fd_sc_hd__o211a_1 _15284_ (.A1(\count_instr[35] ),
    .A2(_12236_),
    .B1(_12237_),
    .C1(_12182_),
    .X(_03900_));
 sky130_fd_sc_hd__a211oi_2 _15285_ (.A1(_12113_),
    .A2(_12180_),
    .B1(_12235_),
    .C1(_12236_),
    .Y(_03899_));
 sky130_vsdinv _15286_ (.A(_12179_),
    .Y(_12238_));
 sky130_fd_sc_hd__o211a_1 _15287_ (.A1(\count_instr[33] ),
    .A2(_12238_),
    .B1(_12237_),
    .C1(_12180_),
    .X(_03898_));
 sky130_fd_sc_hd__a211oi_2 _15288_ (.A1(_12115_),
    .A2(_12178_),
    .B1(_12235_),
    .C1(_12238_),
    .Y(_03897_));
 sky130_vsdinv _15289_ (.A(_12177_),
    .Y(_12239_));
 sky130_fd_sc_hd__o211a_1 _15290_ (.A1(\count_instr[31] ),
    .A2(_12239_),
    .B1(_12237_),
    .C1(_12178_),
    .X(_03896_));
 sky130_fd_sc_hd__a211oi_2 _15291_ (.A1(_12117_),
    .A2(_12176_),
    .B1(_12235_),
    .C1(_12239_),
    .Y(_03895_));
 sky130_vsdinv _15292_ (.A(_12175_),
    .Y(_12240_));
 sky130_fd_sc_hd__o211a_1 _15293_ (.A1(\count_instr[29] ),
    .A2(_12240_),
    .B1(_12237_),
    .C1(_12176_),
    .X(_03894_));
 sky130_fd_sc_hd__buf_2 _15294_ (.A(_12222_),
    .X(_12241_));
 sky130_fd_sc_hd__a211oi_2 _15295_ (.A1(_12119_),
    .A2(_12174_),
    .B1(_12241_),
    .C1(_12240_),
    .Y(_03893_));
 sky130_vsdinv _15296_ (.A(_12173_),
    .Y(_12242_));
 sky130_fd_sc_hd__clkbuf_2 _15297_ (.A(_11787_),
    .X(_12243_));
 sky130_fd_sc_hd__clkbuf_2 _15298_ (.A(_12243_),
    .X(_12244_));
 sky130_fd_sc_hd__o211a_1 _15299_ (.A1(\count_instr[27] ),
    .A2(_12242_),
    .B1(_12244_),
    .C1(_12174_),
    .X(_03892_));
 sky130_fd_sc_hd__a211oi_2 _15300_ (.A1(_12121_),
    .A2(_12172_),
    .B1(_12241_),
    .C1(_12242_),
    .Y(_03891_));
 sky130_vsdinv _15301_ (.A(_12171_),
    .Y(_12245_));
 sky130_fd_sc_hd__o211a_1 _15302_ (.A1(\count_instr[25] ),
    .A2(_12245_),
    .B1(_12244_),
    .C1(_12172_),
    .X(_03890_));
 sky130_fd_sc_hd__a211oi_2 _15303_ (.A1(_12123_),
    .A2(_12170_),
    .B1(_12241_),
    .C1(_12245_),
    .Y(_03889_));
 sky130_vsdinv _15304_ (.A(_12169_),
    .Y(_12246_));
 sky130_fd_sc_hd__o211a_1 _15305_ (.A1(\count_instr[23] ),
    .A2(_12246_),
    .B1(_12244_),
    .C1(_12170_),
    .X(_03888_));
 sky130_fd_sc_hd__a211oi_2 _15306_ (.A1(_12125_),
    .A2(_12168_),
    .B1(_12241_),
    .C1(_12246_),
    .Y(_03887_));
 sky130_vsdinv _15307_ (.A(_12167_),
    .Y(_12247_));
 sky130_fd_sc_hd__o211a_1 _15308_ (.A1(\count_instr[21] ),
    .A2(_12247_),
    .B1(_12244_),
    .C1(_12168_),
    .X(_03886_));
 sky130_fd_sc_hd__buf_1 _15309_ (.A(_11848_),
    .X(_12248_));
 sky130_fd_sc_hd__buf_2 _15310_ (.A(_12248_),
    .X(_12249_));
 sky130_fd_sc_hd__a211oi_2 _15311_ (.A1(_12127_),
    .A2(_12166_),
    .B1(_12249_),
    .C1(_12247_),
    .Y(_03885_));
 sky130_vsdinv _15312_ (.A(_12165_),
    .Y(_12250_));
 sky130_fd_sc_hd__clkbuf_2 _15313_ (.A(_12243_),
    .X(_12251_));
 sky130_fd_sc_hd__o211a_1 _15314_ (.A1(\count_instr[19] ),
    .A2(_12250_),
    .B1(_12251_),
    .C1(_12166_),
    .X(_03884_));
 sky130_fd_sc_hd__a211oi_2 _15315_ (.A1(_12129_),
    .A2(_12164_),
    .B1(_12249_),
    .C1(_12250_),
    .Y(_03883_));
 sky130_vsdinv _15316_ (.A(_12163_),
    .Y(_12252_));
 sky130_fd_sc_hd__o211a_1 _15317_ (.A1(\count_instr[17] ),
    .A2(_12252_),
    .B1(_12251_),
    .C1(_12164_),
    .X(_03882_));
 sky130_fd_sc_hd__a211oi_2 _15318_ (.A1(_12131_),
    .A2(_12162_),
    .B1(_12249_),
    .C1(_12252_),
    .Y(_03881_));
 sky130_vsdinv _15319_ (.A(_12161_),
    .Y(_12253_));
 sky130_fd_sc_hd__o211a_1 _15320_ (.A1(\count_instr[15] ),
    .A2(_12253_),
    .B1(_12251_),
    .C1(_12162_),
    .X(_03880_));
 sky130_fd_sc_hd__a211oi_2 _15321_ (.A1(_12133_),
    .A2(_12160_),
    .B1(_12249_),
    .C1(_12253_),
    .Y(_03879_));
 sky130_vsdinv _15322_ (.A(_12159_),
    .Y(_12254_));
 sky130_fd_sc_hd__o211a_1 _15323_ (.A1(\count_instr[13] ),
    .A2(_12254_),
    .B1(_12251_),
    .C1(_12160_),
    .X(_03878_));
 sky130_fd_sc_hd__clkbuf_2 _15324_ (.A(_12248_),
    .X(_12255_));
 sky130_fd_sc_hd__a211oi_1 _15325_ (.A1(_12135_),
    .A2(_12158_),
    .B1(_12255_),
    .C1(_12254_),
    .Y(_03877_));
 sky130_vsdinv _15326_ (.A(_12157_),
    .Y(_12256_));
 sky130_fd_sc_hd__buf_1 _15327_ (.A(_12243_),
    .X(_12257_));
 sky130_fd_sc_hd__o211a_1 _15328_ (.A1(\count_instr[11] ),
    .A2(_12256_),
    .B1(_12257_),
    .C1(_12158_),
    .X(_03876_));
 sky130_fd_sc_hd__a211oi_1 _15329_ (.A1(_12137_),
    .A2(_12156_),
    .B1(_12255_),
    .C1(_12256_),
    .Y(_03875_));
 sky130_vsdinv _15330_ (.A(_12155_),
    .Y(_12258_));
 sky130_fd_sc_hd__o211a_1 _15331_ (.A1(\count_instr[9] ),
    .A2(_12258_),
    .B1(_12257_),
    .C1(_12156_),
    .X(_03874_));
 sky130_fd_sc_hd__a211oi_2 _15332_ (.A1(_12139_),
    .A2(_12154_),
    .B1(_12255_),
    .C1(_12258_),
    .Y(_03873_));
 sky130_vsdinv _15333_ (.A(_12153_),
    .Y(_12259_));
 sky130_fd_sc_hd__o211a_1 _15334_ (.A1(\count_instr[7] ),
    .A2(_12259_),
    .B1(_12257_),
    .C1(_12154_),
    .X(_03872_));
 sky130_fd_sc_hd__a211oi_2 _15335_ (.A1(_12141_),
    .A2(_12152_),
    .B1(_12255_),
    .C1(_12259_),
    .Y(_03871_));
 sky130_vsdinv _15336_ (.A(_12151_),
    .Y(_12260_));
 sky130_fd_sc_hd__o211a_1 _15337_ (.A1(\count_instr[5] ),
    .A2(_12260_),
    .B1(_12257_),
    .C1(_12152_),
    .X(_03870_));
 sky130_fd_sc_hd__buf_2 _15338_ (.A(_12248_),
    .X(_12261_));
 sky130_fd_sc_hd__a211oi_2 _15339_ (.A1(_12143_),
    .A2(_12150_),
    .B1(_12261_),
    .C1(_12260_),
    .Y(_03869_));
 sky130_vsdinv _15340_ (.A(_12149_),
    .Y(_12262_));
 sky130_fd_sc_hd__buf_2 _15341_ (.A(_12243_),
    .X(_12263_));
 sky130_fd_sc_hd__o211a_1 _15342_ (.A1(\count_instr[3] ),
    .A2(_12262_),
    .B1(_12263_),
    .C1(_12150_),
    .X(_03868_));
 sky130_fd_sc_hd__buf_1 _15343_ (.A(_12148_),
    .X(_12264_));
 sky130_fd_sc_hd__o21a_1 _15344_ (.A1(_12146_),
    .A2(_12264_),
    .B1(_12145_),
    .X(_12265_));
 sky130_fd_sc_hd__nor3_1 _15345_ (.A(_12213_),
    .B(_12262_),
    .C(_12265_),
    .Y(_03867_));
 sky130_vsdinv _15346_ (.A(_12264_),
    .Y(_12266_));
 sky130_fd_sc_hd__o221a_1 _15347_ (.A1(_12146_),
    .A2(_12264_),
    .B1(\count_instr[1] ),
    .B2(_12266_),
    .C1(_12084_),
    .X(_03866_));
 sky130_fd_sc_hd__o211a_1 _15348_ (.A1(\count_instr[0] ),
    .A2(_11676_),
    .B1(_12263_),
    .C1(_12264_),
    .X(_03865_));
 sky130_fd_sc_hd__or2_1 _15349_ (.A(_11781_),
    .B(_11735_),
    .X(_12267_));
 sky130_fd_sc_hd__o221a_2 _15350_ (.A1(_11568_),
    .A2(_11570_),
    .B1(_11770_),
    .B2(_11772_),
    .C1(_12267_),
    .X(_12268_));
 sky130_fd_sc_hd__buf_1 _15351_ (.A(_12268_),
    .X(_12269_));
 sky130_fd_sc_hd__buf_1 _15352_ (.A(_12269_),
    .X(_12270_));
 sky130_vsdinv _15353_ (.A(_12268_),
    .Y(_12271_));
 sky130_fd_sc_hd__buf_1 _15354_ (.A(_12271_),
    .X(_12272_));
 sky130_fd_sc_hd__buf_1 _15355_ (.A(_12272_),
    .X(_12273_));
 sky130_fd_sc_hd__buf_2 _15356_ (.A(_11739_),
    .X(_12274_));
 sky130_fd_sc_hd__buf_2 _15357_ (.A(_12274_),
    .X(_12275_));
 sky130_fd_sc_hd__clkbuf_2 _15358_ (.A(_12275_),
    .X(_12276_));
 sky130_fd_sc_hd__nor3_2 _15359_ (.A(_11814_),
    .B(_11653_),
    .C(_12276_),
    .Y(_12277_));
 sky130_fd_sc_hd__buf_1 _15360_ (.A(_12078_),
    .X(_12278_));
 sky130_fd_sc_hd__o221a_1 _15361_ (.A1(net126),
    .A2(_12270_),
    .B1(_12273_),
    .B2(_12277_),
    .C1(_12278_),
    .X(_03864_));
 sky130_fd_sc_hd__buf_1 _15362_ (.A(\irq_pending[30] ),
    .X(_12279_));
 sky130_fd_sc_hd__buf_2 _15363_ (.A(_11571_),
    .X(_12280_));
 sky130_fd_sc_hd__buf_1 _15364_ (.A(_12280_),
    .X(_12281_));
 sky130_fd_sc_hd__and3_1 _15365_ (.A(_11651_),
    .B(_12279_),
    .C(_12281_),
    .X(_12282_));
 sky130_fd_sc_hd__o221a_1 _15366_ (.A1(net125),
    .A2(_12270_),
    .B1(_12273_),
    .B2(_12282_),
    .C1(_12278_),
    .X(_03863_));
 sky130_fd_sc_hd__nor3_2 _15367_ (.A(_11833_),
    .B(_11652_),
    .C(_12276_),
    .Y(_12283_));
 sky130_fd_sc_hd__o221a_1 _15368_ (.A1(net123),
    .A2(_12270_),
    .B1(_12273_),
    .B2(_12283_),
    .C1(_12278_),
    .X(_03862_));
 sky130_fd_sc_hd__buf_1 _15369_ (.A(\irq_pending[28] ),
    .X(_12284_));
 sky130_fd_sc_hd__and3_1 _15370_ (.A(_11650_),
    .B(_12284_),
    .C(_12281_),
    .X(_12285_));
 sky130_fd_sc_hd__o221a_1 _15371_ (.A1(net122),
    .A2(_12270_),
    .B1(_12273_),
    .B2(_12285_),
    .C1(_12278_),
    .X(_03861_));
 sky130_fd_sc_hd__buf_1 _15372_ (.A(_12269_),
    .X(_12286_));
 sky130_fd_sc_hd__buf_1 _15373_ (.A(_12272_),
    .X(_12287_));
 sky130_fd_sc_hd__nor3_1 _15374_ (.A(_11834_),
    .B(_11634_),
    .C(_12276_),
    .Y(_12288_));
 sky130_fd_sc_hd__buf_1 _15375_ (.A(_12078_),
    .X(_12289_));
 sky130_fd_sc_hd__o221a_1 _15376_ (.A1(net121),
    .A2(_12286_),
    .B1(_12287_),
    .B2(_12288_),
    .C1(_12289_),
    .X(_03860_));
 sky130_fd_sc_hd__buf_1 _15377_ (.A(\irq_pending[26] ),
    .X(_12290_));
 sky130_fd_sc_hd__and3_1 _15378_ (.A(_11632_),
    .B(_12290_),
    .C(_12281_),
    .X(_12291_));
 sky130_fd_sc_hd__o221a_1 _15379_ (.A1(net120),
    .A2(_12286_),
    .B1(_12287_),
    .B2(_12291_),
    .C1(_12289_),
    .X(_03859_));
 sky130_fd_sc_hd__nor3_1 _15380_ (.A(_11838_),
    .B(_11633_),
    .C(_12276_),
    .Y(_12292_));
 sky130_fd_sc_hd__o221a_1 _15381_ (.A1(net119),
    .A2(_12286_),
    .B1(_12287_),
    .B2(_12292_),
    .C1(_12289_),
    .X(_03858_));
 sky130_fd_sc_hd__buf_1 _15382_ (.A(\irq_pending[24] ),
    .X(_12293_));
 sky130_fd_sc_hd__and3_1 _15383_ (.A(_11631_),
    .B(_12293_),
    .C(_12281_),
    .X(_12294_));
 sky130_fd_sc_hd__o221a_1 _15384_ (.A1(net118),
    .A2(_12286_),
    .B1(_12287_),
    .B2(_12294_),
    .C1(_12289_),
    .X(_03857_));
 sky130_fd_sc_hd__buf_1 _15385_ (.A(_12269_),
    .X(_12295_));
 sky130_fd_sc_hd__buf_1 _15386_ (.A(_12272_),
    .X(_12296_));
 sky130_fd_sc_hd__clkbuf_2 _15387_ (.A(_12275_),
    .X(_12297_));
 sky130_fd_sc_hd__nor3_1 _15388_ (.A(_11839_),
    .B(_11665_),
    .C(_12297_),
    .Y(_12298_));
 sky130_fd_sc_hd__clkbuf_2 _15389_ (.A(_11544_),
    .X(_12299_));
 sky130_fd_sc_hd__buf_1 _15390_ (.A(_12299_),
    .X(_12300_));
 sky130_fd_sc_hd__o221a_1 _15391_ (.A1(net117),
    .A2(_12295_),
    .B1(_12296_),
    .B2(_12298_),
    .C1(_12300_),
    .X(_03856_));
 sky130_fd_sc_hd__buf_1 _15392_ (.A(\irq_pending[22] ),
    .X(_12301_));
 sky130_fd_sc_hd__clkbuf_4 _15393_ (.A(_11571_),
    .X(_12302_));
 sky130_fd_sc_hd__clkbuf_2 _15394_ (.A(_12302_),
    .X(_12303_));
 sky130_fd_sc_hd__and3_1 _15395_ (.A(_11663_),
    .B(_12301_),
    .C(_12303_),
    .X(_12304_));
 sky130_fd_sc_hd__o221a_1 _15396_ (.A1(net116),
    .A2(_12295_),
    .B1(_12296_),
    .B2(_12304_),
    .C1(_12300_),
    .X(_03855_));
 sky130_fd_sc_hd__nor3_2 _15397_ (.A(_11845_),
    .B(_11664_),
    .C(_12297_),
    .Y(_12305_));
 sky130_fd_sc_hd__o221a_1 _15398_ (.A1(net115),
    .A2(_12295_),
    .B1(_12296_),
    .B2(_12305_),
    .C1(_12300_),
    .X(_03854_));
 sky130_fd_sc_hd__buf_1 _15399_ (.A(\irq_pending[20] ),
    .X(_12306_));
 sky130_fd_sc_hd__and3_1 _15400_ (.A(_11662_),
    .B(_12306_),
    .C(_12303_),
    .X(_12307_));
 sky130_fd_sc_hd__o221a_1 _15401_ (.A1(net114),
    .A2(_12295_),
    .B1(_12296_),
    .B2(_12307_),
    .C1(_12300_),
    .X(_03853_));
 sky130_fd_sc_hd__buf_1 _15402_ (.A(_12269_),
    .X(_12308_));
 sky130_fd_sc_hd__buf_1 _15403_ (.A(_12272_),
    .X(_12309_));
 sky130_fd_sc_hd__nor3_2 _15404_ (.A(_11846_),
    .B(_11626_),
    .C(_12297_),
    .Y(_12310_));
 sky130_fd_sc_hd__buf_1 _15405_ (.A(_12299_),
    .X(_12311_));
 sky130_fd_sc_hd__o221a_1 _15406_ (.A1(net112),
    .A2(_12308_),
    .B1(_12309_),
    .B2(_12310_),
    .C1(_12311_),
    .X(_03852_));
 sky130_vsdinv _15407_ (.A(\irq_mask[18] ),
    .Y(_12312_));
 sky130_fd_sc_hd__buf_1 _15408_ (.A(\irq_pending[18] ),
    .X(_12313_));
 sky130_fd_sc_hd__and3_1 _15409_ (.A(_12312_),
    .B(_12313_),
    .C(_12303_),
    .X(_12314_));
 sky130_fd_sc_hd__o221a_1 _15410_ (.A1(net111),
    .A2(_12308_),
    .B1(_12309_),
    .B2(_12314_),
    .C1(_12311_),
    .X(_03851_));
 sky130_fd_sc_hd__nor3_2 _15411_ (.A(_11852_),
    .B(_11625_),
    .C(_12297_),
    .Y(_12315_));
 sky130_fd_sc_hd__o221a_1 _15412_ (.A1(net110),
    .A2(_12308_),
    .B1(_12309_),
    .B2(_12315_),
    .C1(_12311_),
    .X(_03850_));
 sky130_fd_sc_hd__clkbuf_2 _15413_ (.A(_12275_),
    .X(_12316_));
 sky130_fd_sc_hd__nor3_2 _15414_ (.A(_11853_),
    .B(_11627_),
    .C(_12316_),
    .Y(_12317_));
 sky130_fd_sc_hd__o221a_1 _15415_ (.A1(net109),
    .A2(_12308_),
    .B1(_12309_),
    .B2(_12317_),
    .C1(_12311_),
    .X(_03849_));
 sky130_fd_sc_hd__buf_1 _15416_ (.A(_12268_),
    .X(_12318_));
 sky130_fd_sc_hd__buf_1 _15417_ (.A(_12318_),
    .X(_12319_));
 sky130_fd_sc_hd__clkbuf_2 _15418_ (.A(_12271_),
    .X(_12320_));
 sky130_fd_sc_hd__buf_1 _15419_ (.A(_12320_),
    .X(_12321_));
 sky130_fd_sc_hd__buf_1 _15420_ (.A(\irq_pending[15] ),
    .X(_12322_));
 sky130_fd_sc_hd__and3_1 _15421_ (.A(_11645_),
    .B(_12322_),
    .C(_12303_),
    .X(_12323_));
 sky130_fd_sc_hd__buf_1 _15422_ (.A(_12299_),
    .X(_12324_));
 sky130_fd_sc_hd__o221a_1 _15423_ (.A1(net108),
    .A2(_12319_),
    .B1(_12321_),
    .B2(_12323_),
    .C1(_12324_),
    .X(_03848_));
 sky130_fd_sc_hd__nor3_1 _15424_ (.A(_11858_),
    .B(_11647_),
    .C(_12316_),
    .Y(_12325_));
 sky130_fd_sc_hd__o221a_1 _15425_ (.A1(net107),
    .A2(_12319_),
    .B1(_12321_),
    .B2(_12325_),
    .C1(_12324_),
    .X(_03847_));
 sky130_fd_sc_hd__buf_1 _15426_ (.A(\irq_pending[13] ),
    .X(_12326_));
 sky130_fd_sc_hd__buf_1 _15427_ (.A(_12302_),
    .X(_12327_));
 sky130_fd_sc_hd__and3_1 _15428_ (.A(_11644_),
    .B(_12326_),
    .C(_12327_),
    .X(_12328_));
 sky130_fd_sc_hd__o221a_1 _15429_ (.A1(net106),
    .A2(_12319_),
    .B1(_12321_),
    .B2(_12328_),
    .C1(_12324_),
    .X(_03846_));
 sky130_fd_sc_hd__nor3_1 _15430_ (.A(_11861_),
    .B(_11646_),
    .C(_12316_),
    .Y(_12329_));
 sky130_fd_sc_hd__o221a_1 _15431_ (.A1(net105),
    .A2(_12319_),
    .B1(_12321_),
    .B2(_12329_),
    .C1(_12324_),
    .X(_03845_));
 sky130_fd_sc_hd__buf_1 _15432_ (.A(_12318_),
    .X(_12330_));
 sky130_fd_sc_hd__buf_1 _15433_ (.A(_12320_),
    .X(_12331_));
 sky130_fd_sc_hd__buf_1 _15434_ (.A(\irq_pending[11] ),
    .X(_12332_));
 sky130_fd_sc_hd__and3_1 _15435_ (.A(_11657_),
    .B(_12332_),
    .C(_12327_),
    .X(_12333_));
 sky130_fd_sc_hd__buf_1 _15436_ (.A(_12299_),
    .X(_12334_));
 sky130_fd_sc_hd__o221a_1 _15437_ (.A1(net104),
    .A2(_12330_),
    .B1(_12331_),
    .B2(_12333_),
    .C1(_12334_),
    .X(_03844_));
 sky130_fd_sc_hd__nor3_1 _15438_ (.A(_11864_),
    .B(_11659_),
    .C(_12316_),
    .Y(_12335_));
 sky130_fd_sc_hd__o221a_1 _15439_ (.A1(net103),
    .A2(_12330_),
    .B1(_12331_),
    .B2(_12335_),
    .C1(_12334_),
    .X(_03843_));
 sky130_fd_sc_hd__buf_1 _15440_ (.A(\irq_pending[9] ),
    .X(_12336_));
 sky130_fd_sc_hd__and3_1 _15441_ (.A(_11656_),
    .B(_12336_),
    .C(_12327_),
    .X(_12337_));
 sky130_fd_sc_hd__o221a_1 _15442_ (.A1(net133),
    .A2(_12330_),
    .B1(_12331_),
    .B2(_12337_),
    .C1(_12334_),
    .X(_03842_));
 sky130_fd_sc_hd__clkbuf_2 _15443_ (.A(_12274_),
    .X(_12338_));
 sky130_fd_sc_hd__nor3_1 _15444_ (.A(_11866_),
    .B(_11658_),
    .C(_12338_),
    .Y(_12339_));
 sky130_fd_sc_hd__o221a_1 _15445_ (.A1(net132),
    .A2(_12330_),
    .B1(_12331_),
    .B2(_12339_),
    .C1(_12334_),
    .X(_03841_));
 sky130_fd_sc_hd__buf_1 _15446_ (.A(_12318_),
    .X(_12340_));
 sky130_fd_sc_hd__buf_1 _15447_ (.A(_12320_),
    .X(_12341_));
 sky130_fd_sc_hd__buf_1 _15448_ (.A(\irq_pending[7] ),
    .X(_12342_));
 sky130_fd_sc_hd__and3_1 _15449_ (.A(_11638_),
    .B(_12342_),
    .C(_12327_),
    .X(_12343_));
 sky130_fd_sc_hd__buf_1 _15450_ (.A(_11565_),
    .X(_12344_));
 sky130_fd_sc_hd__o221a_1 _15451_ (.A1(net131),
    .A2(_12340_),
    .B1(_12341_),
    .B2(_12343_),
    .C1(_12344_),
    .X(_03840_));
 sky130_fd_sc_hd__nor3_1 _15452_ (.A(_11870_),
    .B(_11640_),
    .C(_12338_),
    .Y(_12345_));
 sky130_fd_sc_hd__o221a_1 _15453_ (.A1(net130),
    .A2(_12340_),
    .B1(_12341_),
    .B2(_12345_),
    .C1(_12344_),
    .X(_03839_));
 sky130_fd_sc_hd__buf_1 _15454_ (.A(\irq_pending[5] ),
    .X(_12346_));
 sky130_fd_sc_hd__buf_1 _15455_ (.A(_12302_),
    .X(_12347_));
 sky130_fd_sc_hd__and3_1 _15456_ (.A(_11637_),
    .B(_12346_),
    .C(_12347_),
    .X(_12348_));
 sky130_fd_sc_hd__o221a_1 _15457_ (.A1(net129),
    .A2(_12340_),
    .B1(_12341_),
    .B2(_12348_),
    .C1(_12344_),
    .X(_03838_));
 sky130_fd_sc_hd__nor3_1 _15458_ (.A(_11872_),
    .B(_11639_),
    .C(_12338_),
    .Y(_12349_));
 sky130_fd_sc_hd__o221a_1 _15459_ (.A1(net128),
    .A2(_12340_),
    .B1(_12341_),
    .B2(_12349_),
    .C1(_12344_),
    .X(_03837_));
 sky130_fd_sc_hd__buf_1 _15460_ (.A(_12318_),
    .X(_12350_));
 sky130_fd_sc_hd__buf_1 _15461_ (.A(_12320_),
    .X(_12351_));
 sky130_fd_sc_hd__nor3_2 _15462_ (.A(_11873_),
    .B(_11622_),
    .C(_12338_),
    .Y(_12352_));
 sky130_fd_sc_hd__buf_1 _15463_ (.A(_11565_),
    .X(_12353_));
 sky130_fd_sc_hd__o221a_1 _15464_ (.A1(net127),
    .A2(_12350_),
    .B1(_12351_),
    .B2(_12352_),
    .C1(_12353_),
    .X(_03836_));
 sky130_fd_sc_hd__buf_1 _15465_ (.A(_11620_),
    .X(_12354_));
 sky130_fd_sc_hd__buf_1 _15466_ (.A(\irq_pending[2] ),
    .X(_12355_));
 sky130_fd_sc_hd__and3_1 _15467_ (.A(_12354_),
    .B(_12355_),
    .C(_12347_),
    .X(_12356_));
 sky130_fd_sc_hd__o221a_1 _15468_ (.A1(net124),
    .A2(_12350_),
    .B1(_12351_),
    .B2(_12356_),
    .C1(_12353_),
    .X(_03835_));
 sky130_fd_sc_hd__buf_1 _15469_ (.A(_11619_),
    .X(_12357_));
 sky130_fd_sc_hd__buf_1 _15470_ (.A(\irq_pending[1] ),
    .X(_12358_));
 sky130_fd_sc_hd__and3_1 _15471_ (.A(_12357_),
    .B(_12358_),
    .C(_12347_),
    .X(_12359_));
 sky130_fd_sc_hd__o221a_1 _15472_ (.A1(net113),
    .A2(_12350_),
    .B1(_12351_),
    .B2(_12359_),
    .C1(_12353_),
    .X(_03834_));
 sky130_vsdinv _15473_ (.A(\irq_mask[0] ),
    .Y(_12360_));
 sky130_fd_sc_hd__and3_1 _15474_ (.A(_12360_),
    .B(\irq_pending[0] ),
    .C(_12347_),
    .X(_12361_));
 sky130_fd_sc_hd__o221a_1 _15475_ (.A1(net102),
    .A2(_12350_),
    .B1(_12351_),
    .B2(_12361_),
    .C1(_12353_),
    .X(_03833_));
 sky130_vsdinv _15476_ (.A(\cpu_state[3] ),
    .Y(_12362_));
 sky130_fd_sc_hd__or2_1 _15477_ (.A(_12362_),
    .B(_11763_),
    .X(_12363_));
 sky130_fd_sc_hd__clkbuf_2 _15478_ (.A(_12363_),
    .X(_12364_));
 sky130_fd_sc_hd__buf_2 _15479_ (.A(\cpu_state[3] ),
    .X(_12365_));
 sky130_fd_sc_hd__buf_1 _15480_ (.A(_12365_),
    .X(_12366_));
 sky130_fd_sc_hd__clkbuf_4 _15481_ (.A(_12366_),
    .X(_12367_));
 sky130_fd_sc_hd__nor2_4 _15482_ (.A(instr_ecall_ebreak),
    .B(pcpi_timeout),
    .Y(_00311_));
 sky130_fd_sc_hd__nand2_1 _15483_ (.A(_11748_),
    .B(_00311_),
    .Y(_12368_));
 sky130_fd_sc_hd__a31o_1 _15484_ (.A1(_12367_),
    .A2(_00310_),
    .A3(_12368_),
    .B1(_12212_),
    .X(_12369_));
 sky130_fd_sc_hd__a21oi_1 _15485_ (.A1(_11685_),
    .A2(_12364_),
    .B1(_12369_),
    .Y(_03832_));
 sky130_fd_sc_hd__inv_2 _15486_ (.A(_11591_),
    .Y(_00290_));
 sky130_fd_sc_hd__o31a_1 _15487_ (.A1(_11588_),
    .A2(_11590_),
    .A3(net237),
    .B1(_00290_),
    .X(_12370_));
 sky130_fd_sc_hd__a21oi_1 _15488_ (.A1(net237),
    .A2(_11550_),
    .B1(_12370_),
    .Y(_12371_));
 sky130_vsdinv _15489_ (.A(net237),
    .Y(_12372_));
 sky130_fd_sc_hd__o22a_1 _15490_ (.A1(_11582_),
    .A2(_12371_),
    .B1(_12372_),
    .B2(net65),
    .X(_12373_));
 sky130_fd_sc_hd__nor2_1 _15491_ (.A(_11991_),
    .B(_12373_),
    .Y(_03831_));
 sky130_fd_sc_hd__or4_4 _15492_ (.A(\irq_pending[21] ),
    .B(_12306_),
    .C(\irq_pending[23] ),
    .D(_12301_),
    .X(_12374_));
 sky130_fd_sc_hd__or4_4 _15493_ (.A(\irq_pending[17] ),
    .B(\irq_pending[16] ),
    .C(\irq_pending[19] ),
    .D(_12313_),
    .X(_12375_));
 sky130_fd_sc_hd__or4_4 _15494_ (.A(\irq_pending[29] ),
    .B(_12284_),
    .C(\irq_pending[31] ),
    .D(_12279_),
    .X(_12376_));
 sky130_fd_sc_hd__or4_4 _15495_ (.A(\irq_pending[25] ),
    .B(_12293_),
    .C(\irq_pending[27] ),
    .D(_12290_),
    .X(_12377_));
 sky130_fd_sc_hd__or4_4 _15496_ (.A(_12374_),
    .B(_12375_),
    .C(_12376_),
    .D(_12377_),
    .X(_12378_));
 sky130_fd_sc_hd__or4_1 _15497_ (.A(_12346_),
    .B(\irq_pending[4] ),
    .C(_12342_),
    .D(\irq_pending[6] ),
    .X(_12379_));
 sky130_fd_sc_hd__or4_4 _15498_ (.A(_12358_),
    .B(\irq_pending[0] ),
    .C(\irq_pending[3] ),
    .D(_12355_),
    .X(_12380_));
 sky130_fd_sc_hd__or4_4 _15499_ (.A(_12326_),
    .B(\irq_pending[12] ),
    .C(_12322_),
    .D(\irq_pending[14] ),
    .X(_12381_));
 sky130_fd_sc_hd__or4_4 _15500_ (.A(_12336_),
    .B(\irq_pending[8] ),
    .C(_12332_),
    .D(\irq_pending[10] ),
    .X(_12382_));
 sky130_fd_sc_hd__or4_1 _15501_ (.A(_12379_),
    .B(_12380_),
    .C(_12381_),
    .D(_12382_),
    .X(_12383_));
 sky130_fd_sc_hd__or2_2 _15502_ (.A(_12378_),
    .B(_12383_),
    .X(_12384_));
 sky130_fd_sc_hd__inv_2 _15503_ (.A(_12384_),
    .Y(_02410_));
 sky130_fd_sc_hd__clkbuf_2 _15504_ (.A(_11791_),
    .X(_00322_));
 sky130_fd_sc_hd__or2_1 _15505_ (.A(_11578_),
    .B(_11672_),
    .X(_12385_));
 sky130_fd_sc_hd__or2_2 _15506_ (.A(_11673_),
    .B(_12385_),
    .X(_12386_));
 sky130_fd_sc_hd__nor3_1 _15507_ (.A(_00322_),
    .B(_12384_),
    .C(_12386_),
    .Y(_03830_));
 sky130_fd_sc_hd__or3_1 _15508_ (.A(_11891_),
    .B(instr_sltu),
    .C(instr_slt),
    .X(_12387_));
 sky130_fd_sc_hd__clkbuf_4 _15509_ (.A(_11565_),
    .X(_12388_));
 sky130_fd_sc_hd__buf_4 _15510_ (.A(_11942_),
    .X(_12389_));
 sky130_fd_sc_hd__o311a_2 _15511_ (.A1(instr_sltiu),
    .A2(instr_slti),
    .A3(_12387_),
    .B1(_12388_),
    .C1(_12389_),
    .X(_03829_));
 sky130_vsdinv _15512_ (.A(_11806_),
    .Y(_12390_));
 sky130_fd_sc_hd__or2_1 _15513_ (.A(_11545_),
    .B(_11555_),
    .X(_12391_));
 sky130_fd_sc_hd__or2_2 _15514_ (.A(_12390_),
    .B(_12391_),
    .X(_12392_));
 sky130_vsdinv _15515_ (.A(_12392_),
    .Y(_03828_));
 sky130_fd_sc_hd__clkbuf_2 _15516_ (.A(_11978_),
    .X(_12393_));
 sky130_fd_sc_hd__nor2_1 _15517_ (.A(_12393_),
    .B(_12006_),
    .Y(_03827_));
 sky130_fd_sc_hd__clkbuf_2 _15518_ (.A(_11680_),
    .X(_12394_));
 sky130_fd_sc_hd__and2_1 _15519_ (.A(_12394_),
    .B(_02435_),
    .X(_03826_));
 sky130_fd_sc_hd__and2_1 _15520_ (.A(_12394_),
    .B(_02434_),
    .X(_03825_));
 sky130_fd_sc_hd__and2_1 _15521_ (.A(_12394_),
    .B(_02432_),
    .X(_03824_));
 sky130_fd_sc_hd__clkbuf_2 _15522_ (.A(_11678_),
    .X(_12395_));
 sky130_fd_sc_hd__clkbuf_4 _15523_ (.A(_12395_),
    .X(_12396_));
 sky130_fd_sc_hd__buf_1 _15524_ (.A(_12396_),
    .X(_12397_));
 sky130_fd_sc_hd__and2_1 _15525_ (.A(_12397_),
    .B(_02431_),
    .X(_03823_));
 sky130_fd_sc_hd__and2_1 _15526_ (.A(_12397_),
    .B(_02430_),
    .X(_03822_));
 sky130_fd_sc_hd__and2_1 _15527_ (.A(_12397_),
    .B(_02429_),
    .X(_03821_));
 sky130_fd_sc_hd__and2_1 _15528_ (.A(_12397_),
    .B(_02428_),
    .X(_03820_));
 sky130_fd_sc_hd__buf_1 _15529_ (.A(_12396_),
    .X(_12398_));
 sky130_fd_sc_hd__and2_1 _15530_ (.A(_12398_),
    .B(_02427_),
    .X(_03819_));
 sky130_fd_sc_hd__and2_1 _15531_ (.A(_12398_),
    .B(_02426_),
    .X(_03818_));
 sky130_fd_sc_hd__and2_1 _15532_ (.A(_12398_),
    .B(_02425_),
    .X(_03817_));
 sky130_fd_sc_hd__and2_1 _15533_ (.A(_12398_),
    .B(_02424_),
    .X(_03816_));
 sky130_fd_sc_hd__buf_1 _15534_ (.A(_12396_),
    .X(_12399_));
 sky130_fd_sc_hd__and2_1 _15535_ (.A(_12399_),
    .B(_02423_),
    .X(_03815_));
 sky130_fd_sc_hd__and2_1 _15536_ (.A(_12399_),
    .B(_02421_),
    .X(_03814_));
 sky130_fd_sc_hd__and2_1 _15537_ (.A(_12399_),
    .B(_02420_),
    .X(_03813_));
 sky130_fd_sc_hd__and2_1 _15538_ (.A(_12399_),
    .B(_02419_),
    .X(_03812_));
 sky130_fd_sc_hd__buf_1 _15539_ (.A(_12395_),
    .X(_12400_));
 sky130_fd_sc_hd__buf_1 _15540_ (.A(_12400_),
    .X(_12401_));
 sky130_fd_sc_hd__and2_1 _15541_ (.A(_12401_),
    .B(_02418_),
    .X(_03811_));
 sky130_fd_sc_hd__and2_1 _15542_ (.A(_12401_),
    .B(_02417_),
    .X(_03810_));
 sky130_fd_sc_hd__and2_1 _15543_ (.A(_12401_),
    .B(_02416_),
    .X(_03809_));
 sky130_fd_sc_hd__and2_1 _15544_ (.A(_12401_),
    .B(_02415_),
    .X(_03808_));
 sky130_fd_sc_hd__buf_1 _15545_ (.A(_12400_),
    .X(_12402_));
 sky130_fd_sc_hd__and2_1 _15546_ (.A(_12402_),
    .B(_02414_),
    .X(_03807_));
 sky130_fd_sc_hd__and2_1 _15547_ (.A(_12402_),
    .B(_02413_),
    .X(_03806_));
 sky130_fd_sc_hd__and2_1 _15548_ (.A(_12402_),
    .B(_02412_),
    .X(_03805_));
 sky130_fd_sc_hd__and2_1 _15549_ (.A(_12402_),
    .B(_02442_),
    .X(_03804_));
 sky130_fd_sc_hd__buf_1 _15550_ (.A(_12400_),
    .X(_12403_));
 sky130_fd_sc_hd__and2_1 _15551_ (.A(_12403_),
    .B(_02441_),
    .X(_03803_));
 sky130_fd_sc_hd__and2_1 _15552_ (.A(_12403_),
    .B(_02440_),
    .X(_03802_));
 sky130_fd_sc_hd__and2_1 _15553_ (.A(_12403_),
    .B(_02439_),
    .X(_03801_));
 sky130_fd_sc_hd__and2_1 _15554_ (.A(_12403_),
    .B(_02438_),
    .X(_03800_));
 sky130_fd_sc_hd__buf_1 _15555_ (.A(_12400_),
    .X(_12404_));
 sky130_fd_sc_hd__and2_1 _15556_ (.A(_12404_),
    .B(_02437_),
    .X(_03799_));
 sky130_fd_sc_hd__and2_1 _15557_ (.A(_12404_),
    .B(_02436_),
    .X(_03798_));
 sky130_fd_sc_hd__and2_1 _15558_ (.A(_12404_),
    .B(_02433_),
    .X(_03797_));
 sky130_fd_sc_hd__and2_1 _15559_ (.A(_12404_),
    .B(_02422_),
    .X(_03796_));
 sky130_fd_sc_hd__buf_1 _15560_ (.A(_12395_),
    .X(_12405_));
 sky130_fd_sc_hd__clkbuf_4 _15561_ (.A(_12405_),
    .X(_12406_));
 sky130_fd_sc_hd__and2_1 _15562_ (.A(_12406_),
    .B(_02411_),
    .X(_03795_));
 sky130_vsdinv _15563_ (.A(\count_cycle[62] ),
    .Y(_12407_));
 sky130_vsdinv _15564_ (.A(\count_cycle[61] ),
    .Y(_12408_));
 sky130_vsdinv _15565_ (.A(\count_cycle[60] ),
    .Y(_12409_));
 sky130_vsdinv _15566_ (.A(\count_cycle[59] ),
    .Y(_12410_));
 sky130_vsdinv _15567_ (.A(\count_cycle[58] ),
    .Y(_12411_));
 sky130_vsdinv _15568_ (.A(\count_cycle[57] ),
    .Y(_12412_));
 sky130_vsdinv _15569_ (.A(\count_cycle[56] ),
    .Y(_12413_));
 sky130_vsdinv _15570_ (.A(\count_cycle[55] ),
    .Y(_12414_));
 sky130_vsdinv _15571_ (.A(\count_cycle[54] ),
    .Y(_12415_));
 sky130_vsdinv _15572_ (.A(\count_cycle[53] ),
    .Y(_12416_));
 sky130_vsdinv _15573_ (.A(\count_cycle[52] ),
    .Y(_12417_));
 sky130_vsdinv _15574_ (.A(\count_cycle[51] ),
    .Y(_12418_));
 sky130_vsdinv _15575_ (.A(\count_cycle[50] ),
    .Y(_12419_));
 sky130_vsdinv _15576_ (.A(\count_cycle[49] ),
    .Y(_12420_));
 sky130_vsdinv _15577_ (.A(\count_cycle[48] ),
    .Y(_12421_));
 sky130_vsdinv _15578_ (.A(\count_cycle[47] ),
    .Y(_12422_));
 sky130_vsdinv _15579_ (.A(\count_cycle[46] ),
    .Y(_12423_));
 sky130_vsdinv _15580_ (.A(\count_cycle[45] ),
    .Y(_12424_));
 sky130_vsdinv _15581_ (.A(\count_cycle[44] ),
    .Y(_12425_));
 sky130_vsdinv _15582_ (.A(\count_cycle[43] ),
    .Y(_12426_));
 sky130_vsdinv _15583_ (.A(\count_cycle[42] ),
    .Y(_12427_));
 sky130_vsdinv _15584_ (.A(\count_cycle[41] ),
    .Y(_12428_));
 sky130_vsdinv _15585_ (.A(\count_cycle[40] ),
    .Y(_12429_));
 sky130_vsdinv _15586_ (.A(\count_cycle[39] ),
    .Y(_12430_));
 sky130_vsdinv _15587_ (.A(\count_cycle[38] ),
    .Y(_12431_));
 sky130_vsdinv _15588_ (.A(\count_cycle[37] ),
    .Y(_12432_));
 sky130_vsdinv _15589_ (.A(\count_cycle[36] ),
    .Y(_12433_));
 sky130_vsdinv _15590_ (.A(\count_cycle[35] ),
    .Y(_12434_));
 sky130_vsdinv _15591_ (.A(\count_cycle[34] ),
    .Y(_12435_));
 sky130_vsdinv _15592_ (.A(\count_cycle[33] ),
    .Y(_12436_));
 sky130_vsdinv _15593_ (.A(\count_cycle[32] ),
    .Y(_12437_));
 sky130_vsdinv _15594_ (.A(\count_cycle[31] ),
    .Y(_02055_));
 sky130_fd_sc_hd__inv_2 _15595_ (.A(\count_cycle[30] ),
    .Y(_02046_));
 sky130_vsdinv _15596_ (.A(\count_cycle[29] ),
    .Y(_02037_));
 sky130_fd_sc_hd__inv_2 _15597_ (.A(\count_cycle[28] ),
    .Y(_02028_));
 sky130_vsdinv _15598_ (.A(\count_cycle[27] ),
    .Y(_02019_));
 sky130_fd_sc_hd__inv_2 _15599_ (.A(\count_cycle[26] ),
    .Y(_02010_));
 sky130_vsdinv _15600_ (.A(\count_cycle[25] ),
    .Y(_02001_));
 sky130_fd_sc_hd__inv_2 _15601_ (.A(\count_cycle[24] ),
    .Y(_01992_));
 sky130_vsdinv _15602_ (.A(\count_cycle[23] ),
    .Y(_01983_));
 sky130_fd_sc_hd__inv_2 _15603_ (.A(\count_cycle[22] ),
    .Y(_01974_));
 sky130_vsdinv _15604_ (.A(\count_cycle[21] ),
    .Y(_01965_));
 sky130_fd_sc_hd__inv_2 _15605_ (.A(\count_cycle[20] ),
    .Y(_01956_));
 sky130_vsdinv _15606_ (.A(\count_cycle[19] ),
    .Y(_01947_));
 sky130_fd_sc_hd__inv_2 _15607_ (.A(\count_cycle[18] ),
    .Y(_01938_));
 sky130_vsdinv _15608_ (.A(\count_cycle[17] ),
    .Y(_01929_));
 sky130_fd_sc_hd__inv_2 _15609_ (.A(\count_cycle[16] ),
    .Y(_01920_));
 sky130_vsdinv _15610_ (.A(\count_cycle[15] ),
    .Y(_01911_));
 sky130_fd_sc_hd__inv_2 _15611_ (.A(\count_cycle[14] ),
    .Y(_01898_));
 sky130_vsdinv _15612_ (.A(\count_cycle[13] ),
    .Y(_01885_));
 sky130_fd_sc_hd__inv_2 _15613_ (.A(\count_cycle[12] ),
    .Y(_01872_));
 sky130_vsdinv _15614_ (.A(\count_cycle[11] ),
    .Y(_01859_));
 sky130_fd_sc_hd__inv_2 _15615_ (.A(\count_cycle[10] ),
    .Y(_01846_));
 sky130_vsdinv _15616_ (.A(\count_cycle[9] ),
    .Y(_01833_));
 sky130_fd_sc_hd__inv_2 _15617_ (.A(\count_cycle[8] ),
    .Y(_01820_));
 sky130_vsdinv _15618_ (.A(\count_cycle[7] ),
    .Y(_01806_));
 sky130_fd_sc_hd__inv_2 _15619_ (.A(\count_cycle[6] ),
    .Y(_01793_));
 sky130_vsdinv _15620_ (.A(\count_cycle[5] ),
    .Y(_01780_));
 sky130_vsdinv _15621_ (.A(\count_cycle[4] ),
    .Y(_01767_));
 sky130_vsdinv _15622_ (.A(\count_cycle[0] ),
    .Y(_12438_));
 sky130_vsdinv _15623_ (.A(\count_cycle[1] ),
    .Y(_12439_));
 sky130_vsdinv _15624_ (.A(\count_cycle[2] ),
    .Y(_12440_));
 sky130_fd_sc_hd__inv_2 _15625_ (.A(\count_cycle[3] ),
    .Y(_01754_));
 sky130_fd_sc_hd__or4_4 _15626_ (.A(_12438_),
    .B(_12439_),
    .C(_12440_),
    .D(_01754_),
    .X(_12441_));
 sky130_fd_sc_hd__or2_1 _15627_ (.A(_01767_),
    .B(_12441_),
    .X(_12442_));
 sky130_fd_sc_hd__or2_1 _15628_ (.A(_01780_),
    .B(_12442_),
    .X(_12443_));
 sky130_fd_sc_hd__or2_1 _15629_ (.A(_01793_),
    .B(_12443_),
    .X(_12444_));
 sky130_fd_sc_hd__or2_1 _15630_ (.A(_01806_),
    .B(_12444_),
    .X(_12445_));
 sky130_fd_sc_hd__or2_1 _15631_ (.A(_01820_),
    .B(_12445_),
    .X(_12446_));
 sky130_fd_sc_hd__or2_2 _15632_ (.A(_01833_),
    .B(_12446_),
    .X(_12447_));
 sky130_fd_sc_hd__or2_1 _15633_ (.A(_01846_),
    .B(_12447_),
    .X(_12448_));
 sky130_fd_sc_hd__or2_1 _15634_ (.A(_01859_),
    .B(_12448_),
    .X(_12449_));
 sky130_fd_sc_hd__or2_1 _15635_ (.A(_01872_),
    .B(_12449_),
    .X(_12450_));
 sky130_fd_sc_hd__or2_2 _15636_ (.A(_01885_),
    .B(_12450_),
    .X(_12451_));
 sky130_fd_sc_hd__or2_1 _15637_ (.A(_01898_),
    .B(_12451_),
    .X(_12452_));
 sky130_fd_sc_hd__or2_2 _15638_ (.A(_01911_),
    .B(_12452_),
    .X(_12453_));
 sky130_fd_sc_hd__or2_1 _15639_ (.A(_01920_),
    .B(_12453_),
    .X(_12454_));
 sky130_fd_sc_hd__or2_2 _15640_ (.A(_01929_),
    .B(_12454_),
    .X(_12455_));
 sky130_fd_sc_hd__or2_1 _15641_ (.A(_01938_),
    .B(_12455_),
    .X(_12456_));
 sky130_fd_sc_hd__or2_2 _15642_ (.A(_01947_),
    .B(_12456_),
    .X(_12457_));
 sky130_fd_sc_hd__or2_1 _15643_ (.A(_01956_),
    .B(_12457_),
    .X(_12458_));
 sky130_fd_sc_hd__or2_2 _15644_ (.A(_01965_),
    .B(_12458_),
    .X(_12459_));
 sky130_fd_sc_hd__or2_1 _15645_ (.A(_01974_),
    .B(_12459_),
    .X(_12460_));
 sky130_fd_sc_hd__or2_2 _15646_ (.A(_01983_),
    .B(_12460_),
    .X(_12461_));
 sky130_fd_sc_hd__or2_1 _15647_ (.A(_01992_),
    .B(_12461_),
    .X(_12462_));
 sky130_fd_sc_hd__or2_2 _15648_ (.A(_02001_),
    .B(_12462_),
    .X(_12463_));
 sky130_fd_sc_hd__or2_1 _15649_ (.A(_02010_),
    .B(_12463_),
    .X(_12464_));
 sky130_fd_sc_hd__or2_2 _15650_ (.A(_02019_),
    .B(_12464_),
    .X(_12465_));
 sky130_fd_sc_hd__or2_1 _15651_ (.A(_02028_),
    .B(_12465_),
    .X(_12466_));
 sky130_fd_sc_hd__or2_1 _15652_ (.A(_02037_),
    .B(_12466_),
    .X(_12467_));
 sky130_fd_sc_hd__or2_1 _15653_ (.A(_02046_),
    .B(_12467_),
    .X(_12468_));
 sky130_fd_sc_hd__or2_1 _15654_ (.A(_02055_),
    .B(_12468_),
    .X(_12469_));
 sky130_fd_sc_hd__or2_1 _15655_ (.A(_12437_),
    .B(_12469_),
    .X(_12470_));
 sky130_fd_sc_hd__or2_1 _15656_ (.A(_12436_),
    .B(_12470_),
    .X(_12471_));
 sky130_fd_sc_hd__or2_1 _15657_ (.A(_12435_),
    .B(_12471_),
    .X(_12472_));
 sky130_fd_sc_hd__or2_2 _15658_ (.A(_12434_),
    .B(_12472_),
    .X(_12473_));
 sky130_fd_sc_hd__or2_1 _15659_ (.A(_12433_),
    .B(_12473_),
    .X(_12474_));
 sky130_fd_sc_hd__or2_2 _15660_ (.A(_12432_),
    .B(_12474_),
    .X(_12475_));
 sky130_fd_sc_hd__or2_1 _15661_ (.A(_12431_),
    .B(_12475_),
    .X(_12476_));
 sky130_fd_sc_hd__or2_2 _15662_ (.A(_12430_),
    .B(_12476_),
    .X(_12477_));
 sky130_fd_sc_hd__or2_1 _15663_ (.A(_12429_),
    .B(_12477_),
    .X(_12478_));
 sky130_fd_sc_hd__or2_2 _15664_ (.A(_12428_),
    .B(_12478_),
    .X(_12479_));
 sky130_fd_sc_hd__or2_1 _15665_ (.A(_12427_),
    .B(_12479_),
    .X(_12480_));
 sky130_fd_sc_hd__or2_2 _15666_ (.A(_12426_),
    .B(_12480_),
    .X(_12481_));
 sky130_fd_sc_hd__or2_1 _15667_ (.A(_12425_),
    .B(_12481_),
    .X(_12482_));
 sky130_fd_sc_hd__or2_1 _15668_ (.A(_12424_),
    .B(_12482_),
    .X(_12483_));
 sky130_fd_sc_hd__or2_1 _15669_ (.A(_12423_),
    .B(_12483_),
    .X(_12484_));
 sky130_fd_sc_hd__or2_2 _15670_ (.A(_12422_),
    .B(_12484_),
    .X(_12485_));
 sky130_fd_sc_hd__or2_1 _15671_ (.A(_12421_),
    .B(_12485_),
    .X(_12486_));
 sky130_fd_sc_hd__or2_2 _15672_ (.A(_12420_),
    .B(_12486_),
    .X(_12487_));
 sky130_fd_sc_hd__or2_1 _15673_ (.A(_12419_),
    .B(_12487_),
    .X(_12488_));
 sky130_fd_sc_hd__or2_2 _15674_ (.A(_12418_),
    .B(_12488_),
    .X(_12489_));
 sky130_fd_sc_hd__or2_1 _15675_ (.A(_12417_),
    .B(_12489_),
    .X(_12490_));
 sky130_fd_sc_hd__or2_1 _15676_ (.A(_12416_),
    .B(_12490_),
    .X(_12491_));
 sky130_fd_sc_hd__or2_1 _15677_ (.A(_12415_),
    .B(_12491_),
    .X(_12492_));
 sky130_fd_sc_hd__or2_2 _15678_ (.A(_12414_),
    .B(_12492_),
    .X(_12493_));
 sky130_fd_sc_hd__or2_1 _15679_ (.A(_12413_),
    .B(_12493_),
    .X(_12494_));
 sky130_fd_sc_hd__or2_2 _15680_ (.A(_12412_),
    .B(_12494_),
    .X(_12495_));
 sky130_fd_sc_hd__or2_1 _15681_ (.A(_12411_),
    .B(_12495_),
    .X(_12496_));
 sky130_fd_sc_hd__or2_2 _15682_ (.A(_12410_),
    .B(_12496_),
    .X(_12497_));
 sky130_fd_sc_hd__or2_1 _15683_ (.A(_12409_),
    .B(_12497_),
    .X(_12498_));
 sky130_fd_sc_hd__or2_2 _15684_ (.A(_12408_),
    .B(_12498_),
    .X(_12499_));
 sky130_fd_sc_hd__or2_1 _15685_ (.A(_12407_),
    .B(_12499_),
    .X(_12500_));
 sky130_vsdinv _15686_ (.A(_12500_),
    .Y(_12501_));
 sky130_vsdinv _15687_ (.A(\count_cycle[63] ),
    .Y(_12502_));
 sky130_fd_sc_hd__o221a_1 _15688_ (.A1(\count_cycle[63] ),
    .A2(_12501_),
    .B1(_12502_),
    .B2(_12500_),
    .C1(_12388_),
    .X(_03794_));
 sky130_fd_sc_hd__a211oi_2 _15689_ (.A1(_12407_),
    .A2(_12499_),
    .B1(_12261_),
    .C1(_12501_),
    .Y(_03793_));
 sky130_vsdinv _15690_ (.A(_12498_),
    .Y(_12503_));
 sky130_fd_sc_hd__o211a_1 _15691_ (.A1(\count_cycle[61] ),
    .A2(_12503_),
    .B1(_12263_),
    .C1(_12499_),
    .X(_03792_));
 sky130_fd_sc_hd__a211oi_2 _15692_ (.A1(_12409_),
    .A2(_12497_),
    .B1(_12261_),
    .C1(_12503_),
    .Y(_03791_));
 sky130_vsdinv _15693_ (.A(_12496_),
    .Y(_12504_));
 sky130_fd_sc_hd__o211a_1 _15694_ (.A1(\count_cycle[59] ),
    .A2(_12504_),
    .B1(_12263_),
    .C1(_12497_),
    .X(_03790_));
 sky130_fd_sc_hd__a211oi_2 _15695_ (.A1(_12411_),
    .A2(_12495_),
    .B1(_12261_),
    .C1(_12504_),
    .Y(_03789_));
 sky130_vsdinv _15696_ (.A(_12494_),
    .Y(_12505_));
 sky130_fd_sc_hd__clkbuf_2 _15697_ (.A(_11787_),
    .X(_12506_));
 sky130_fd_sc_hd__clkbuf_2 _15698_ (.A(_12506_),
    .X(_12507_));
 sky130_fd_sc_hd__o211a_1 _15699_ (.A1(\count_cycle[57] ),
    .A2(_12505_),
    .B1(_12507_),
    .C1(_12495_),
    .X(_03788_));
 sky130_fd_sc_hd__clkbuf_2 _15700_ (.A(_12248_),
    .X(_12508_));
 sky130_fd_sc_hd__a211oi_2 _15701_ (.A1(_12413_),
    .A2(_12493_),
    .B1(_12508_),
    .C1(_12505_),
    .Y(_03787_));
 sky130_vsdinv _15702_ (.A(_12492_),
    .Y(_12509_));
 sky130_fd_sc_hd__o211a_1 _15703_ (.A1(\count_cycle[55] ),
    .A2(_12509_),
    .B1(_12507_),
    .C1(_12493_),
    .X(_03786_));
 sky130_fd_sc_hd__a211oi_1 _15704_ (.A1(_12415_),
    .A2(_12491_),
    .B1(_12508_),
    .C1(_12509_),
    .Y(_03785_));
 sky130_vsdinv _15705_ (.A(_12490_),
    .Y(_12510_));
 sky130_fd_sc_hd__o211a_1 _15706_ (.A1(\count_cycle[53] ),
    .A2(_12510_),
    .B1(_12507_),
    .C1(_12491_),
    .X(_03784_));
 sky130_fd_sc_hd__a211oi_2 _15707_ (.A1(_12417_),
    .A2(_12489_),
    .B1(_12508_),
    .C1(_12510_),
    .Y(_03783_));
 sky130_vsdinv _15708_ (.A(_12488_),
    .Y(_12511_));
 sky130_fd_sc_hd__o211a_1 _15709_ (.A1(\count_cycle[51] ),
    .A2(_12511_),
    .B1(_12507_),
    .C1(_12489_),
    .X(_03782_));
 sky130_fd_sc_hd__a211oi_2 _15710_ (.A1(_12419_),
    .A2(_12487_),
    .B1(_12508_),
    .C1(_12511_),
    .Y(_03781_));
 sky130_vsdinv _15711_ (.A(_12486_),
    .Y(_12512_));
 sky130_fd_sc_hd__clkbuf_2 _15712_ (.A(_12506_),
    .X(_12513_));
 sky130_fd_sc_hd__o211a_1 _15713_ (.A1(\count_cycle[49] ),
    .A2(_12512_),
    .B1(_12513_),
    .C1(_12487_),
    .X(_03780_));
 sky130_fd_sc_hd__clkbuf_2 _15714_ (.A(_11848_),
    .X(_12514_));
 sky130_fd_sc_hd__buf_2 _15715_ (.A(_12514_),
    .X(_12515_));
 sky130_fd_sc_hd__a211oi_2 _15716_ (.A1(_12421_),
    .A2(_12485_),
    .B1(_12515_),
    .C1(_12512_),
    .Y(_03779_));
 sky130_vsdinv _15717_ (.A(_12484_),
    .Y(_12516_));
 sky130_fd_sc_hd__o211a_1 _15718_ (.A1(\count_cycle[47] ),
    .A2(_12516_),
    .B1(_12513_),
    .C1(_12485_),
    .X(_03778_));
 sky130_fd_sc_hd__a211oi_2 _15719_ (.A1(_12423_),
    .A2(_12483_),
    .B1(_12515_),
    .C1(_12516_),
    .Y(_03777_));
 sky130_vsdinv _15720_ (.A(_12482_),
    .Y(_12517_));
 sky130_fd_sc_hd__o211a_1 _15721_ (.A1(\count_cycle[45] ),
    .A2(_12517_),
    .B1(_12513_),
    .C1(_12483_),
    .X(_03776_));
 sky130_fd_sc_hd__a211oi_1 _15722_ (.A1(_12425_),
    .A2(_12481_),
    .B1(_12515_),
    .C1(_12517_),
    .Y(_03775_));
 sky130_vsdinv _15723_ (.A(_12480_),
    .Y(_12518_));
 sky130_fd_sc_hd__o211a_1 _15724_ (.A1(\count_cycle[43] ),
    .A2(_12518_),
    .B1(_12513_),
    .C1(_12481_),
    .X(_03774_));
 sky130_fd_sc_hd__a211oi_2 _15725_ (.A1(_12427_),
    .A2(_12479_),
    .B1(_12515_),
    .C1(_12518_),
    .Y(_03773_));
 sky130_vsdinv _15726_ (.A(_12478_),
    .Y(_12519_));
 sky130_fd_sc_hd__buf_1 _15727_ (.A(_12506_),
    .X(_12520_));
 sky130_fd_sc_hd__o211a_1 _15728_ (.A1(\count_cycle[41] ),
    .A2(_12519_),
    .B1(_12520_),
    .C1(_12479_),
    .X(_03772_));
 sky130_fd_sc_hd__clkbuf_2 _15729_ (.A(_12514_),
    .X(_12521_));
 sky130_fd_sc_hd__a211oi_2 _15730_ (.A1(_12429_),
    .A2(_12477_),
    .B1(_12521_),
    .C1(_12519_),
    .Y(_03771_));
 sky130_vsdinv _15731_ (.A(_12476_),
    .Y(_12522_));
 sky130_fd_sc_hd__o211a_1 _15732_ (.A1(\count_cycle[39] ),
    .A2(_12522_),
    .B1(_12520_),
    .C1(_12477_),
    .X(_03770_));
 sky130_fd_sc_hd__a211oi_2 _15733_ (.A1(_12431_),
    .A2(_12475_),
    .B1(_12521_),
    .C1(_12522_),
    .Y(_03769_));
 sky130_vsdinv _15734_ (.A(_12474_),
    .Y(_12523_));
 sky130_fd_sc_hd__o211a_1 _15735_ (.A1(\count_cycle[37] ),
    .A2(_12523_),
    .B1(_12520_),
    .C1(_12475_),
    .X(_03768_));
 sky130_fd_sc_hd__a211oi_2 _15736_ (.A1(_12433_),
    .A2(_12473_),
    .B1(_12521_),
    .C1(_12523_),
    .Y(_03767_));
 sky130_vsdinv _15737_ (.A(_12472_),
    .Y(_12524_));
 sky130_fd_sc_hd__o211a_1 _15738_ (.A1(\count_cycle[35] ),
    .A2(_12524_),
    .B1(_12520_),
    .C1(_12473_),
    .X(_03766_));
 sky130_fd_sc_hd__a211oi_1 _15739_ (.A1(_12435_),
    .A2(_12471_),
    .B1(_12521_),
    .C1(_12524_),
    .Y(_03765_));
 sky130_vsdinv _15740_ (.A(_12470_),
    .Y(_12525_));
 sky130_fd_sc_hd__clkbuf_2 _15741_ (.A(_12506_),
    .X(_12526_));
 sky130_fd_sc_hd__o211a_1 _15742_ (.A1(\count_cycle[33] ),
    .A2(_12525_),
    .B1(_12526_),
    .C1(_12471_),
    .X(_03764_));
 sky130_fd_sc_hd__clkbuf_2 _15743_ (.A(_12514_),
    .X(_12527_));
 sky130_fd_sc_hd__a211oi_1 _15744_ (.A1(_12437_),
    .A2(_12469_),
    .B1(_12527_),
    .C1(_12525_),
    .Y(_03763_));
 sky130_vsdinv _15745_ (.A(_12468_),
    .Y(_12528_));
 sky130_fd_sc_hd__o211a_1 _15746_ (.A1(\count_cycle[31] ),
    .A2(_12528_),
    .B1(_12526_),
    .C1(_12469_),
    .X(_03762_));
 sky130_fd_sc_hd__a211oi_2 _15747_ (.A1(_02046_),
    .A2(_12467_),
    .B1(_12527_),
    .C1(_12528_),
    .Y(_03761_));
 sky130_vsdinv _15748_ (.A(_12466_),
    .Y(_12529_));
 sky130_fd_sc_hd__o211a_1 _15749_ (.A1(\count_cycle[29] ),
    .A2(_12529_),
    .B1(_12526_),
    .C1(_12467_),
    .X(_03760_));
 sky130_fd_sc_hd__a211oi_2 _15750_ (.A1(_02028_),
    .A2(_12465_),
    .B1(_12527_),
    .C1(_12529_),
    .Y(_03759_));
 sky130_vsdinv _15751_ (.A(_12464_),
    .Y(_12530_));
 sky130_fd_sc_hd__o211a_1 _15752_ (.A1(\count_cycle[27] ),
    .A2(_12530_),
    .B1(_12526_),
    .C1(_12465_),
    .X(_03758_));
 sky130_fd_sc_hd__a211oi_1 _15753_ (.A1(_02010_),
    .A2(_12463_),
    .B1(_12527_),
    .C1(_12530_),
    .Y(_03757_));
 sky130_vsdinv _15754_ (.A(_12462_),
    .Y(_12531_));
 sky130_fd_sc_hd__clkbuf_2 _15755_ (.A(_11788_),
    .X(_12532_));
 sky130_fd_sc_hd__o211a_1 _15756_ (.A1(\count_cycle[25] ),
    .A2(_12531_),
    .B1(_12532_),
    .C1(_12463_),
    .X(_03756_));
 sky130_fd_sc_hd__buf_2 _15757_ (.A(_12514_),
    .X(_12533_));
 sky130_fd_sc_hd__a211oi_2 _15758_ (.A1(_01992_),
    .A2(_12461_),
    .B1(_12533_),
    .C1(_12531_),
    .Y(_03755_));
 sky130_vsdinv _15759_ (.A(_12460_),
    .Y(_12534_));
 sky130_fd_sc_hd__o211a_1 _15760_ (.A1(\count_cycle[23] ),
    .A2(_12534_),
    .B1(_12532_),
    .C1(_12461_),
    .X(_03754_));
 sky130_fd_sc_hd__a211oi_2 _15761_ (.A1(_01974_),
    .A2(_12459_),
    .B1(_12533_),
    .C1(_12534_),
    .Y(_03753_));
 sky130_vsdinv _15762_ (.A(_12458_),
    .Y(_12535_));
 sky130_fd_sc_hd__o211a_1 _15763_ (.A1(\count_cycle[21] ),
    .A2(_12535_),
    .B1(_12532_),
    .C1(_12459_),
    .X(_03752_));
 sky130_fd_sc_hd__a211oi_2 _15764_ (.A1(_01956_),
    .A2(_12457_),
    .B1(_12533_),
    .C1(_12535_),
    .Y(_03751_));
 sky130_vsdinv _15765_ (.A(_12456_),
    .Y(_12536_));
 sky130_fd_sc_hd__o211a_1 _15766_ (.A1(\count_cycle[19] ),
    .A2(_12536_),
    .B1(_12532_),
    .C1(_12457_),
    .X(_03750_));
 sky130_fd_sc_hd__a211oi_2 _15767_ (.A1(_01938_),
    .A2(_12455_),
    .B1(_12533_),
    .C1(_12536_),
    .Y(_03749_));
 sky130_vsdinv _15768_ (.A(_12454_),
    .Y(_12537_));
 sky130_fd_sc_hd__clkbuf_2 _15769_ (.A(_11788_),
    .X(_12538_));
 sky130_fd_sc_hd__o211a_1 _15770_ (.A1(\count_cycle[17] ),
    .A2(_12537_),
    .B1(_12538_),
    .C1(_12455_),
    .X(_03748_));
 sky130_fd_sc_hd__buf_2 _15771_ (.A(_12212_),
    .X(_12539_));
 sky130_fd_sc_hd__a211oi_2 _15772_ (.A1(_01920_),
    .A2(_12453_),
    .B1(_12539_),
    .C1(_12537_),
    .Y(_03747_));
 sky130_vsdinv _15773_ (.A(_12452_),
    .Y(_12540_));
 sky130_fd_sc_hd__o211a_1 _15774_ (.A1(\count_cycle[15] ),
    .A2(_12540_),
    .B1(_12538_),
    .C1(_12453_),
    .X(_03746_));
 sky130_fd_sc_hd__a211oi_2 _15775_ (.A1(_01898_),
    .A2(_12451_),
    .B1(_12539_),
    .C1(_12540_),
    .Y(_03745_));
 sky130_vsdinv _15776_ (.A(_12450_),
    .Y(_12541_));
 sky130_fd_sc_hd__o211a_1 _15777_ (.A1(\count_cycle[13] ),
    .A2(_12541_),
    .B1(_12538_),
    .C1(_12451_),
    .X(_03744_));
 sky130_fd_sc_hd__a211oi_1 _15778_ (.A1(_01872_),
    .A2(_12449_),
    .B1(_12539_),
    .C1(_12541_),
    .Y(_03743_));
 sky130_vsdinv _15779_ (.A(_12448_),
    .Y(_12542_));
 sky130_fd_sc_hd__o211a_1 _15780_ (.A1(\count_cycle[11] ),
    .A2(_12542_),
    .B1(_12538_),
    .C1(_12449_),
    .X(_03742_));
 sky130_fd_sc_hd__a211oi_1 _15781_ (.A1(_01846_),
    .A2(_12447_),
    .B1(_12539_),
    .C1(_12542_),
    .Y(_03741_));
 sky130_vsdinv _15782_ (.A(_12446_),
    .Y(_12543_));
 sky130_fd_sc_hd__buf_1 _15783_ (.A(_11788_),
    .X(_12544_));
 sky130_fd_sc_hd__o211a_1 _15784_ (.A1(\count_cycle[9] ),
    .A2(_12543_),
    .B1(_12544_),
    .C1(_12447_),
    .X(_03740_));
 sky130_fd_sc_hd__clkbuf_2 _15785_ (.A(_12212_),
    .X(_12545_));
 sky130_fd_sc_hd__a211oi_1 _15786_ (.A1(_01820_),
    .A2(_12445_),
    .B1(_12545_),
    .C1(_12543_),
    .Y(_03739_));
 sky130_vsdinv _15787_ (.A(_12444_),
    .Y(_12546_));
 sky130_fd_sc_hd__o211a_1 _15788_ (.A1(\count_cycle[7] ),
    .A2(_12546_),
    .B1(_12544_),
    .C1(_12445_),
    .X(_03738_));
 sky130_fd_sc_hd__a211oi_1 _15789_ (.A1(_01793_),
    .A2(_12443_),
    .B1(_12545_),
    .C1(_12546_),
    .Y(_03737_));
 sky130_vsdinv _15790_ (.A(_12442_),
    .Y(_12547_));
 sky130_fd_sc_hd__o211a_1 _15791_ (.A1(\count_cycle[5] ),
    .A2(_12547_),
    .B1(_12544_),
    .C1(_12443_),
    .X(_03736_));
 sky130_vsdinv _15792_ (.A(_12441_),
    .Y(_12548_));
 sky130_fd_sc_hd__o211a_1 _15793_ (.A1(\count_cycle[4] ),
    .A2(_12548_),
    .B1(_12544_),
    .C1(_12442_),
    .X(_03735_));
 sky130_fd_sc_hd__buf_1 _15794_ (.A(_12440_),
    .X(_01741_));
 sky130_fd_sc_hd__o31a_1 _15795_ (.A1(_12438_),
    .A2(_12439_),
    .A3(_01741_),
    .B1(_01754_),
    .X(_12549_));
 sky130_fd_sc_hd__nor3_1 _15796_ (.A(_12213_),
    .B(_12548_),
    .C(_12549_),
    .Y(_03734_));
 sky130_fd_sc_hd__buf_1 _15797_ (.A(_12438_),
    .X(_02559_));
 sky130_fd_sc_hd__buf_1 _15798_ (.A(_12439_),
    .X(_01728_));
 sky130_fd_sc_hd__o21ai_1 _15799_ (.A1(_02559_),
    .A2(_01728_),
    .B1(_01741_),
    .Y(_12550_));
 sky130_fd_sc_hd__o311a_1 _15800_ (.A1(_02559_),
    .A2(_01728_),
    .A3(_01741_),
    .B1(_11789_),
    .C1(_12550_),
    .X(_03733_));
 sky130_fd_sc_hd__o221a_1 _15801_ (.A1(_02559_),
    .A2(_01728_),
    .B1(\count_cycle[0] ),
    .B2(\count_cycle[1] ),
    .C1(_12388_),
    .X(_03732_));
 sky130_fd_sc_hd__nor2_1 _15802_ (.A(_12393_),
    .B(\count_cycle[0] ),
    .Y(_03731_));
 sky130_vsdinv _15803_ (.A(\cpu_state[0] ),
    .Y(_12551_));
 sky130_fd_sc_hd__nor2_1 _15804_ (.A(_12393_),
    .B(_12551_),
    .Y(_03730_));
 sky130_fd_sc_hd__and2_1 _15805_ (.A(_12406_),
    .B(\pcpi_mul.active[0] ),
    .X(_03729_));
 sky130_fd_sc_hd__buf_1 _15806_ (.A(_11710_),
    .X(_03728_));
 sky130_fd_sc_hd__buf_1 _15807_ (.A(\latched_rd[4] ),
    .X(_12552_));
 sky130_fd_sc_hd__buf_1 _15808_ (.A(\latched_rd[3] ),
    .X(_12553_));
 sky130_fd_sc_hd__buf_1 _15809_ (.A(\latched_rd[2] ),
    .X(_12554_));
 sky130_vsdinv _15810_ (.A(_12554_),
    .Y(_12555_));
 sky130_fd_sc_hd__or3_1 _15811_ (.A(_12552_),
    .B(_12553_),
    .C(_12555_),
    .X(_12556_));
 sky130_fd_sc_hd__buf_2 _15812_ (.A(\latched_rd[0] ),
    .X(_12557_));
 sky130_vsdinv _15813_ (.A(latched_branch),
    .Y(_12558_));
 sky130_vsdinv _15814_ (.A(latched_store),
    .Y(_12559_));
 sky130_fd_sc_hd__and4_1 _15815_ (.A(_11778_),
    .B(_11776_),
    .C(_12558_),
    .D(_12559_),
    .X(_12560_));
 sky130_fd_sc_hd__or3_4 _15816_ (.A(\latched_rd[4] ),
    .B(\latched_rd[3] ),
    .C(\latched_rd[2] ),
    .X(_12561_));
 sky130_fd_sc_hd__nor3_4 _15817_ (.A(\latched_rd[0] ),
    .B(\latched_rd[1] ),
    .C(_12561_),
    .Y(_12562_));
 sky130_fd_sc_hd__or4_4 _15818_ (.A(_11577_),
    .B(_11772_),
    .C(_12560_),
    .D(_12562_),
    .X(_12563_));
 sky130_fd_sc_hd__buf_2 _15819_ (.A(\latched_rd[1] ),
    .X(_12564_));
 sky130_fd_sc_hd__or2b_1 _15820_ (.A(_12563_),
    .B_N(_12564_),
    .X(_12565_));
 sky130_fd_sc_hd__or2_1 _15821_ (.A(_12557_),
    .B(_12565_),
    .X(_12566_));
 sky130_fd_sc_hd__buf_1 _15822_ (.A(_12566_),
    .X(_12567_));
 sky130_fd_sc_hd__or2_2 _15823_ (.A(_12556_),
    .B(_12567_),
    .X(_12568_));
 sky130_fd_sc_hd__clkbuf_4 _15824_ (.A(_12568_),
    .X(_12569_));
 sky130_fd_sc_hd__buf_1 _15825_ (.A(_12569_),
    .X(_12570_));
 sky130_fd_sc_hd__clkbuf_2 _15826_ (.A(\cpuregs_wrdata[31] ),
    .X(_12571_));
 sky130_fd_sc_hd__buf_1 _15827_ (.A(_12571_),
    .X(_12572_));
 sky130_vsdinv _15828_ (.A(_12568_),
    .Y(_12573_));
 sky130_fd_sc_hd__clkbuf_4 _15829_ (.A(_12573_),
    .X(_12574_));
 sky130_fd_sc_hd__buf_1 _15830_ (.A(_12574_),
    .X(_12575_));
 sky130_fd_sc_hd__a22o_1 _15831_ (.A1(\cpuregs[6][31] ),
    .A2(_12570_),
    .B1(_12572_),
    .B2(_12575_),
    .X(_03727_));
 sky130_fd_sc_hd__clkbuf_2 _15832_ (.A(\cpuregs_wrdata[30] ),
    .X(_12576_));
 sky130_fd_sc_hd__buf_1 _15833_ (.A(_12576_),
    .X(_12577_));
 sky130_fd_sc_hd__a22o_1 _15834_ (.A1(\cpuregs[6][30] ),
    .A2(_12570_),
    .B1(_12577_),
    .B2(_12575_),
    .X(_03726_));
 sky130_fd_sc_hd__clkbuf_2 _15835_ (.A(\cpuregs_wrdata[29] ),
    .X(_12578_));
 sky130_fd_sc_hd__buf_1 _15836_ (.A(_12578_),
    .X(_12579_));
 sky130_fd_sc_hd__a22o_1 _15837_ (.A1(\cpuregs[6][29] ),
    .A2(_12570_),
    .B1(_12579_),
    .B2(_12575_),
    .X(_03725_));
 sky130_fd_sc_hd__clkbuf_2 _15838_ (.A(\cpuregs_wrdata[28] ),
    .X(_12580_));
 sky130_fd_sc_hd__buf_1 _15839_ (.A(_12580_),
    .X(_12581_));
 sky130_fd_sc_hd__a22o_1 _15840_ (.A1(\cpuregs[6][28] ),
    .A2(_12570_),
    .B1(_12581_),
    .B2(_12575_),
    .X(_03724_));
 sky130_fd_sc_hd__buf_1 _15841_ (.A(_12569_),
    .X(_12582_));
 sky130_fd_sc_hd__clkbuf_2 _15842_ (.A(\cpuregs_wrdata[27] ),
    .X(_12583_));
 sky130_fd_sc_hd__clkbuf_2 _15843_ (.A(_12583_),
    .X(_12584_));
 sky130_fd_sc_hd__buf_1 _15844_ (.A(_12574_),
    .X(_12585_));
 sky130_fd_sc_hd__a22o_1 _15845_ (.A1(\cpuregs[6][27] ),
    .A2(_12582_),
    .B1(_12584_),
    .B2(_12585_),
    .X(_03723_));
 sky130_fd_sc_hd__clkbuf_2 _15846_ (.A(\cpuregs_wrdata[26] ),
    .X(_12586_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _15847_ (.A(_12586_),
    .X(_12587_));
 sky130_fd_sc_hd__a22o_1 _15848_ (.A1(\cpuregs[6][26] ),
    .A2(_12582_),
    .B1(_12587_),
    .B2(_12585_),
    .X(_03722_));
 sky130_fd_sc_hd__clkbuf_2 _15849_ (.A(\cpuregs_wrdata[25] ),
    .X(_12588_));
 sky130_fd_sc_hd__clkbuf_2 _15850_ (.A(_12588_),
    .X(_12589_));
 sky130_fd_sc_hd__a22o_1 _15851_ (.A1(\cpuregs[6][25] ),
    .A2(_12582_),
    .B1(_12589_),
    .B2(_12585_),
    .X(_03721_));
 sky130_fd_sc_hd__clkbuf_2 _15852_ (.A(\cpuregs_wrdata[24] ),
    .X(_12590_));
 sky130_fd_sc_hd__buf_1 _15853_ (.A(_12590_),
    .X(_12591_));
 sky130_fd_sc_hd__a22o_1 _15854_ (.A1(\cpuregs[6][24] ),
    .A2(_12582_),
    .B1(_12591_),
    .B2(_12585_),
    .X(_03720_));
 sky130_fd_sc_hd__buf_1 _15855_ (.A(_12569_),
    .X(_12592_));
 sky130_fd_sc_hd__buf_1 _15856_ (.A(\cpuregs_wrdata[23] ),
    .X(_12593_));
 sky130_fd_sc_hd__clkbuf_2 _15857_ (.A(_12593_),
    .X(_12594_));
 sky130_fd_sc_hd__buf_1 _15858_ (.A(_12574_),
    .X(_12595_));
 sky130_fd_sc_hd__a22o_1 _15859_ (.A1(\cpuregs[6][23] ),
    .A2(_12592_),
    .B1(_12594_),
    .B2(_12595_),
    .X(_03719_));
 sky130_fd_sc_hd__buf_1 _15860_ (.A(\cpuregs_wrdata[22] ),
    .X(_12596_));
 sky130_fd_sc_hd__clkbuf_2 _15861_ (.A(_12596_),
    .X(_12597_));
 sky130_fd_sc_hd__a22o_1 _15862_ (.A1(\cpuregs[6][22] ),
    .A2(_12592_),
    .B1(_12597_),
    .B2(_12595_),
    .X(_03718_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _15863_ (.A(\cpuregs_wrdata[21] ),
    .X(_12598_));
 sky130_fd_sc_hd__clkbuf_2 _15864_ (.A(_12598_),
    .X(_12599_));
 sky130_fd_sc_hd__a22o_1 _15865_ (.A1(\cpuregs[6][21] ),
    .A2(_12592_),
    .B1(_12599_),
    .B2(_12595_),
    .X(_03717_));
 sky130_fd_sc_hd__clkbuf_2 _15866_ (.A(\cpuregs_wrdata[20] ),
    .X(_12600_));
 sky130_fd_sc_hd__clkbuf_2 _15867_ (.A(_12600_),
    .X(_12601_));
 sky130_fd_sc_hd__a22o_1 _15868_ (.A1(\cpuregs[6][20] ),
    .A2(_12592_),
    .B1(_12601_),
    .B2(_12595_),
    .X(_03716_));
 sky130_fd_sc_hd__buf_1 _15869_ (.A(_12569_),
    .X(_12602_));
 sky130_fd_sc_hd__clkbuf_2 _15870_ (.A(\cpuregs_wrdata[19] ),
    .X(_12603_));
 sky130_fd_sc_hd__clkbuf_2 _15871_ (.A(_12603_),
    .X(_12604_));
 sky130_fd_sc_hd__buf_1 _15872_ (.A(_12574_),
    .X(_12605_));
 sky130_fd_sc_hd__a22o_1 _15873_ (.A1(\cpuregs[6][19] ),
    .A2(_12602_),
    .B1(_12604_),
    .B2(_12605_),
    .X(_03715_));
 sky130_fd_sc_hd__clkbuf_2 _15874_ (.A(\cpuregs_wrdata[18] ),
    .X(_12606_));
 sky130_fd_sc_hd__clkbuf_2 _15875_ (.A(_12606_),
    .X(_12607_));
 sky130_fd_sc_hd__a22o_1 _15876_ (.A1(\cpuregs[6][18] ),
    .A2(_12602_),
    .B1(_12607_),
    .B2(_12605_),
    .X(_03714_));
 sky130_fd_sc_hd__clkbuf_2 _15877_ (.A(\cpuregs_wrdata[17] ),
    .X(_12608_));
 sky130_fd_sc_hd__clkbuf_2 _15878_ (.A(_12608_),
    .X(_12609_));
 sky130_fd_sc_hd__a22o_1 _15879_ (.A1(\cpuregs[6][17] ),
    .A2(_12602_),
    .B1(_12609_),
    .B2(_12605_),
    .X(_03713_));
 sky130_fd_sc_hd__clkbuf_2 _15880_ (.A(\cpuregs_wrdata[16] ),
    .X(_12610_));
 sky130_fd_sc_hd__clkbuf_2 _15881_ (.A(_12610_),
    .X(_12611_));
 sky130_fd_sc_hd__a22o_1 _15882_ (.A1(\cpuregs[6][16] ),
    .A2(_12602_),
    .B1(_12611_),
    .B2(_12605_),
    .X(_03712_));
 sky130_fd_sc_hd__clkbuf_2 _15883_ (.A(_12568_),
    .X(_12612_));
 sky130_fd_sc_hd__buf_1 _15884_ (.A(_12612_),
    .X(_12613_));
 sky130_fd_sc_hd__clkbuf_2 _15885_ (.A(\cpuregs_wrdata[15] ),
    .X(_12614_));
 sky130_fd_sc_hd__buf_1 _15886_ (.A(_12614_),
    .X(_12615_));
 sky130_fd_sc_hd__clkbuf_2 _15887_ (.A(_12573_),
    .X(_12616_));
 sky130_fd_sc_hd__buf_1 _15888_ (.A(_12616_),
    .X(_12617_));
 sky130_fd_sc_hd__a22o_1 _15889_ (.A1(\cpuregs[6][15] ),
    .A2(_12613_),
    .B1(_12615_),
    .B2(_12617_),
    .X(_03711_));
 sky130_fd_sc_hd__clkbuf_2 _15890_ (.A(\cpuregs_wrdata[14] ),
    .X(_12618_));
 sky130_fd_sc_hd__clkbuf_2 _15891_ (.A(_12618_),
    .X(_12619_));
 sky130_fd_sc_hd__a22o_1 _15892_ (.A1(\cpuregs[6][14] ),
    .A2(_12613_),
    .B1(_12619_),
    .B2(_12617_),
    .X(_03710_));
 sky130_fd_sc_hd__clkbuf_2 _15893_ (.A(\cpuregs_wrdata[13] ),
    .X(_12620_));
 sky130_fd_sc_hd__clkbuf_2 _15894_ (.A(_12620_),
    .X(_12621_));
 sky130_fd_sc_hd__a22o_1 _15895_ (.A1(\cpuregs[6][13] ),
    .A2(_12613_),
    .B1(_12621_),
    .B2(_12617_),
    .X(_03709_));
 sky130_fd_sc_hd__clkbuf_2 _15896_ (.A(\cpuregs_wrdata[12] ),
    .X(_12622_));
 sky130_fd_sc_hd__clkbuf_2 _15897_ (.A(_12622_),
    .X(_12623_));
 sky130_fd_sc_hd__a22o_1 _15898_ (.A1(\cpuregs[6][12] ),
    .A2(_12613_),
    .B1(_12623_),
    .B2(_12617_),
    .X(_03708_));
 sky130_fd_sc_hd__buf_1 _15899_ (.A(_12612_),
    .X(_12624_));
 sky130_fd_sc_hd__clkbuf_2 _15900_ (.A(\cpuregs_wrdata[11] ),
    .X(_12625_));
 sky130_fd_sc_hd__buf_1 _15901_ (.A(_12625_),
    .X(_12626_));
 sky130_fd_sc_hd__buf_1 _15902_ (.A(_12616_),
    .X(_12627_));
 sky130_fd_sc_hd__a22o_1 _15903_ (.A1(\cpuregs[6][11] ),
    .A2(_12624_),
    .B1(_12626_),
    .B2(_12627_),
    .X(_03707_));
 sky130_fd_sc_hd__clkbuf_2 _15904_ (.A(\cpuregs_wrdata[10] ),
    .X(_12628_));
 sky130_fd_sc_hd__buf_1 _15905_ (.A(_12628_),
    .X(_12629_));
 sky130_fd_sc_hd__a22o_1 _15906_ (.A1(\cpuregs[6][10] ),
    .A2(_12624_),
    .B1(_12629_),
    .B2(_12627_),
    .X(_03706_));
 sky130_fd_sc_hd__clkbuf_2 _15907_ (.A(\cpuregs_wrdata[9] ),
    .X(_12630_));
 sky130_fd_sc_hd__buf_1 _15908_ (.A(_12630_),
    .X(_12631_));
 sky130_fd_sc_hd__a22o_1 _15909_ (.A1(\cpuregs[6][9] ),
    .A2(_12624_),
    .B1(_12631_),
    .B2(_12627_),
    .X(_03705_));
 sky130_fd_sc_hd__clkbuf_2 _15910_ (.A(\cpuregs_wrdata[8] ),
    .X(_12632_));
 sky130_fd_sc_hd__buf_1 _15911_ (.A(_12632_),
    .X(_12633_));
 sky130_fd_sc_hd__a22o_1 _15912_ (.A1(\cpuregs[6][8] ),
    .A2(_12624_),
    .B1(_12633_),
    .B2(_12627_),
    .X(_03704_));
 sky130_fd_sc_hd__buf_1 _15913_ (.A(_12612_),
    .X(_12634_));
 sky130_fd_sc_hd__buf_2 _15914_ (.A(\cpuregs_wrdata[7] ),
    .X(_12635_));
 sky130_fd_sc_hd__clkbuf_2 _15915_ (.A(_12635_),
    .X(_12636_));
 sky130_fd_sc_hd__buf_1 _15916_ (.A(_12616_),
    .X(_12637_));
 sky130_fd_sc_hd__a22o_1 _15917_ (.A1(\cpuregs[6][7] ),
    .A2(_12634_),
    .B1(_12636_),
    .B2(_12637_),
    .X(_03703_));
 sky130_fd_sc_hd__clkbuf_2 _15918_ (.A(\cpuregs_wrdata[6] ),
    .X(_12638_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _15919_ (.A(_12638_),
    .X(_12639_));
 sky130_fd_sc_hd__a22o_1 _15920_ (.A1(\cpuregs[6][6] ),
    .A2(_12634_),
    .B1(_12639_),
    .B2(_12637_),
    .X(_03702_));
 sky130_fd_sc_hd__clkbuf_2 _15921_ (.A(\cpuregs_wrdata[5] ),
    .X(_12640_));
 sky130_fd_sc_hd__clkbuf_2 _15922_ (.A(_12640_),
    .X(_12641_));
 sky130_fd_sc_hd__a22o_1 _15923_ (.A1(\cpuregs[6][5] ),
    .A2(_12634_),
    .B1(_12641_),
    .B2(_12637_),
    .X(_03701_));
 sky130_fd_sc_hd__buf_2 _15924_ (.A(\cpuregs_wrdata[4] ),
    .X(_12642_));
 sky130_fd_sc_hd__clkbuf_2 _15925_ (.A(_12642_),
    .X(_12643_));
 sky130_fd_sc_hd__a22o_1 _15926_ (.A1(\cpuregs[6][4] ),
    .A2(_12634_),
    .B1(_12643_),
    .B2(_12637_),
    .X(_03700_));
 sky130_fd_sc_hd__buf_1 _15927_ (.A(_12612_),
    .X(_12644_));
 sky130_fd_sc_hd__clkbuf_2 _15928_ (.A(\cpuregs_wrdata[3] ),
    .X(_12645_));
 sky130_fd_sc_hd__clkbuf_2 _15929_ (.A(_12645_),
    .X(_12646_));
 sky130_fd_sc_hd__buf_1 _15930_ (.A(_12616_),
    .X(_12647_));
 sky130_fd_sc_hd__a22o_1 _15931_ (.A1(\cpuregs[6][3] ),
    .A2(_12644_),
    .B1(_12646_),
    .B2(_12647_),
    .X(_03699_));
 sky130_fd_sc_hd__clkbuf_2 _15932_ (.A(\cpuregs_wrdata[2] ),
    .X(_12648_));
 sky130_fd_sc_hd__clkbuf_2 _15933_ (.A(_12648_),
    .X(_12649_));
 sky130_fd_sc_hd__a22o_1 _15934_ (.A1(\cpuregs[6][2] ),
    .A2(_12644_),
    .B1(_12649_),
    .B2(_12647_),
    .X(_03698_));
 sky130_fd_sc_hd__clkbuf_2 _15935_ (.A(\cpuregs_wrdata[1] ),
    .X(_12650_));
 sky130_fd_sc_hd__clkbuf_2 _15936_ (.A(_12650_),
    .X(_12651_));
 sky130_fd_sc_hd__a22o_1 _15937_ (.A1(\cpuregs[6][1] ),
    .A2(_12644_),
    .B1(_12651_),
    .B2(_12647_),
    .X(_03697_));
 sky130_fd_sc_hd__clkbuf_2 _15938_ (.A(\cpuregs_wrdata[0] ),
    .X(_12652_));
 sky130_fd_sc_hd__clkbuf_2 _15939_ (.A(_12652_),
    .X(_12653_));
 sky130_fd_sc_hd__a22o_1 _15940_ (.A1(\cpuregs[6][0] ),
    .A2(_12644_),
    .B1(_12653_),
    .B2(_12647_),
    .X(_03696_));
 sky130_vsdinv _15941_ (.A(_12553_),
    .Y(_12654_));
 sky130_fd_sc_hd__or3_4 _15942_ (.A(\latched_rd[4] ),
    .B(_12654_),
    .C(_12554_),
    .X(_12655_));
 sky130_vsdinv _15943_ (.A(_12557_),
    .Y(_12656_));
 sky130_fd_sc_hd__or3_1 _15944_ (.A(_12656_),
    .B(_12564_),
    .C(_12563_),
    .X(_12657_));
 sky130_fd_sc_hd__buf_1 _15945_ (.A(_12657_),
    .X(_12658_));
 sky130_fd_sc_hd__or2_2 _15946_ (.A(_12655_),
    .B(_12658_),
    .X(_12659_));
 sky130_fd_sc_hd__clkbuf_4 _15947_ (.A(_12659_),
    .X(_12660_));
 sky130_fd_sc_hd__buf_1 _15948_ (.A(_12660_),
    .X(_12661_));
 sky130_vsdinv _15949_ (.A(_12659_),
    .Y(_12662_));
 sky130_fd_sc_hd__clkbuf_4 _15950_ (.A(_12662_),
    .X(_12663_));
 sky130_fd_sc_hd__buf_1 _15951_ (.A(_12663_),
    .X(_12664_));
 sky130_fd_sc_hd__a22o_1 _15952_ (.A1(\cpuregs[9][31] ),
    .A2(_12661_),
    .B1(_12572_),
    .B2(_12664_),
    .X(_03695_));
 sky130_fd_sc_hd__a22o_1 _15953_ (.A1(\cpuregs[9][30] ),
    .A2(_12661_),
    .B1(_12577_),
    .B2(_12664_),
    .X(_03694_));
 sky130_fd_sc_hd__a22o_1 _15954_ (.A1(\cpuregs[9][29] ),
    .A2(_12661_),
    .B1(_12579_),
    .B2(_12664_),
    .X(_03693_));
 sky130_fd_sc_hd__a22o_1 _15955_ (.A1(\cpuregs[9][28] ),
    .A2(_12661_),
    .B1(_12581_),
    .B2(_12664_),
    .X(_03692_));
 sky130_fd_sc_hd__buf_1 _15956_ (.A(_12660_),
    .X(_12665_));
 sky130_fd_sc_hd__buf_1 _15957_ (.A(_12663_),
    .X(_12666_));
 sky130_fd_sc_hd__a22o_1 _15958_ (.A1(\cpuregs[9][27] ),
    .A2(_12665_),
    .B1(_12584_),
    .B2(_12666_),
    .X(_03691_));
 sky130_fd_sc_hd__a22o_1 _15959_ (.A1(\cpuregs[9][26] ),
    .A2(_12665_),
    .B1(_12587_),
    .B2(_12666_),
    .X(_03690_));
 sky130_fd_sc_hd__a22o_1 _15960_ (.A1(\cpuregs[9][25] ),
    .A2(_12665_),
    .B1(_12589_),
    .B2(_12666_),
    .X(_03689_));
 sky130_fd_sc_hd__a22o_1 _15961_ (.A1(\cpuregs[9][24] ),
    .A2(_12665_),
    .B1(_12591_),
    .B2(_12666_),
    .X(_03688_));
 sky130_fd_sc_hd__buf_1 _15962_ (.A(_12660_),
    .X(_12667_));
 sky130_fd_sc_hd__buf_1 _15963_ (.A(_12663_),
    .X(_12668_));
 sky130_fd_sc_hd__a22o_1 _15964_ (.A1(\cpuregs[9][23] ),
    .A2(_12667_),
    .B1(_12594_),
    .B2(_12668_),
    .X(_03687_));
 sky130_fd_sc_hd__a22o_1 _15965_ (.A1(\cpuregs[9][22] ),
    .A2(_12667_),
    .B1(_12597_),
    .B2(_12668_),
    .X(_03686_));
 sky130_fd_sc_hd__a22o_1 _15966_ (.A1(\cpuregs[9][21] ),
    .A2(_12667_),
    .B1(_12599_),
    .B2(_12668_),
    .X(_03685_));
 sky130_fd_sc_hd__a22o_1 _15967_ (.A1(\cpuregs[9][20] ),
    .A2(_12667_),
    .B1(_12601_),
    .B2(_12668_),
    .X(_03684_));
 sky130_fd_sc_hd__buf_1 _15968_ (.A(_12660_),
    .X(_12669_));
 sky130_fd_sc_hd__buf_1 _15969_ (.A(_12663_),
    .X(_12670_));
 sky130_fd_sc_hd__a22o_1 _15970_ (.A1(\cpuregs[9][19] ),
    .A2(_12669_),
    .B1(_12604_),
    .B2(_12670_),
    .X(_03683_));
 sky130_fd_sc_hd__a22o_1 _15971_ (.A1(\cpuregs[9][18] ),
    .A2(_12669_),
    .B1(_12607_),
    .B2(_12670_),
    .X(_03682_));
 sky130_fd_sc_hd__a22o_1 _15972_ (.A1(\cpuregs[9][17] ),
    .A2(_12669_),
    .B1(_12609_),
    .B2(_12670_),
    .X(_03681_));
 sky130_fd_sc_hd__a22o_1 _15973_ (.A1(\cpuregs[9][16] ),
    .A2(_12669_),
    .B1(_12611_),
    .B2(_12670_),
    .X(_03680_));
 sky130_fd_sc_hd__clkbuf_2 _15974_ (.A(_12659_),
    .X(_12671_));
 sky130_fd_sc_hd__buf_1 _15975_ (.A(_12671_),
    .X(_12672_));
 sky130_fd_sc_hd__clkbuf_2 _15976_ (.A(_12662_),
    .X(_12673_));
 sky130_fd_sc_hd__buf_1 _15977_ (.A(_12673_),
    .X(_12674_));
 sky130_fd_sc_hd__a22o_1 _15978_ (.A1(\cpuregs[9][15] ),
    .A2(_12672_),
    .B1(_12615_),
    .B2(_12674_),
    .X(_03679_));
 sky130_fd_sc_hd__a22o_1 _15979_ (.A1(\cpuregs[9][14] ),
    .A2(_12672_),
    .B1(_12619_),
    .B2(_12674_),
    .X(_03678_));
 sky130_fd_sc_hd__a22o_1 _15980_ (.A1(\cpuregs[9][13] ),
    .A2(_12672_),
    .B1(_12621_),
    .B2(_12674_),
    .X(_03677_));
 sky130_fd_sc_hd__a22o_1 _15981_ (.A1(\cpuregs[9][12] ),
    .A2(_12672_),
    .B1(_12623_),
    .B2(_12674_),
    .X(_03676_));
 sky130_fd_sc_hd__buf_1 _15982_ (.A(_12671_),
    .X(_12675_));
 sky130_fd_sc_hd__buf_1 _15983_ (.A(_12673_),
    .X(_12676_));
 sky130_fd_sc_hd__a22o_1 _15984_ (.A1(\cpuregs[9][11] ),
    .A2(_12675_),
    .B1(_12626_),
    .B2(_12676_),
    .X(_03675_));
 sky130_fd_sc_hd__a22o_1 _15985_ (.A1(\cpuregs[9][10] ),
    .A2(_12675_),
    .B1(_12629_),
    .B2(_12676_),
    .X(_03674_));
 sky130_fd_sc_hd__a22o_1 _15986_ (.A1(\cpuregs[9][9] ),
    .A2(_12675_),
    .B1(_12631_),
    .B2(_12676_),
    .X(_03673_));
 sky130_fd_sc_hd__a22o_1 _15987_ (.A1(\cpuregs[9][8] ),
    .A2(_12675_),
    .B1(_12633_),
    .B2(_12676_),
    .X(_03672_));
 sky130_fd_sc_hd__buf_1 _15988_ (.A(_12671_),
    .X(_12677_));
 sky130_fd_sc_hd__buf_1 _15989_ (.A(_12673_),
    .X(_12678_));
 sky130_fd_sc_hd__a22o_1 _15990_ (.A1(\cpuregs[9][7] ),
    .A2(_12677_),
    .B1(_12636_),
    .B2(_12678_),
    .X(_03671_));
 sky130_fd_sc_hd__a22o_1 _15991_ (.A1(\cpuregs[9][6] ),
    .A2(_12677_),
    .B1(_12639_),
    .B2(_12678_),
    .X(_03670_));
 sky130_fd_sc_hd__a22o_1 _15992_ (.A1(\cpuregs[9][5] ),
    .A2(_12677_),
    .B1(_12641_),
    .B2(_12678_),
    .X(_03669_));
 sky130_fd_sc_hd__a22o_1 _15993_ (.A1(\cpuregs[9][4] ),
    .A2(_12677_),
    .B1(_12643_),
    .B2(_12678_),
    .X(_03668_));
 sky130_fd_sc_hd__buf_1 _15994_ (.A(_12671_),
    .X(_12679_));
 sky130_fd_sc_hd__buf_1 _15995_ (.A(_12673_),
    .X(_12680_));
 sky130_fd_sc_hd__a22o_1 _15996_ (.A1(\cpuregs[9][3] ),
    .A2(_12679_),
    .B1(_12646_),
    .B2(_12680_),
    .X(_03667_));
 sky130_fd_sc_hd__a22o_1 _15997_ (.A1(\cpuregs[9][2] ),
    .A2(_12679_),
    .B1(_12649_),
    .B2(_12680_),
    .X(_03666_));
 sky130_fd_sc_hd__a22o_1 _15998_ (.A1(\cpuregs[9][1] ),
    .A2(_12679_),
    .B1(_12651_),
    .B2(_12680_),
    .X(_03665_));
 sky130_fd_sc_hd__a22o_1 _15999_ (.A1(\cpuregs[9][0] ),
    .A2(_12679_),
    .B1(_12653_),
    .B2(_12680_),
    .X(_03664_));
 sky130_fd_sc_hd__o21ai_4 _16000_ (.A1(_11739_),
    .A2(_12365_),
    .B1(_11543_),
    .Y(_12681_));
 sky130_fd_sc_hd__clkbuf_4 _16001_ (.A(_12681_),
    .X(_12682_));
 sky130_vsdinv _16002_ (.A(_12681_),
    .Y(_12683_));
 sky130_fd_sc_hd__buf_2 _16003_ (.A(_12683_),
    .X(_12684_));
 sky130_fd_sc_hd__clkbuf_2 _16004_ (.A(_12684_),
    .X(_12685_));
 sky130_fd_sc_hd__a22o_1 _16005_ (.A1(_11712_),
    .A2(_12682_),
    .B1(_02467_),
    .B2(_12685_),
    .X(_03663_));
 sky130_fd_sc_hd__clkbuf_4 _16006_ (.A(net361),
    .X(_12686_));
 sky130_fd_sc_hd__a22o_1 _16007_ (.A1(_12686_),
    .A2(_12682_),
    .B1(_02466_),
    .B2(_12685_),
    .X(_03662_));
 sky130_fd_sc_hd__buf_2 _16008_ (.A(net359),
    .X(_12687_));
 sky130_fd_sc_hd__a22o_1 _16009_ (.A1(_12687_),
    .A2(_12682_),
    .B1(_02464_),
    .B2(_12685_),
    .X(_03661_));
 sky130_fd_sc_hd__clkbuf_4 _16010_ (.A(net358),
    .X(_12688_));
 sky130_fd_sc_hd__buf_2 _16011_ (.A(_12681_),
    .X(_12689_));
 sky130_fd_sc_hd__buf_1 _16012_ (.A(_12689_),
    .X(_12690_));
 sky130_fd_sc_hd__a22o_1 _16013_ (.A1(_12688_),
    .A2(_12690_),
    .B1(_02463_),
    .B2(_12685_),
    .X(_03660_));
 sky130_fd_sc_hd__buf_2 _16014_ (.A(net357),
    .X(_12691_));
 sky130_fd_sc_hd__buf_1 _16015_ (.A(_12684_),
    .X(_12692_));
 sky130_fd_sc_hd__a22o_1 _16016_ (.A1(_12691_),
    .A2(_12690_),
    .B1(_02462_),
    .B2(_12692_),
    .X(_03659_));
 sky130_fd_sc_hd__clkbuf_4 _16017_ (.A(net356),
    .X(_12693_));
 sky130_fd_sc_hd__a22o_1 _16018_ (.A1(_12693_),
    .A2(_12690_),
    .B1(_02461_),
    .B2(_12692_),
    .X(_03658_));
 sky130_fd_sc_hd__clkbuf_4 _16019_ (.A(net355),
    .X(_12694_));
 sky130_fd_sc_hd__a22o_1 _16020_ (.A1(_12694_),
    .A2(_12690_),
    .B1(_02460_),
    .B2(_12692_),
    .X(_03657_));
 sky130_fd_sc_hd__clkbuf_4 _16021_ (.A(net354),
    .X(_12695_));
 sky130_fd_sc_hd__buf_1 _16022_ (.A(_12689_),
    .X(_12696_));
 sky130_fd_sc_hd__a22o_1 _16023_ (.A1(_12695_),
    .A2(_12696_),
    .B1(_02459_),
    .B2(_12692_),
    .X(_03656_));
 sky130_fd_sc_hd__clkbuf_4 _16024_ (.A(net353),
    .X(_12697_));
 sky130_fd_sc_hd__buf_1 _16025_ (.A(_12684_),
    .X(_12698_));
 sky130_fd_sc_hd__a22o_1 _16026_ (.A1(_12697_),
    .A2(_12696_),
    .B1(_02458_),
    .B2(_12698_),
    .X(_03655_));
 sky130_fd_sc_hd__buf_4 _16027_ (.A(net352),
    .X(_12699_));
 sky130_fd_sc_hd__a22o_1 _16028_ (.A1(_12699_),
    .A2(_12696_),
    .B1(_02457_),
    .B2(_12698_),
    .X(_03654_));
 sky130_fd_sc_hd__clkbuf_4 _16029_ (.A(net351),
    .X(_12700_));
 sky130_fd_sc_hd__a22o_1 _16030_ (.A1(_12700_),
    .A2(_12696_),
    .B1(_02456_),
    .B2(_12698_),
    .X(_03653_));
 sky130_fd_sc_hd__buf_4 _16031_ (.A(net350),
    .X(_12701_));
 sky130_fd_sc_hd__clkbuf_2 _16032_ (.A(_12689_),
    .X(_12702_));
 sky130_fd_sc_hd__a22o_1 _16033_ (.A1(_12701_),
    .A2(_12702_),
    .B1(_02455_),
    .B2(_12698_),
    .X(_03652_));
 sky130_fd_sc_hd__buf_4 _16034_ (.A(net348),
    .X(_12703_));
 sky130_fd_sc_hd__buf_1 _16035_ (.A(_12684_),
    .X(_12704_));
 sky130_fd_sc_hd__a22o_1 _16036_ (.A1(_12703_),
    .A2(_12702_),
    .B1(_02453_),
    .B2(_12704_),
    .X(_03651_));
 sky130_fd_sc_hd__buf_4 _16037_ (.A(net347),
    .X(_12705_));
 sky130_fd_sc_hd__a22o_1 _16038_ (.A1(_12705_),
    .A2(_12702_),
    .B1(_02452_),
    .B2(_12704_),
    .X(_03650_));
 sky130_fd_sc_hd__clkbuf_4 _16039_ (.A(net346),
    .X(_12706_));
 sky130_fd_sc_hd__a22o_1 _16040_ (.A1(_12706_),
    .A2(_12702_),
    .B1(_02451_),
    .B2(_12704_),
    .X(_03649_));
 sky130_fd_sc_hd__clkbuf_4 _16041_ (.A(net345),
    .X(_12707_));
 sky130_fd_sc_hd__clkbuf_2 _16042_ (.A(_12681_),
    .X(_12708_));
 sky130_fd_sc_hd__clkbuf_2 _16043_ (.A(_12708_),
    .X(_12709_));
 sky130_fd_sc_hd__a22o_1 _16044_ (.A1(_12707_),
    .A2(_12709_),
    .B1(_02450_),
    .B2(_12704_),
    .X(_03648_));
 sky130_fd_sc_hd__clkbuf_2 _16045_ (.A(net344),
    .X(_12710_));
 sky130_fd_sc_hd__clkbuf_4 _16046_ (.A(_12710_),
    .X(_12711_));
 sky130_fd_sc_hd__clkbuf_2 _16047_ (.A(_12683_),
    .X(_12712_));
 sky130_fd_sc_hd__buf_1 _16048_ (.A(_12712_),
    .X(_12713_));
 sky130_fd_sc_hd__a22o_1 _16049_ (.A1(_12711_),
    .A2(_12709_),
    .B1(_02449_),
    .B2(_12713_),
    .X(_03647_));
 sky130_fd_sc_hd__clkbuf_4 _16050_ (.A(net343),
    .X(_12714_));
 sky130_fd_sc_hd__a22o_1 _16051_ (.A1(_12714_),
    .A2(_12709_),
    .B1(_02448_),
    .B2(_12713_),
    .X(_03646_));
 sky130_fd_sc_hd__clkbuf_2 _16052_ (.A(net342),
    .X(_12715_));
 sky130_fd_sc_hd__buf_2 _16053_ (.A(_12715_),
    .X(_12716_));
 sky130_fd_sc_hd__a22o_1 _16054_ (.A1(_12716_),
    .A2(_12709_),
    .B1(_02447_),
    .B2(_12713_),
    .X(_03645_));
 sky130_fd_sc_hd__buf_2 _16055_ (.A(net341),
    .X(_12717_));
 sky130_fd_sc_hd__buf_1 _16056_ (.A(_12708_),
    .X(_12718_));
 sky130_fd_sc_hd__a22o_1 _16057_ (.A1(_12717_),
    .A2(_12718_),
    .B1(_02446_),
    .B2(_12713_),
    .X(_03644_));
 sky130_fd_sc_hd__clkbuf_2 _16058_ (.A(net340),
    .X(_12719_));
 sky130_fd_sc_hd__buf_2 _16059_ (.A(_12719_),
    .X(_12720_));
 sky130_fd_sc_hd__buf_1 _16060_ (.A(_12712_),
    .X(_12721_));
 sky130_fd_sc_hd__a22o_1 _16061_ (.A1(_12720_),
    .A2(_12718_),
    .B1(_02445_),
    .B2(_12721_),
    .X(_03643_));
 sky130_fd_sc_hd__buf_2 _16062_ (.A(net339),
    .X(_12722_));
 sky130_fd_sc_hd__a22o_1 _16063_ (.A1(_12722_),
    .A2(_12718_),
    .B1(_02444_),
    .B2(_12721_),
    .X(_03642_));
 sky130_fd_sc_hd__clkbuf_2 _16064_ (.A(net369),
    .X(_12723_));
 sky130_fd_sc_hd__clkbuf_2 _16065_ (.A(_12723_),
    .X(_12724_));
 sky130_fd_sc_hd__a22o_1 _16066_ (.A1(_12724_),
    .A2(_12718_),
    .B1(_02474_),
    .B2(_12721_),
    .X(_03641_));
 sky130_fd_sc_hd__buf_2 _16067_ (.A(net368),
    .X(_12725_));
 sky130_fd_sc_hd__buf_1 _16068_ (.A(_12708_),
    .X(_12726_));
 sky130_fd_sc_hd__a22o_1 _16069_ (.A1(_12725_),
    .A2(_12726_),
    .B1(_02473_),
    .B2(_12721_),
    .X(_03640_));
 sky130_fd_sc_hd__buf_2 _16070_ (.A(net229),
    .X(_12727_));
 sky130_fd_sc_hd__clkbuf_2 _16071_ (.A(_12727_),
    .X(_12728_));
 sky130_fd_sc_hd__buf_1 _16072_ (.A(_12712_),
    .X(_12729_));
 sky130_fd_sc_hd__a22o_1 _16073_ (.A1(_12728_),
    .A2(_12726_),
    .B1(_02472_),
    .B2(_12729_),
    .X(_03639_));
 sky130_fd_sc_hd__clkbuf_2 _16074_ (.A(net228),
    .X(_12730_));
 sky130_fd_sc_hd__clkbuf_2 _16075_ (.A(_12730_),
    .X(_12731_));
 sky130_fd_sc_hd__a22o_1 _16076_ (.A1(_12731_),
    .A2(_12726_),
    .B1(_02471_),
    .B2(_12729_),
    .X(_03638_));
 sky130_fd_sc_hd__buf_2 _16077_ (.A(net227),
    .X(_12732_));
 sky130_fd_sc_hd__clkbuf_2 _16078_ (.A(_12732_),
    .X(_12733_));
 sky130_fd_sc_hd__a22o_1 _16079_ (.A1(_12733_),
    .A2(_12726_),
    .B1(_02470_),
    .B2(_12729_),
    .X(_03637_));
 sky130_fd_sc_hd__clkbuf_2 _16080_ (.A(net226),
    .X(_12734_));
 sky130_fd_sc_hd__buf_2 _16081_ (.A(_12734_),
    .X(_12735_));
 sky130_fd_sc_hd__buf_1 _16082_ (.A(_12708_),
    .X(_12736_));
 sky130_fd_sc_hd__a22o_1 _16083_ (.A1(_12735_),
    .A2(_12736_),
    .B1(_02469_),
    .B2(_12729_),
    .X(_03636_));
 sky130_fd_sc_hd__clkbuf_2 _16084_ (.A(net225),
    .X(_12737_));
 sky130_fd_sc_hd__clkbuf_2 _16085_ (.A(_12737_),
    .X(_12738_));
 sky130_fd_sc_hd__buf_1 _16086_ (.A(_12712_),
    .X(_12739_));
 sky130_fd_sc_hd__a22o_1 _16087_ (.A1(_12738_),
    .A2(_12736_),
    .B1(_02468_),
    .B2(_12739_),
    .X(_03635_));
 sky130_fd_sc_hd__clkbuf_2 _16088_ (.A(net222),
    .X(_12740_));
 sky130_fd_sc_hd__clkbuf_2 _16089_ (.A(_12740_),
    .X(_12741_));
 sky130_fd_sc_hd__a22o_1 _16090_ (.A1(_12741_),
    .A2(_12736_),
    .B1(_02465_),
    .B2(_12739_),
    .X(_03634_));
 sky130_fd_sc_hd__clkbuf_2 _16091_ (.A(net211),
    .X(_12742_));
 sky130_fd_sc_hd__buf_2 _16092_ (.A(_12742_),
    .X(_12743_));
 sky130_fd_sc_hd__a22o_1 _16093_ (.A1(_12743_),
    .A2(_12736_),
    .B1(_02454_),
    .B2(_12739_),
    .X(_03633_));
 sky130_fd_sc_hd__clkbuf_2 _16094_ (.A(net200),
    .X(_12744_));
 sky130_fd_sc_hd__clkbuf_2 _16095_ (.A(_12744_),
    .X(_12745_));
 sky130_fd_sc_hd__a22o_1 _16096_ (.A1(_12745_),
    .A2(_12689_),
    .B1(_02443_),
    .B2(_12739_),
    .X(_03632_));
 sky130_fd_sc_hd__or3_4 _16097_ (.A(_12557_),
    .B(_12564_),
    .C(_12563_),
    .X(_12746_));
 sky130_fd_sc_hd__or2_2 _16098_ (.A(_12556_),
    .B(_12746_),
    .X(_12747_));
 sky130_fd_sc_hd__clkbuf_4 _16099_ (.A(_12747_),
    .X(_12748_));
 sky130_fd_sc_hd__buf_1 _16100_ (.A(_12748_),
    .X(_12749_));
 sky130_vsdinv _16101_ (.A(_12747_),
    .Y(_12750_));
 sky130_fd_sc_hd__clkbuf_4 _16102_ (.A(_12750_),
    .X(_12751_));
 sky130_fd_sc_hd__buf_1 _16103_ (.A(_12751_),
    .X(_12752_));
 sky130_fd_sc_hd__a22o_1 _16104_ (.A1(\cpuregs[4][31] ),
    .A2(_12749_),
    .B1(_12572_),
    .B2(_12752_),
    .X(_03631_));
 sky130_fd_sc_hd__a22o_1 _16105_ (.A1(\cpuregs[4][30] ),
    .A2(_12749_),
    .B1(_12577_),
    .B2(_12752_),
    .X(_03630_));
 sky130_fd_sc_hd__a22o_1 _16106_ (.A1(\cpuregs[4][29] ),
    .A2(_12749_),
    .B1(_12579_),
    .B2(_12752_),
    .X(_03629_));
 sky130_fd_sc_hd__a22o_1 _16107_ (.A1(\cpuregs[4][28] ),
    .A2(_12749_),
    .B1(_12581_),
    .B2(_12752_),
    .X(_03628_));
 sky130_fd_sc_hd__buf_1 _16108_ (.A(_12748_),
    .X(_12753_));
 sky130_fd_sc_hd__buf_1 _16109_ (.A(_12751_),
    .X(_12754_));
 sky130_fd_sc_hd__a22o_1 _16110_ (.A1(\cpuregs[4][27] ),
    .A2(_12753_),
    .B1(_12584_),
    .B2(_12754_),
    .X(_03627_));
 sky130_fd_sc_hd__a22o_1 _16111_ (.A1(\cpuregs[4][26] ),
    .A2(_12753_),
    .B1(_12587_),
    .B2(_12754_),
    .X(_03626_));
 sky130_fd_sc_hd__a22o_1 _16112_ (.A1(\cpuregs[4][25] ),
    .A2(_12753_),
    .B1(_12589_),
    .B2(_12754_),
    .X(_03625_));
 sky130_fd_sc_hd__a22o_1 _16113_ (.A1(\cpuregs[4][24] ),
    .A2(_12753_),
    .B1(_12591_),
    .B2(_12754_),
    .X(_03624_));
 sky130_fd_sc_hd__buf_1 _16114_ (.A(_12748_),
    .X(_12755_));
 sky130_fd_sc_hd__buf_1 _16115_ (.A(_12751_),
    .X(_12756_));
 sky130_fd_sc_hd__a22o_1 _16116_ (.A1(\cpuregs[4][23] ),
    .A2(_12755_),
    .B1(_12594_),
    .B2(_12756_),
    .X(_03623_));
 sky130_fd_sc_hd__a22o_1 _16117_ (.A1(\cpuregs[4][22] ),
    .A2(_12755_),
    .B1(_12597_),
    .B2(_12756_),
    .X(_03622_));
 sky130_fd_sc_hd__a22o_1 _16118_ (.A1(\cpuregs[4][21] ),
    .A2(_12755_),
    .B1(_12599_),
    .B2(_12756_),
    .X(_03621_));
 sky130_fd_sc_hd__a22o_1 _16119_ (.A1(\cpuregs[4][20] ),
    .A2(_12755_),
    .B1(_12601_),
    .B2(_12756_),
    .X(_03620_));
 sky130_fd_sc_hd__buf_1 _16120_ (.A(_12748_),
    .X(_12757_));
 sky130_fd_sc_hd__buf_1 _16121_ (.A(_12751_),
    .X(_12758_));
 sky130_fd_sc_hd__a22o_1 _16122_ (.A1(\cpuregs[4][19] ),
    .A2(_12757_),
    .B1(_12604_),
    .B2(_12758_),
    .X(_03619_));
 sky130_fd_sc_hd__a22o_1 _16123_ (.A1(\cpuregs[4][18] ),
    .A2(_12757_),
    .B1(_12607_),
    .B2(_12758_),
    .X(_03618_));
 sky130_fd_sc_hd__a22o_1 _16124_ (.A1(\cpuregs[4][17] ),
    .A2(_12757_),
    .B1(_12609_),
    .B2(_12758_),
    .X(_03617_));
 sky130_fd_sc_hd__a22o_1 _16125_ (.A1(\cpuregs[4][16] ),
    .A2(_12757_),
    .B1(_12611_),
    .B2(_12758_),
    .X(_03616_));
 sky130_fd_sc_hd__clkbuf_2 _16126_ (.A(_12747_),
    .X(_12759_));
 sky130_fd_sc_hd__buf_1 _16127_ (.A(_12759_),
    .X(_12760_));
 sky130_fd_sc_hd__buf_2 _16128_ (.A(_12750_),
    .X(_12761_));
 sky130_fd_sc_hd__buf_1 _16129_ (.A(_12761_),
    .X(_12762_));
 sky130_fd_sc_hd__a22o_1 _16130_ (.A1(\cpuregs[4][15] ),
    .A2(_12760_),
    .B1(_12615_),
    .B2(_12762_),
    .X(_03615_));
 sky130_fd_sc_hd__a22o_1 _16131_ (.A1(\cpuregs[4][14] ),
    .A2(_12760_),
    .B1(_12619_),
    .B2(_12762_),
    .X(_03614_));
 sky130_fd_sc_hd__a22o_1 _16132_ (.A1(\cpuregs[4][13] ),
    .A2(_12760_),
    .B1(_12621_),
    .B2(_12762_),
    .X(_03613_));
 sky130_fd_sc_hd__a22o_1 _16133_ (.A1(\cpuregs[4][12] ),
    .A2(_12760_),
    .B1(_12623_),
    .B2(_12762_),
    .X(_03612_));
 sky130_fd_sc_hd__buf_1 _16134_ (.A(_12759_),
    .X(_12763_));
 sky130_fd_sc_hd__buf_1 _16135_ (.A(_12761_),
    .X(_12764_));
 sky130_fd_sc_hd__a22o_1 _16136_ (.A1(\cpuregs[4][11] ),
    .A2(_12763_),
    .B1(_12626_),
    .B2(_12764_),
    .X(_03611_));
 sky130_fd_sc_hd__a22o_1 _16137_ (.A1(\cpuregs[4][10] ),
    .A2(_12763_),
    .B1(_12629_),
    .B2(_12764_),
    .X(_03610_));
 sky130_fd_sc_hd__a22o_1 _16138_ (.A1(\cpuregs[4][9] ),
    .A2(_12763_),
    .B1(_12631_),
    .B2(_12764_),
    .X(_03609_));
 sky130_fd_sc_hd__a22o_1 _16139_ (.A1(\cpuregs[4][8] ),
    .A2(_12763_),
    .B1(_12633_),
    .B2(_12764_),
    .X(_03608_));
 sky130_fd_sc_hd__buf_1 _16140_ (.A(_12759_),
    .X(_12765_));
 sky130_fd_sc_hd__buf_1 _16141_ (.A(_12761_),
    .X(_12766_));
 sky130_fd_sc_hd__a22o_1 _16142_ (.A1(\cpuregs[4][7] ),
    .A2(_12765_),
    .B1(_12636_),
    .B2(_12766_),
    .X(_03607_));
 sky130_fd_sc_hd__a22o_1 _16143_ (.A1(\cpuregs[4][6] ),
    .A2(_12765_),
    .B1(_12639_),
    .B2(_12766_),
    .X(_03606_));
 sky130_fd_sc_hd__a22o_1 _16144_ (.A1(\cpuregs[4][5] ),
    .A2(_12765_),
    .B1(_12641_),
    .B2(_12766_),
    .X(_03605_));
 sky130_fd_sc_hd__a22o_1 _16145_ (.A1(\cpuregs[4][4] ),
    .A2(_12765_),
    .B1(_12643_),
    .B2(_12766_),
    .X(_03604_));
 sky130_fd_sc_hd__buf_1 _16146_ (.A(_12759_),
    .X(_12767_));
 sky130_fd_sc_hd__buf_1 _16147_ (.A(_12761_),
    .X(_12768_));
 sky130_fd_sc_hd__a22o_1 _16148_ (.A1(\cpuregs[4][3] ),
    .A2(_12767_),
    .B1(_12646_),
    .B2(_12768_),
    .X(_03603_));
 sky130_fd_sc_hd__a22o_1 _16149_ (.A1(\cpuregs[4][2] ),
    .A2(_12767_),
    .B1(_12649_),
    .B2(_12768_),
    .X(_03602_));
 sky130_fd_sc_hd__a22o_1 _16150_ (.A1(\cpuregs[4][1] ),
    .A2(_12767_),
    .B1(_12651_),
    .B2(_12768_),
    .X(_03601_));
 sky130_fd_sc_hd__a22o_1 _16151_ (.A1(\cpuregs[4][0] ),
    .A2(_12767_),
    .B1(_12653_),
    .B2(_12768_),
    .X(_03600_));
 sky130_vsdinv _16152_ (.A(_12552_),
    .Y(_12769_));
 sky130_fd_sc_hd__buf_2 _16153_ (.A(_12554_),
    .X(_12770_));
 sky130_fd_sc_hd__buf_2 _16154_ (.A(_12553_),
    .X(_12771_));
 sky130_fd_sc_hd__or2_1 _16155_ (.A(_12656_),
    .B(_12565_),
    .X(_12772_));
 sky130_fd_sc_hd__or4_4 _16156_ (.A(_12769_),
    .B(_12770_),
    .C(_12771_),
    .D(_12772_),
    .X(_12773_));
 sky130_fd_sc_hd__clkbuf_4 _16157_ (.A(_12773_),
    .X(_12774_));
 sky130_fd_sc_hd__buf_1 _16158_ (.A(_12774_),
    .X(_12775_));
 sky130_vsdinv _16159_ (.A(_12773_),
    .Y(_12776_));
 sky130_fd_sc_hd__clkbuf_4 _16160_ (.A(_12776_),
    .X(_12777_));
 sky130_fd_sc_hd__buf_1 _16161_ (.A(_12777_),
    .X(_12778_));
 sky130_fd_sc_hd__a22o_1 _16162_ (.A1(\cpuregs[19][31] ),
    .A2(_12775_),
    .B1(_12572_),
    .B2(_12778_),
    .X(_03599_));
 sky130_fd_sc_hd__a22o_1 _16163_ (.A1(\cpuregs[19][30] ),
    .A2(_12775_),
    .B1(_12577_),
    .B2(_12778_),
    .X(_03598_));
 sky130_fd_sc_hd__a22o_1 _16164_ (.A1(\cpuregs[19][29] ),
    .A2(_12775_),
    .B1(_12579_),
    .B2(_12778_),
    .X(_03597_));
 sky130_fd_sc_hd__a22o_1 _16165_ (.A1(\cpuregs[19][28] ),
    .A2(_12775_),
    .B1(_12581_),
    .B2(_12778_),
    .X(_03596_));
 sky130_fd_sc_hd__buf_1 _16166_ (.A(_12774_),
    .X(_12779_));
 sky130_fd_sc_hd__buf_1 _16167_ (.A(_12777_),
    .X(_12780_));
 sky130_fd_sc_hd__a22o_1 _16168_ (.A1(\cpuregs[19][27] ),
    .A2(_12779_),
    .B1(_12584_),
    .B2(_12780_),
    .X(_03595_));
 sky130_fd_sc_hd__a22o_1 _16169_ (.A1(\cpuregs[19][26] ),
    .A2(_12779_),
    .B1(_12587_),
    .B2(_12780_),
    .X(_03594_));
 sky130_fd_sc_hd__a22o_1 _16170_ (.A1(\cpuregs[19][25] ),
    .A2(_12779_),
    .B1(_12589_),
    .B2(_12780_),
    .X(_03593_));
 sky130_fd_sc_hd__a22o_1 _16171_ (.A1(\cpuregs[19][24] ),
    .A2(_12779_),
    .B1(_12591_),
    .B2(_12780_),
    .X(_03592_));
 sky130_fd_sc_hd__buf_1 _16172_ (.A(_12774_),
    .X(_12781_));
 sky130_fd_sc_hd__buf_1 _16173_ (.A(_12777_),
    .X(_12782_));
 sky130_fd_sc_hd__a22o_1 _16174_ (.A1(\cpuregs[19][23] ),
    .A2(_12781_),
    .B1(_12594_),
    .B2(_12782_),
    .X(_03591_));
 sky130_fd_sc_hd__a22o_1 _16175_ (.A1(\cpuregs[19][22] ),
    .A2(_12781_),
    .B1(_12597_),
    .B2(_12782_),
    .X(_03590_));
 sky130_fd_sc_hd__a22o_1 _16176_ (.A1(\cpuregs[19][21] ),
    .A2(_12781_),
    .B1(_12599_),
    .B2(_12782_),
    .X(_03589_));
 sky130_fd_sc_hd__a22o_1 _16177_ (.A1(\cpuregs[19][20] ),
    .A2(_12781_),
    .B1(_12601_),
    .B2(_12782_),
    .X(_03588_));
 sky130_fd_sc_hd__buf_1 _16178_ (.A(_12774_),
    .X(_12783_));
 sky130_fd_sc_hd__buf_1 _16179_ (.A(_12777_),
    .X(_12784_));
 sky130_fd_sc_hd__a22o_1 _16180_ (.A1(\cpuregs[19][19] ),
    .A2(_12783_),
    .B1(_12604_),
    .B2(_12784_),
    .X(_03587_));
 sky130_fd_sc_hd__a22o_1 _16181_ (.A1(\cpuregs[19][18] ),
    .A2(_12783_),
    .B1(_12607_),
    .B2(_12784_),
    .X(_03586_));
 sky130_fd_sc_hd__a22o_1 _16182_ (.A1(\cpuregs[19][17] ),
    .A2(_12783_),
    .B1(_12609_),
    .B2(_12784_),
    .X(_03585_));
 sky130_fd_sc_hd__a22o_1 _16183_ (.A1(\cpuregs[19][16] ),
    .A2(_12783_),
    .B1(_12611_),
    .B2(_12784_),
    .X(_03584_));
 sky130_fd_sc_hd__buf_2 _16184_ (.A(_12773_),
    .X(_12785_));
 sky130_fd_sc_hd__buf_1 _16185_ (.A(_12785_),
    .X(_12786_));
 sky130_fd_sc_hd__buf_2 _16186_ (.A(_12776_),
    .X(_12787_));
 sky130_fd_sc_hd__buf_1 _16187_ (.A(_12787_),
    .X(_12788_));
 sky130_fd_sc_hd__a22o_1 _16188_ (.A1(\cpuregs[19][15] ),
    .A2(_12786_),
    .B1(_12615_),
    .B2(_12788_),
    .X(_03583_));
 sky130_fd_sc_hd__a22o_1 _16189_ (.A1(\cpuregs[19][14] ),
    .A2(_12786_),
    .B1(_12619_),
    .B2(_12788_),
    .X(_03582_));
 sky130_fd_sc_hd__a22o_1 _16190_ (.A1(\cpuregs[19][13] ),
    .A2(_12786_),
    .B1(_12621_),
    .B2(_12788_),
    .X(_03581_));
 sky130_fd_sc_hd__a22o_1 _16191_ (.A1(\cpuregs[19][12] ),
    .A2(_12786_),
    .B1(_12623_),
    .B2(_12788_),
    .X(_03580_));
 sky130_fd_sc_hd__buf_1 _16192_ (.A(_12785_),
    .X(_12789_));
 sky130_fd_sc_hd__buf_1 _16193_ (.A(_12787_),
    .X(_12790_));
 sky130_fd_sc_hd__a22o_1 _16194_ (.A1(\cpuregs[19][11] ),
    .A2(_12789_),
    .B1(_12626_),
    .B2(_12790_),
    .X(_03579_));
 sky130_fd_sc_hd__a22o_1 _16195_ (.A1(\cpuregs[19][10] ),
    .A2(_12789_),
    .B1(_12629_),
    .B2(_12790_),
    .X(_03578_));
 sky130_fd_sc_hd__a22o_1 _16196_ (.A1(\cpuregs[19][9] ),
    .A2(_12789_),
    .B1(_12631_),
    .B2(_12790_),
    .X(_03577_));
 sky130_fd_sc_hd__a22o_1 _16197_ (.A1(\cpuregs[19][8] ),
    .A2(_12789_),
    .B1(_12633_),
    .B2(_12790_),
    .X(_03576_));
 sky130_fd_sc_hd__buf_1 _16198_ (.A(_12785_),
    .X(_12791_));
 sky130_fd_sc_hd__buf_1 _16199_ (.A(_12787_),
    .X(_12792_));
 sky130_fd_sc_hd__a22o_1 _16200_ (.A1(\cpuregs[19][7] ),
    .A2(_12791_),
    .B1(_12636_),
    .B2(_12792_),
    .X(_03575_));
 sky130_fd_sc_hd__a22o_1 _16201_ (.A1(\cpuregs[19][6] ),
    .A2(_12791_),
    .B1(_12639_),
    .B2(_12792_),
    .X(_03574_));
 sky130_fd_sc_hd__a22o_1 _16202_ (.A1(\cpuregs[19][5] ),
    .A2(_12791_),
    .B1(_12641_),
    .B2(_12792_),
    .X(_03573_));
 sky130_fd_sc_hd__a22o_1 _16203_ (.A1(\cpuregs[19][4] ),
    .A2(_12791_),
    .B1(_12643_),
    .B2(_12792_),
    .X(_03572_));
 sky130_fd_sc_hd__buf_1 _16204_ (.A(_12785_),
    .X(_12793_));
 sky130_fd_sc_hd__buf_1 _16205_ (.A(_12787_),
    .X(_12794_));
 sky130_fd_sc_hd__a22o_1 _16206_ (.A1(\cpuregs[19][3] ),
    .A2(_12793_),
    .B1(_12646_),
    .B2(_12794_),
    .X(_03571_));
 sky130_fd_sc_hd__a22o_1 _16207_ (.A1(\cpuregs[19][2] ),
    .A2(_12793_),
    .B1(_12649_),
    .B2(_12794_),
    .X(_03570_));
 sky130_fd_sc_hd__a22o_1 _16208_ (.A1(\cpuregs[19][1] ),
    .A2(_12793_),
    .B1(_12651_),
    .B2(_12794_),
    .X(_03569_));
 sky130_fd_sc_hd__a22o_1 _16209_ (.A1(\cpuregs[19][0] ),
    .A2(_12793_),
    .B1(_12653_),
    .B2(_12794_),
    .X(_03568_));
 sky130_fd_sc_hd__or3_1 _16210_ (.A(_11579_),
    .B(_11591_),
    .C(_11878_),
    .X(_12795_));
 sky130_fd_sc_hd__or2_4 _16211_ (.A(_11582_),
    .B(_12795_),
    .X(_12796_));
 sky130_fd_sc_hd__buf_1 _16212_ (.A(_12796_),
    .X(_12797_));
 sky130_fd_sc_hd__buf_1 _16213_ (.A(_12797_),
    .X(_12798_));
 sky130_vsdinv _16214_ (.A(_12796_),
    .Y(_12799_));
 sky130_fd_sc_hd__buf_1 _16215_ (.A(_12799_),
    .X(_12800_));
 sky130_fd_sc_hd__buf_1 _16216_ (.A(_12800_),
    .X(_12801_));
 sky130_fd_sc_hd__a22o_1 _16217_ (.A1(net262),
    .A2(_12798_),
    .B1(net224),
    .B2(_12801_),
    .X(_03567_));
 sky130_fd_sc_hd__a22o_1 _16218_ (.A1(net261),
    .A2(_12798_),
    .B1(net223),
    .B2(_12801_),
    .X(_03566_));
 sky130_fd_sc_hd__a22o_1 _16219_ (.A1(net259),
    .A2(_12798_),
    .B1(net221),
    .B2(_12801_),
    .X(_03565_));
 sky130_fd_sc_hd__a22o_1 _16220_ (.A1(net258),
    .A2(_12798_),
    .B1(net220),
    .B2(_12801_),
    .X(_03564_));
 sky130_fd_sc_hd__buf_1 _16221_ (.A(_12797_),
    .X(_12802_));
 sky130_fd_sc_hd__buf_1 _16222_ (.A(_12800_),
    .X(_12803_));
 sky130_fd_sc_hd__a22o_1 _16223_ (.A1(net257),
    .A2(_12802_),
    .B1(net219),
    .B2(_12803_),
    .X(_03563_));
 sky130_fd_sc_hd__a22o_1 _16224_ (.A1(net256),
    .A2(_12802_),
    .B1(net218),
    .B2(_12803_),
    .X(_03562_));
 sky130_fd_sc_hd__a22o_1 _16225_ (.A1(net255),
    .A2(_12802_),
    .B1(net217),
    .B2(_12803_),
    .X(_03561_));
 sky130_fd_sc_hd__a22o_1 _16226_ (.A1(net254),
    .A2(_12802_),
    .B1(net216),
    .B2(_12803_),
    .X(_03560_));
 sky130_fd_sc_hd__buf_1 _16227_ (.A(_12797_),
    .X(_12804_));
 sky130_fd_sc_hd__buf_1 _16228_ (.A(_12800_),
    .X(_12805_));
 sky130_fd_sc_hd__a22o_1 _16229_ (.A1(net253),
    .A2(_12804_),
    .B1(net215),
    .B2(_12805_),
    .X(_03559_));
 sky130_fd_sc_hd__a22o_1 _16230_ (.A1(net252),
    .A2(_12804_),
    .B1(net214),
    .B2(_12805_),
    .X(_03558_));
 sky130_fd_sc_hd__a22o_1 _16231_ (.A1(net251),
    .A2(_12804_),
    .B1(net213),
    .B2(_12805_),
    .X(_03557_));
 sky130_fd_sc_hd__a22o_1 _16232_ (.A1(net250),
    .A2(_12804_),
    .B1(net212),
    .B2(_12805_),
    .X(_03556_));
 sky130_fd_sc_hd__clkbuf_2 _16233_ (.A(_12797_),
    .X(_12806_));
 sky130_fd_sc_hd__clkbuf_2 _16234_ (.A(_12800_),
    .X(_12807_));
 sky130_fd_sc_hd__a22o_1 _16235_ (.A1(net248),
    .A2(_12806_),
    .B1(net210),
    .B2(_12807_),
    .X(_03555_));
 sky130_fd_sc_hd__a22o_1 _16236_ (.A1(net247),
    .A2(_12806_),
    .B1(net209),
    .B2(_12807_),
    .X(_03554_));
 sky130_fd_sc_hd__a22o_1 _16237_ (.A1(net246),
    .A2(_12806_),
    .B1(net208),
    .B2(_12807_),
    .X(_03553_));
 sky130_fd_sc_hd__a22o_1 _16238_ (.A1(net245),
    .A2(_12806_),
    .B1(net207),
    .B2(_12807_),
    .X(_03552_));
 sky130_fd_sc_hd__buf_1 _16239_ (.A(_12796_),
    .X(_12808_));
 sky130_fd_sc_hd__buf_1 _16240_ (.A(_12808_),
    .X(_12809_));
 sky130_fd_sc_hd__buf_1 _16241_ (.A(_12799_),
    .X(_12810_));
 sky130_fd_sc_hd__buf_1 _16242_ (.A(_12810_),
    .X(_12811_));
 sky130_fd_sc_hd__a22o_1 _16243_ (.A1(net244),
    .A2(_12809_),
    .B1(net206),
    .B2(_12811_),
    .X(_03551_));
 sky130_fd_sc_hd__a22o_1 _16244_ (.A1(net243),
    .A2(_12809_),
    .B1(net205),
    .B2(_12811_),
    .X(_03550_));
 sky130_fd_sc_hd__a22o_1 _16245_ (.A1(net242),
    .A2(_12809_),
    .B1(net204),
    .B2(_12811_),
    .X(_03549_));
 sky130_fd_sc_hd__a22o_1 _16246_ (.A1(net241),
    .A2(_12809_),
    .B1(net203),
    .B2(_12811_),
    .X(_03548_));
 sky130_fd_sc_hd__clkbuf_2 _16247_ (.A(_12808_),
    .X(_12812_));
 sky130_fd_sc_hd__clkbuf_2 _16248_ (.A(_12810_),
    .X(_12813_));
 sky130_fd_sc_hd__a22o_1 _16249_ (.A1(net240),
    .A2(_12812_),
    .B1(net202),
    .B2(_12813_),
    .X(_03547_));
 sky130_fd_sc_hd__a22o_1 _16250_ (.A1(net239),
    .A2(_12812_),
    .B1(net201),
    .B2(_12813_),
    .X(_03546_));
 sky130_fd_sc_hd__a22o_1 _16251_ (.A1(net269),
    .A2(_12812_),
    .B1(net231),
    .B2(_12813_),
    .X(_03545_));
 sky130_fd_sc_hd__a22o_1 _16252_ (.A1(net268),
    .A2(_12812_),
    .B1(net230),
    .B2(_12813_),
    .X(_03544_));
 sky130_fd_sc_hd__clkbuf_2 _16253_ (.A(_12808_),
    .X(_12814_));
 sky130_fd_sc_hd__clkbuf_2 _16254_ (.A(_12810_),
    .X(_12815_));
 sky130_fd_sc_hd__a22o_1 _16255_ (.A1(net267),
    .A2(_12814_),
    .B1(_12728_),
    .B2(_12815_),
    .X(_03543_));
 sky130_fd_sc_hd__a22o_1 _16256_ (.A1(net266),
    .A2(_12814_),
    .B1(_12731_),
    .B2(_12815_),
    .X(_03542_));
 sky130_fd_sc_hd__a22o_1 _16257_ (.A1(net265),
    .A2(_12814_),
    .B1(_12733_),
    .B2(_12815_),
    .X(_03541_));
 sky130_fd_sc_hd__a22o_1 _16258_ (.A1(net264),
    .A2(_12814_),
    .B1(_12735_),
    .B2(_12815_),
    .X(_03540_));
 sky130_fd_sc_hd__buf_1 _16259_ (.A(_12808_),
    .X(_12816_));
 sky130_fd_sc_hd__buf_1 _16260_ (.A(_12810_),
    .X(_12817_));
 sky130_fd_sc_hd__a22o_1 _16261_ (.A1(net263),
    .A2(_12816_),
    .B1(_12738_),
    .B2(_12817_),
    .X(_03539_));
 sky130_fd_sc_hd__a22o_1 _16262_ (.A1(net260),
    .A2(_12816_),
    .B1(_12741_),
    .B2(_12817_),
    .X(_03538_));
 sky130_fd_sc_hd__a22o_1 _16263_ (.A1(net249),
    .A2(_12816_),
    .B1(_12743_),
    .B2(_12817_),
    .X(_03537_));
 sky130_fd_sc_hd__a22o_1 _16264_ (.A1(net238),
    .A2(_12816_),
    .B1(_12745_),
    .B2(_12817_),
    .X(_03536_));
 sky130_fd_sc_hd__buf_1 _16265_ (.A(_12772_),
    .X(_12818_));
 sky130_fd_sc_hd__or2_2 _16266_ (.A(_12556_),
    .B(_12818_),
    .X(_12819_));
 sky130_fd_sc_hd__clkbuf_4 _16267_ (.A(_12819_),
    .X(_12820_));
 sky130_fd_sc_hd__buf_1 _16268_ (.A(_12820_),
    .X(_12821_));
 sky130_fd_sc_hd__buf_2 _16269_ (.A(\cpuregs_wrdata[31] ),
    .X(_12822_));
 sky130_vsdinv _16270_ (.A(_12819_),
    .Y(_12823_));
 sky130_fd_sc_hd__clkbuf_4 _16271_ (.A(_12823_),
    .X(_12824_));
 sky130_fd_sc_hd__buf_1 _16272_ (.A(_12824_),
    .X(_12825_));
 sky130_fd_sc_hd__a22o_1 _16273_ (.A1(\cpuregs[7][31] ),
    .A2(_12821_),
    .B1(_12822_),
    .B2(_12825_),
    .X(_03535_));
 sky130_fd_sc_hd__buf_2 _16274_ (.A(\cpuregs_wrdata[30] ),
    .X(_12826_));
 sky130_fd_sc_hd__a22o_1 _16275_ (.A1(\cpuregs[7][30] ),
    .A2(_12821_),
    .B1(_12826_),
    .B2(_12825_),
    .X(_03534_));
 sky130_fd_sc_hd__buf_2 _16276_ (.A(\cpuregs_wrdata[29] ),
    .X(_12827_));
 sky130_fd_sc_hd__a22o_1 _16277_ (.A1(\cpuregs[7][29] ),
    .A2(_12821_),
    .B1(_12827_),
    .B2(_12825_),
    .X(_03533_));
 sky130_fd_sc_hd__buf_2 _16278_ (.A(\cpuregs_wrdata[28] ),
    .X(_12828_));
 sky130_fd_sc_hd__a22o_1 _16279_ (.A1(\cpuregs[7][28] ),
    .A2(_12821_),
    .B1(_12828_),
    .B2(_12825_),
    .X(_03532_));
 sky130_fd_sc_hd__buf_1 _16280_ (.A(_12820_),
    .X(_12829_));
 sky130_fd_sc_hd__clkbuf_2 _16281_ (.A(\cpuregs_wrdata[27] ),
    .X(_12830_));
 sky130_fd_sc_hd__buf_1 _16282_ (.A(_12824_),
    .X(_12831_));
 sky130_fd_sc_hd__a22o_1 _16283_ (.A1(\cpuregs[7][27] ),
    .A2(_12829_),
    .B1(_12830_),
    .B2(_12831_),
    .X(_03531_));
 sky130_fd_sc_hd__clkbuf_2 _16284_ (.A(\cpuregs_wrdata[26] ),
    .X(_12832_));
 sky130_fd_sc_hd__a22o_1 _16285_ (.A1(\cpuregs[7][26] ),
    .A2(_12829_),
    .B1(_12832_),
    .B2(_12831_),
    .X(_03530_));
 sky130_fd_sc_hd__clkbuf_2 _16286_ (.A(\cpuregs_wrdata[25] ),
    .X(_12833_));
 sky130_fd_sc_hd__a22o_1 _16287_ (.A1(\cpuregs[7][25] ),
    .A2(_12829_),
    .B1(_12833_),
    .B2(_12831_),
    .X(_03529_));
 sky130_fd_sc_hd__clkbuf_2 _16288_ (.A(\cpuregs_wrdata[24] ),
    .X(_12834_));
 sky130_fd_sc_hd__a22o_1 _16289_ (.A1(\cpuregs[7][24] ),
    .A2(_12829_),
    .B1(_12834_),
    .B2(_12831_),
    .X(_03528_));
 sky130_fd_sc_hd__buf_1 _16290_ (.A(_12820_),
    .X(_12835_));
 sky130_fd_sc_hd__clkbuf_2 _16291_ (.A(\cpuregs_wrdata[23] ),
    .X(_12836_));
 sky130_fd_sc_hd__buf_1 _16292_ (.A(_12824_),
    .X(_12837_));
 sky130_fd_sc_hd__a22o_1 _16293_ (.A1(\cpuregs[7][23] ),
    .A2(_12835_),
    .B1(_12836_),
    .B2(_12837_),
    .X(_03527_));
 sky130_fd_sc_hd__clkbuf_2 _16294_ (.A(\cpuregs_wrdata[22] ),
    .X(_12838_));
 sky130_fd_sc_hd__a22o_1 _16295_ (.A1(\cpuregs[7][22] ),
    .A2(_12835_),
    .B1(_12838_),
    .B2(_12837_),
    .X(_03526_));
 sky130_fd_sc_hd__clkbuf_2 _16296_ (.A(\cpuregs_wrdata[21] ),
    .X(_12839_));
 sky130_fd_sc_hd__a22o_1 _16297_ (.A1(\cpuregs[7][21] ),
    .A2(_12835_),
    .B1(_12839_),
    .B2(_12837_),
    .X(_03525_));
 sky130_fd_sc_hd__clkbuf_2 _16298_ (.A(\cpuregs_wrdata[20] ),
    .X(_12840_));
 sky130_fd_sc_hd__a22o_1 _16299_ (.A1(\cpuregs[7][20] ),
    .A2(_12835_),
    .B1(_12840_),
    .B2(_12837_),
    .X(_03524_));
 sky130_fd_sc_hd__buf_1 _16300_ (.A(_12820_),
    .X(_12841_));
 sky130_fd_sc_hd__clkbuf_2 _16301_ (.A(\cpuregs_wrdata[19] ),
    .X(_12842_));
 sky130_fd_sc_hd__buf_1 _16302_ (.A(_12824_),
    .X(_12843_));
 sky130_fd_sc_hd__a22o_1 _16303_ (.A1(\cpuregs[7][19] ),
    .A2(_12841_),
    .B1(_12842_),
    .B2(_12843_),
    .X(_03523_));
 sky130_fd_sc_hd__clkbuf_2 _16304_ (.A(\cpuregs_wrdata[18] ),
    .X(_12844_));
 sky130_fd_sc_hd__a22o_1 _16305_ (.A1(\cpuregs[7][18] ),
    .A2(_12841_),
    .B1(_12844_),
    .B2(_12843_),
    .X(_03522_));
 sky130_fd_sc_hd__clkbuf_2 _16306_ (.A(\cpuregs_wrdata[17] ),
    .X(_12845_));
 sky130_fd_sc_hd__a22o_1 _16307_ (.A1(\cpuregs[7][17] ),
    .A2(_12841_),
    .B1(_12845_),
    .B2(_12843_),
    .X(_03521_));
 sky130_fd_sc_hd__clkbuf_2 _16308_ (.A(\cpuregs_wrdata[16] ),
    .X(_12846_));
 sky130_fd_sc_hd__a22o_1 _16309_ (.A1(\cpuregs[7][16] ),
    .A2(_12841_),
    .B1(_12846_),
    .B2(_12843_),
    .X(_03520_));
 sky130_fd_sc_hd__buf_2 _16310_ (.A(_12819_),
    .X(_12847_));
 sky130_fd_sc_hd__buf_1 _16311_ (.A(_12847_),
    .X(_12848_));
 sky130_fd_sc_hd__buf_2 _16312_ (.A(\cpuregs_wrdata[15] ),
    .X(_12849_));
 sky130_fd_sc_hd__buf_2 _16313_ (.A(_12823_),
    .X(_12850_));
 sky130_fd_sc_hd__buf_1 _16314_ (.A(_12850_),
    .X(_12851_));
 sky130_fd_sc_hd__a22o_1 _16315_ (.A1(\cpuregs[7][15] ),
    .A2(_12848_),
    .B1(_12849_),
    .B2(_12851_),
    .X(_03519_));
 sky130_fd_sc_hd__buf_2 _16316_ (.A(\cpuregs_wrdata[14] ),
    .X(_12852_));
 sky130_fd_sc_hd__a22o_1 _16317_ (.A1(\cpuregs[7][14] ),
    .A2(_12848_),
    .B1(_12852_),
    .B2(_12851_),
    .X(_03518_));
 sky130_fd_sc_hd__buf_2 _16318_ (.A(\cpuregs_wrdata[13] ),
    .X(_12853_));
 sky130_fd_sc_hd__a22o_1 _16319_ (.A1(\cpuregs[7][13] ),
    .A2(_12848_),
    .B1(_12853_),
    .B2(_12851_),
    .X(_03517_));
 sky130_fd_sc_hd__buf_2 _16320_ (.A(\cpuregs_wrdata[12] ),
    .X(_12854_));
 sky130_fd_sc_hd__a22o_1 _16321_ (.A1(\cpuregs[7][12] ),
    .A2(_12848_),
    .B1(_12854_),
    .B2(_12851_),
    .X(_03516_));
 sky130_fd_sc_hd__buf_1 _16322_ (.A(_12847_),
    .X(_12855_));
 sky130_fd_sc_hd__clkbuf_2 _16323_ (.A(\cpuregs_wrdata[11] ),
    .X(_12856_));
 sky130_fd_sc_hd__buf_1 _16324_ (.A(_12850_),
    .X(_12857_));
 sky130_fd_sc_hd__a22o_1 _16325_ (.A1(\cpuregs[7][11] ),
    .A2(_12855_),
    .B1(_12856_),
    .B2(_12857_),
    .X(_03515_));
 sky130_fd_sc_hd__clkbuf_2 _16326_ (.A(\cpuregs_wrdata[10] ),
    .X(_12858_));
 sky130_fd_sc_hd__a22o_1 _16327_ (.A1(\cpuregs[7][10] ),
    .A2(_12855_),
    .B1(_12858_),
    .B2(_12857_),
    .X(_03514_));
 sky130_fd_sc_hd__clkbuf_2 _16328_ (.A(\cpuregs_wrdata[9] ),
    .X(_12859_));
 sky130_fd_sc_hd__a22o_1 _16329_ (.A1(\cpuregs[7][9] ),
    .A2(_12855_),
    .B1(_12859_),
    .B2(_12857_),
    .X(_03513_));
 sky130_fd_sc_hd__clkbuf_2 _16330_ (.A(\cpuregs_wrdata[8] ),
    .X(_12860_));
 sky130_fd_sc_hd__a22o_1 _16331_ (.A1(\cpuregs[7][8] ),
    .A2(_12855_),
    .B1(_12860_),
    .B2(_12857_),
    .X(_03512_));
 sky130_fd_sc_hd__buf_1 _16332_ (.A(_12847_),
    .X(_12861_));
 sky130_fd_sc_hd__buf_2 _16333_ (.A(\cpuregs_wrdata[7] ),
    .X(_12862_));
 sky130_fd_sc_hd__buf_1 _16334_ (.A(_12850_),
    .X(_12863_));
 sky130_fd_sc_hd__a22o_1 _16335_ (.A1(\cpuregs[7][7] ),
    .A2(_12861_),
    .B1(_12862_),
    .B2(_12863_),
    .X(_03511_));
 sky130_fd_sc_hd__clkbuf_2 _16336_ (.A(\cpuregs_wrdata[6] ),
    .X(_12864_));
 sky130_fd_sc_hd__a22o_1 _16337_ (.A1(\cpuregs[7][6] ),
    .A2(_12861_),
    .B1(_12864_),
    .B2(_12863_),
    .X(_03510_));
 sky130_fd_sc_hd__buf_2 _16338_ (.A(\cpuregs_wrdata[5] ),
    .X(_12865_));
 sky130_fd_sc_hd__a22o_1 _16339_ (.A1(\cpuregs[7][5] ),
    .A2(_12861_),
    .B1(_12865_),
    .B2(_12863_),
    .X(_03509_));
 sky130_fd_sc_hd__buf_2 _16340_ (.A(\cpuregs_wrdata[4] ),
    .X(_12866_));
 sky130_fd_sc_hd__a22o_1 _16341_ (.A1(\cpuregs[7][4] ),
    .A2(_12861_),
    .B1(_12866_),
    .B2(_12863_),
    .X(_03508_));
 sky130_fd_sc_hd__buf_1 _16342_ (.A(_12847_),
    .X(_12867_));
 sky130_fd_sc_hd__clkbuf_2 _16343_ (.A(\cpuregs_wrdata[3] ),
    .X(_12868_));
 sky130_fd_sc_hd__buf_1 _16344_ (.A(_12850_),
    .X(_12869_));
 sky130_fd_sc_hd__a22o_1 _16345_ (.A1(\cpuregs[7][3] ),
    .A2(_12867_),
    .B1(_12868_),
    .B2(_12869_),
    .X(_03507_));
 sky130_fd_sc_hd__clkbuf_2 _16346_ (.A(\cpuregs_wrdata[2] ),
    .X(_12870_));
 sky130_fd_sc_hd__a22o_1 _16347_ (.A1(\cpuregs[7][2] ),
    .A2(_12867_),
    .B1(_12870_),
    .B2(_12869_),
    .X(_03506_));
 sky130_fd_sc_hd__clkbuf_2 _16348_ (.A(\cpuregs_wrdata[1] ),
    .X(_12871_));
 sky130_fd_sc_hd__a22o_1 _16349_ (.A1(\cpuregs[7][1] ),
    .A2(_12867_),
    .B1(_12871_),
    .B2(_12869_),
    .X(_03505_));
 sky130_fd_sc_hd__clkbuf_2 _16350_ (.A(\cpuregs_wrdata[0] ),
    .X(_12872_));
 sky130_fd_sc_hd__a22o_1 _16351_ (.A1(\cpuregs[7][0] ),
    .A2(_12867_),
    .B1(_12872_),
    .B2(_12869_),
    .X(_03504_));
 sky130_vsdinv _16352_ (.A(instr_setq),
    .Y(_12873_));
 sky130_fd_sc_hd__and3_2 _16353_ (.A(\cpu_state[4] ),
    .B(_11728_),
    .C(_00302_),
    .X(_12874_));
 sky130_fd_sc_hd__a2111o_4 _16354_ (.A1(_12873_),
    .A2(_12274_),
    .B1(_11767_),
    .C1(_00331_),
    .D1(_12874_),
    .X(_12875_));
 sky130_fd_sc_hd__mux2_1 _16355_ (.A0(_14282_),
    .A1(_12552_),
    .S(_12875_),
    .X(_03503_));
 sky130_fd_sc_hd__or3_1 _16356_ (.A(_12552_),
    .B(_12654_),
    .C(_12555_),
    .X(_12876_));
 sky130_fd_sc_hd__or2_1 _16357_ (.A(_12818_),
    .B(_12876_),
    .X(_12877_));
 sky130_fd_sc_hd__clkbuf_4 _16358_ (.A(_12877_),
    .X(_12878_));
 sky130_fd_sc_hd__buf_1 _16359_ (.A(_12878_),
    .X(_12879_));
 sky130_vsdinv _16360_ (.A(_12877_),
    .Y(_12880_));
 sky130_fd_sc_hd__buf_4 _16361_ (.A(_12880_),
    .X(_12881_));
 sky130_fd_sc_hd__buf_1 _16362_ (.A(_12881_),
    .X(_12882_));
 sky130_fd_sc_hd__a22o_1 _16363_ (.A1(\cpuregs[15][31] ),
    .A2(_12879_),
    .B1(_12822_),
    .B2(_12882_),
    .X(_03502_));
 sky130_fd_sc_hd__a22o_1 _16364_ (.A1(\cpuregs[15][30] ),
    .A2(_12879_),
    .B1(_12826_),
    .B2(_12882_),
    .X(_03501_));
 sky130_fd_sc_hd__a22o_1 _16365_ (.A1(\cpuregs[15][29] ),
    .A2(_12879_),
    .B1(_12827_),
    .B2(_12882_),
    .X(_03500_));
 sky130_fd_sc_hd__a22o_1 _16366_ (.A1(\cpuregs[15][28] ),
    .A2(_12879_),
    .B1(_12828_),
    .B2(_12882_),
    .X(_03499_));
 sky130_fd_sc_hd__buf_1 _16367_ (.A(_12878_),
    .X(_12883_));
 sky130_fd_sc_hd__buf_1 _16368_ (.A(_12881_),
    .X(_12884_));
 sky130_fd_sc_hd__a22o_1 _16369_ (.A1(\cpuregs[15][27] ),
    .A2(_12883_),
    .B1(_12830_),
    .B2(_12884_),
    .X(_03498_));
 sky130_fd_sc_hd__a22o_1 _16370_ (.A1(\cpuregs[15][26] ),
    .A2(_12883_),
    .B1(_12832_),
    .B2(_12884_),
    .X(_03497_));
 sky130_fd_sc_hd__a22o_1 _16371_ (.A1(\cpuregs[15][25] ),
    .A2(_12883_),
    .B1(_12833_),
    .B2(_12884_),
    .X(_03496_));
 sky130_fd_sc_hd__a22o_1 _16372_ (.A1(\cpuregs[15][24] ),
    .A2(_12883_),
    .B1(_12834_),
    .B2(_12884_),
    .X(_03495_));
 sky130_fd_sc_hd__buf_1 _16373_ (.A(_12878_),
    .X(_12885_));
 sky130_fd_sc_hd__buf_1 _16374_ (.A(_12881_),
    .X(_12886_));
 sky130_fd_sc_hd__a22o_1 _16375_ (.A1(\cpuregs[15][23] ),
    .A2(_12885_),
    .B1(_12836_),
    .B2(_12886_),
    .X(_03494_));
 sky130_fd_sc_hd__a22o_1 _16376_ (.A1(\cpuregs[15][22] ),
    .A2(_12885_),
    .B1(_12838_),
    .B2(_12886_),
    .X(_03493_));
 sky130_fd_sc_hd__a22o_1 _16377_ (.A1(\cpuregs[15][21] ),
    .A2(_12885_),
    .B1(_12839_),
    .B2(_12886_),
    .X(_03492_));
 sky130_fd_sc_hd__a22o_1 _16378_ (.A1(\cpuregs[15][20] ),
    .A2(_12885_),
    .B1(_12840_),
    .B2(_12886_),
    .X(_03491_));
 sky130_fd_sc_hd__buf_1 _16379_ (.A(_12878_),
    .X(_12887_));
 sky130_fd_sc_hd__buf_1 _16380_ (.A(_12881_),
    .X(_12888_));
 sky130_fd_sc_hd__a22o_1 _16381_ (.A1(\cpuregs[15][19] ),
    .A2(_12887_),
    .B1(_12842_),
    .B2(_12888_),
    .X(_03490_));
 sky130_fd_sc_hd__a22o_1 _16382_ (.A1(\cpuregs[15][18] ),
    .A2(_12887_),
    .B1(_12844_),
    .B2(_12888_),
    .X(_03489_));
 sky130_fd_sc_hd__a22o_1 _16383_ (.A1(\cpuregs[15][17] ),
    .A2(_12887_),
    .B1(_12845_),
    .B2(_12888_),
    .X(_03488_));
 sky130_fd_sc_hd__a22o_1 _16384_ (.A1(\cpuregs[15][16] ),
    .A2(_12887_),
    .B1(_12846_),
    .B2(_12888_),
    .X(_03487_));
 sky130_fd_sc_hd__buf_2 _16385_ (.A(_12877_),
    .X(_12889_));
 sky130_fd_sc_hd__buf_1 _16386_ (.A(_12889_),
    .X(_12890_));
 sky130_fd_sc_hd__buf_2 _16387_ (.A(_12880_),
    .X(_12891_));
 sky130_fd_sc_hd__buf_1 _16388_ (.A(_12891_),
    .X(_12892_));
 sky130_fd_sc_hd__a22o_1 _16389_ (.A1(\cpuregs[15][15] ),
    .A2(_12890_),
    .B1(_12849_),
    .B2(_12892_),
    .X(_03486_));
 sky130_fd_sc_hd__a22o_1 _16390_ (.A1(\cpuregs[15][14] ),
    .A2(_12890_),
    .B1(_12852_),
    .B2(_12892_),
    .X(_03485_));
 sky130_fd_sc_hd__a22o_1 _16391_ (.A1(\cpuregs[15][13] ),
    .A2(_12890_),
    .B1(_12853_),
    .B2(_12892_),
    .X(_03484_));
 sky130_fd_sc_hd__a22o_1 _16392_ (.A1(\cpuregs[15][12] ),
    .A2(_12890_),
    .B1(_12854_),
    .B2(_12892_),
    .X(_03483_));
 sky130_fd_sc_hd__buf_1 _16393_ (.A(_12889_),
    .X(_12893_));
 sky130_fd_sc_hd__buf_1 _16394_ (.A(_12891_),
    .X(_12894_));
 sky130_fd_sc_hd__a22o_1 _16395_ (.A1(\cpuregs[15][11] ),
    .A2(_12893_),
    .B1(_12856_),
    .B2(_12894_),
    .X(_03482_));
 sky130_fd_sc_hd__a22o_1 _16396_ (.A1(\cpuregs[15][10] ),
    .A2(_12893_),
    .B1(_12858_),
    .B2(_12894_),
    .X(_03481_));
 sky130_fd_sc_hd__a22o_1 _16397_ (.A1(\cpuregs[15][9] ),
    .A2(_12893_),
    .B1(_12859_),
    .B2(_12894_),
    .X(_03480_));
 sky130_fd_sc_hd__a22o_1 _16398_ (.A1(\cpuregs[15][8] ),
    .A2(_12893_),
    .B1(_12860_),
    .B2(_12894_),
    .X(_03479_));
 sky130_fd_sc_hd__buf_1 _16399_ (.A(_12889_),
    .X(_12895_));
 sky130_fd_sc_hd__buf_1 _16400_ (.A(_12891_),
    .X(_12896_));
 sky130_fd_sc_hd__a22o_1 _16401_ (.A1(\cpuregs[15][7] ),
    .A2(_12895_),
    .B1(_12862_),
    .B2(_12896_),
    .X(_03478_));
 sky130_fd_sc_hd__a22o_1 _16402_ (.A1(\cpuregs[15][6] ),
    .A2(_12895_),
    .B1(_12864_),
    .B2(_12896_),
    .X(_03477_));
 sky130_fd_sc_hd__a22o_1 _16403_ (.A1(\cpuregs[15][5] ),
    .A2(_12895_),
    .B1(_12865_),
    .B2(_12896_),
    .X(_03476_));
 sky130_fd_sc_hd__a22o_1 _16404_ (.A1(\cpuregs[15][4] ),
    .A2(_12895_),
    .B1(_12866_),
    .B2(_12896_),
    .X(_03475_));
 sky130_fd_sc_hd__buf_1 _16405_ (.A(_12889_),
    .X(_12897_));
 sky130_fd_sc_hd__buf_1 _16406_ (.A(_12891_),
    .X(_12898_));
 sky130_fd_sc_hd__a22o_1 _16407_ (.A1(\cpuregs[15][3] ),
    .A2(_12897_),
    .B1(_12868_),
    .B2(_12898_),
    .X(_03474_));
 sky130_fd_sc_hd__a22o_1 _16408_ (.A1(\cpuregs[15][2] ),
    .A2(_12897_),
    .B1(_12870_),
    .B2(_12898_),
    .X(_03473_));
 sky130_fd_sc_hd__a22o_1 _16409_ (.A1(\cpuregs[15][1] ),
    .A2(_12897_),
    .B1(_12871_),
    .B2(_12898_),
    .X(_03472_));
 sky130_fd_sc_hd__a22o_1 _16410_ (.A1(\cpuregs[15][0] ),
    .A2(_12897_),
    .B1(_12872_),
    .B2(_12898_),
    .X(_03471_));
 sky130_fd_sc_hd__or2_2 _16411_ (.A(_12655_),
    .B(_12818_),
    .X(_12899_));
 sky130_fd_sc_hd__clkbuf_4 _16412_ (.A(_12899_),
    .X(_12900_));
 sky130_fd_sc_hd__buf_1 _16413_ (.A(_12900_),
    .X(_12901_));
 sky130_vsdinv _16414_ (.A(_12899_),
    .Y(_12902_));
 sky130_fd_sc_hd__clkbuf_4 _16415_ (.A(_12902_),
    .X(_12903_));
 sky130_fd_sc_hd__buf_1 _16416_ (.A(_12903_),
    .X(_12904_));
 sky130_fd_sc_hd__a22o_1 _16417_ (.A1(\cpuregs[11][31] ),
    .A2(_12901_),
    .B1(_12822_),
    .B2(_12904_),
    .X(_03470_));
 sky130_fd_sc_hd__a22o_1 _16418_ (.A1(\cpuregs[11][30] ),
    .A2(_12901_),
    .B1(_12826_),
    .B2(_12904_),
    .X(_03469_));
 sky130_fd_sc_hd__a22o_1 _16419_ (.A1(\cpuregs[11][29] ),
    .A2(_12901_),
    .B1(_12827_),
    .B2(_12904_),
    .X(_03468_));
 sky130_fd_sc_hd__a22o_1 _16420_ (.A1(\cpuregs[11][28] ),
    .A2(_12901_),
    .B1(_12828_),
    .B2(_12904_),
    .X(_03467_));
 sky130_fd_sc_hd__buf_1 _16421_ (.A(_12900_),
    .X(_12905_));
 sky130_fd_sc_hd__buf_1 _16422_ (.A(_12903_),
    .X(_12906_));
 sky130_fd_sc_hd__a22o_1 _16423_ (.A1(\cpuregs[11][27] ),
    .A2(_12905_),
    .B1(_12830_),
    .B2(_12906_),
    .X(_03466_));
 sky130_fd_sc_hd__a22o_1 _16424_ (.A1(\cpuregs[11][26] ),
    .A2(_12905_),
    .B1(_12832_),
    .B2(_12906_),
    .X(_03465_));
 sky130_fd_sc_hd__a22o_1 _16425_ (.A1(\cpuregs[11][25] ),
    .A2(_12905_),
    .B1(_12833_),
    .B2(_12906_),
    .X(_03464_));
 sky130_fd_sc_hd__a22o_1 _16426_ (.A1(\cpuregs[11][24] ),
    .A2(_12905_),
    .B1(_12834_),
    .B2(_12906_),
    .X(_03463_));
 sky130_fd_sc_hd__buf_1 _16427_ (.A(_12900_),
    .X(_12907_));
 sky130_fd_sc_hd__buf_1 _16428_ (.A(_12903_),
    .X(_12908_));
 sky130_fd_sc_hd__a22o_1 _16429_ (.A1(\cpuregs[11][23] ),
    .A2(_12907_),
    .B1(_12836_),
    .B2(_12908_),
    .X(_03462_));
 sky130_fd_sc_hd__a22o_1 _16430_ (.A1(\cpuregs[11][22] ),
    .A2(_12907_),
    .B1(_12838_),
    .B2(_12908_),
    .X(_03461_));
 sky130_fd_sc_hd__a22o_1 _16431_ (.A1(\cpuregs[11][21] ),
    .A2(_12907_),
    .B1(_12839_),
    .B2(_12908_),
    .X(_03460_));
 sky130_fd_sc_hd__a22o_1 _16432_ (.A1(\cpuregs[11][20] ),
    .A2(_12907_),
    .B1(_12840_),
    .B2(_12908_),
    .X(_03459_));
 sky130_fd_sc_hd__buf_1 _16433_ (.A(_12900_),
    .X(_12909_));
 sky130_fd_sc_hd__buf_1 _16434_ (.A(_12903_),
    .X(_12910_));
 sky130_fd_sc_hd__a22o_1 _16435_ (.A1(\cpuregs[11][19] ),
    .A2(_12909_),
    .B1(_12842_),
    .B2(_12910_),
    .X(_03458_));
 sky130_fd_sc_hd__a22o_1 _16436_ (.A1(\cpuregs[11][18] ),
    .A2(_12909_),
    .B1(_12844_),
    .B2(_12910_),
    .X(_03457_));
 sky130_fd_sc_hd__a22o_1 _16437_ (.A1(\cpuregs[11][17] ),
    .A2(_12909_),
    .B1(_12845_),
    .B2(_12910_),
    .X(_03456_));
 sky130_fd_sc_hd__a22o_1 _16438_ (.A1(\cpuregs[11][16] ),
    .A2(_12909_),
    .B1(_12846_),
    .B2(_12910_),
    .X(_03455_));
 sky130_fd_sc_hd__clkbuf_2 _16439_ (.A(_12899_),
    .X(_12911_));
 sky130_fd_sc_hd__buf_1 _16440_ (.A(_12911_),
    .X(_12912_));
 sky130_fd_sc_hd__clkbuf_2 _16441_ (.A(_12902_),
    .X(_12913_));
 sky130_fd_sc_hd__buf_1 _16442_ (.A(_12913_),
    .X(_12914_));
 sky130_fd_sc_hd__a22o_1 _16443_ (.A1(\cpuregs[11][15] ),
    .A2(_12912_),
    .B1(_12849_),
    .B2(_12914_),
    .X(_03454_));
 sky130_fd_sc_hd__a22o_1 _16444_ (.A1(\cpuregs[11][14] ),
    .A2(_12912_),
    .B1(_12852_),
    .B2(_12914_),
    .X(_03453_));
 sky130_fd_sc_hd__a22o_1 _16445_ (.A1(\cpuregs[11][13] ),
    .A2(_12912_),
    .B1(_12853_),
    .B2(_12914_),
    .X(_03452_));
 sky130_fd_sc_hd__a22o_1 _16446_ (.A1(\cpuregs[11][12] ),
    .A2(_12912_),
    .B1(_12854_),
    .B2(_12914_),
    .X(_03451_));
 sky130_fd_sc_hd__clkbuf_2 _16447_ (.A(_12911_),
    .X(_12915_));
 sky130_fd_sc_hd__clkbuf_2 _16448_ (.A(_12913_),
    .X(_12916_));
 sky130_fd_sc_hd__a22o_1 _16449_ (.A1(\cpuregs[11][11] ),
    .A2(_12915_),
    .B1(_12856_),
    .B2(_12916_),
    .X(_03450_));
 sky130_fd_sc_hd__a22o_1 _16450_ (.A1(\cpuregs[11][10] ),
    .A2(_12915_),
    .B1(_12858_),
    .B2(_12916_),
    .X(_03449_));
 sky130_fd_sc_hd__a22o_1 _16451_ (.A1(\cpuregs[11][9] ),
    .A2(_12915_),
    .B1(_12859_),
    .B2(_12916_),
    .X(_03448_));
 sky130_fd_sc_hd__a22o_1 _16452_ (.A1(\cpuregs[11][8] ),
    .A2(_12915_),
    .B1(_12860_),
    .B2(_12916_),
    .X(_03447_));
 sky130_fd_sc_hd__buf_1 _16453_ (.A(_12911_),
    .X(_12917_));
 sky130_fd_sc_hd__buf_1 _16454_ (.A(_12913_),
    .X(_12918_));
 sky130_fd_sc_hd__a22o_1 _16455_ (.A1(\cpuregs[11][7] ),
    .A2(_12917_),
    .B1(_12862_),
    .B2(_12918_),
    .X(_03446_));
 sky130_fd_sc_hd__a22o_1 _16456_ (.A1(\cpuregs[11][6] ),
    .A2(_12917_),
    .B1(_12864_),
    .B2(_12918_),
    .X(_03445_));
 sky130_fd_sc_hd__a22o_1 _16457_ (.A1(\cpuregs[11][5] ),
    .A2(_12917_),
    .B1(_12865_),
    .B2(_12918_),
    .X(_03444_));
 sky130_fd_sc_hd__a22o_1 _16458_ (.A1(\cpuregs[11][4] ),
    .A2(_12917_),
    .B1(_12866_),
    .B2(_12918_),
    .X(_03443_));
 sky130_fd_sc_hd__buf_1 _16459_ (.A(_12911_),
    .X(_12919_));
 sky130_fd_sc_hd__buf_1 _16460_ (.A(_12913_),
    .X(_12920_));
 sky130_fd_sc_hd__a22o_1 _16461_ (.A1(\cpuregs[11][3] ),
    .A2(_12919_),
    .B1(_12868_),
    .B2(_12920_),
    .X(_03442_));
 sky130_fd_sc_hd__a22o_1 _16462_ (.A1(\cpuregs[11][2] ),
    .A2(_12919_),
    .B1(_12870_),
    .B2(_12920_),
    .X(_03441_));
 sky130_fd_sc_hd__a22o_1 _16463_ (.A1(\cpuregs[11][1] ),
    .A2(_12919_),
    .B1(_12871_),
    .B2(_12920_),
    .X(_03440_));
 sky130_fd_sc_hd__a22o_1 _16464_ (.A1(\cpuregs[11][0] ),
    .A2(_12919_),
    .B1(_12872_),
    .B2(_12920_),
    .X(_03439_));
 sky130_fd_sc_hd__or2_1 _16465_ (.A(_12561_),
    .B(_12818_),
    .X(_12921_));
 sky130_fd_sc_hd__buf_4 _16466_ (.A(_12921_),
    .X(_12922_));
 sky130_fd_sc_hd__buf_1 _16467_ (.A(_12922_),
    .X(_12923_));
 sky130_vsdinv _16468_ (.A(_12921_),
    .Y(_12924_));
 sky130_fd_sc_hd__buf_4 _16469_ (.A(_12924_),
    .X(_12925_));
 sky130_fd_sc_hd__buf_1 _16470_ (.A(_12925_),
    .X(_12926_));
 sky130_fd_sc_hd__a22o_1 _16471_ (.A1(\cpuregs[3][31] ),
    .A2(_12923_),
    .B1(_12822_),
    .B2(_12926_),
    .X(_03438_));
 sky130_fd_sc_hd__a22o_1 _16472_ (.A1(\cpuregs[3][30] ),
    .A2(_12923_),
    .B1(_12826_),
    .B2(_12926_),
    .X(_03437_));
 sky130_fd_sc_hd__a22o_1 _16473_ (.A1(\cpuregs[3][29] ),
    .A2(_12923_),
    .B1(_12827_),
    .B2(_12926_),
    .X(_03436_));
 sky130_fd_sc_hd__a22o_1 _16474_ (.A1(\cpuregs[3][28] ),
    .A2(_12923_),
    .B1(_12828_),
    .B2(_12926_),
    .X(_03435_));
 sky130_fd_sc_hd__buf_1 _16475_ (.A(_12922_),
    .X(_12927_));
 sky130_fd_sc_hd__buf_1 _16476_ (.A(_12925_),
    .X(_12928_));
 sky130_fd_sc_hd__a22o_1 _16477_ (.A1(\cpuregs[3][27] ),
    .A2(_12927_),
    .B1(_12830_),
    .B2(_12928_),
    .X(_03434_));
 sky130_fd_sc_hd__a22o_1 _16478_ (.A1(\cpuregs[3][26] ),
    .A2(_12927_),
    .B1(_12832_),
    .B2(_12928_),
    .X(_03433_));
 sky130_fd_sc_hd__a22o_1 _16479_ (.A1(\cpuregs[3][25] ),
    .A2(_12927_),
    .B1(_12833_),
    .B2(_12928_),
    .X(_03432_));
 sky130_fd_sc_hd__a22o_1 _16480_ (.A1(\cpuregs[3][24] ),
    .A2(_12927_),
    .B1(_12834_),
    .B2(_12928_),
    .X(_03431_));
 sky130_fd_sc_hd__buf_1 _16481_ (.A(_12922_),
    .X(_12929_));
 sky130_fd_sc_hd__buf_1 _16482_ (.A(_12925_),
    .X(_12930_));
 sky130_fd_sc_hd__a22o_1 _16483_ (.A1(\cpuregs[3][23] ),
    .A2(_12929_),
    .B1(_12836_),
    .B2(_12930_),
    .X(_03430_));
 sky130_fd_sc_hd__a22o_1 _16484_ (.A1(\cpuregs[3][22] ),
    .A2(_12929_),
    .B1(_12838_),
    .B2(_12930_),
    .X(_03429_));
 sky130_fd_sc_hd__a22o_1 _16485_ (.A1(\cpuregs[3][21] ),
    .A2(_12929_),
    .B1(_12839_),
    .B2(_12930_),
    .X(_03428_));
 sky130_fd_sc_hd__a22o_1 _16486_ (.A1(\cpuregs[3][20] ),
    .A2(_12929_),
    .B1(_12840_),
    .B2(_12930_),
    .X(_03427_));
 sky130_fd_sc_hd__buf_1 _16487_ (.A(_12922_),
    .X(_12931_));
 sky130_fd_sc_hd__buf_1 _16488_ (.A(_12925_),
    .X(_12932_));
 sky130_fd_sc_hd__a22o_1 _16489_ (.A1(\cpuregs[3][19] ),
    .A2(_12931_),
    .B1(_12842_),
    .B2(_12932_),
    .X(_03426_));
 sky130_fd_sc_hd__a22o_1 _16490_ (.A1(\cpuregs[3][18] ),
    .A2(_12931_),
    .B1(_12844_),
    .B2(_12932_),
    .X(_03425_));
 sky130_fd_sc_hd__a22o_1 _16491_ (.A1(\cpuregs[3][17] ),
    .A2(_12931_),
    .B1(_12845_),
    .B2(_12932_),
    .X(_03424_));
 sky130_fd_sc_hd__a22o_1 _16492_ (.A1(\cpuregs[3][16] ),
    .A2(_12931_),
    .B1(_12846_),
    .B2(_12932_),
    .X(_03423_));
 sky130_fd_sc_hd__clkbuf_4 _16493_ (.A(_12921_),
    .X(_12933_));
 sky130_fd_sc_hd__buf_1 _16494_ (.A(_12933_),
    .X(_12934_));
 sky130_fd_sc_hd__clkbuf_4 _16495_ (.A(_12924_),
    .X(_12935_));
 sky130_fd_sc_hd__buf_1 _16496_ (.A(_12935_),
    .X(_12936_));
 sky130_fd_sc_hd__a22o_1 _16497_ (.A1(\cpuregs[3][15] ),
    .A2(_12934_),
    .B1(_12849_),
    .B2(_12936_),
    .X(_03422_));
 sky130_fd_sc_hd__a22o_1 _16498_ (.A1(\cpuregs[3][14] ),
    .A2(_12934_),
    .B1(_12852_),
    .B2(_12936_),
    .X(_03421_));
 sky130_fd_sc_hd__a22o_1 _16499_ (.A1(\cpuregs[3][13] ),
    .A2(_12934_),
    .B1(_12853_),
    .B2(_12936_),
    .X(_03420_));
 sky130_fd_sc_hd__a22o_1 _16500_ (.A1(\cpuregs[3][12] ),
    .A2(_12934_),
    .B1(_12854_),
    .B2(_12936_),
    .X(_03419_));
 sky130_fd_sc_hd__buf_1 _16501_ (.A(_12933_),
    .X(_12937_));
 sky130_fd_sc_hd__buf_1 _16502_ (.A(_12935_),
    .X(_12938_));
 sky130_fd_sc_hd__a22o_1 _16503_ (.A1(\cpuregs[3][11] ),
    .A2(_12937_),
    .B1(_12856_),
    .B2(_12938_),
    .X(_03418_));
 sky130_fd_sc_hd__a22o_1 _16504_ (.A1(\cpuregs[3][10] ),
    .A2(_12937_),
    .B1(_12858_),
    .B2(_12938_),
    .X(_03417_));
 sky130_fd_sc_hd__a22o_1 _16505_ (.A1(\cpuregs[3][9] ),
    .A2(_12937_),
    .B1(_12859_),
    .B2(_12938_),
    .X(_03416_));
 sky130_fd_sc_hd__a22o_1 _16506_ (.A1(\cpuregs[3][8] ),
    .A2(_12937_),
    .B1(_12860_),
    .B2(_12938_),
    .X(_03415_));
 sky130_fd_sc_hd__buf_1 _16507_ (.A(_12933_),
    .X(_12939_));
 sky130_fd_sc_hd__buf_1 _16508_ (.A(_12935_),
    .X(_12940_));
 sky130_fd_sc_hd__a22o_1 _16509_ (.A1(\cpuregs[3][7] ),
    .A2(_12939_),
    .B1(_12862_),
    .B2(_12940_),
    .X(_03414_));
 sky130_fd_sc_hd__a22o_1 _16510_ (.A1(\cpuregs[3][6] ),
    .A2(_12939_),
    .B1(_12864_),
    .B2(_12940_),
    .X(_03413_));
 sky130_fd_sc_hd__a22o_1 _16511_ (.A1(\cpuregs[3][5] ),
    .A2(_12939_),
    .B1(_12865_),
    .B2(_12940_),
    .X(_03412_));
 sky130_fd_sc_hd__a22o_1 _16512_ (.A1(\cpuregs[3][4] ),
    .A2(_12939_),
    .B1(_12866_),
    .B2(_12940_),
    .X(_03411_));
 sky130_fd_sc_hd__buf_1 _16513_ (.A(_12933_),
    .X(_12941_));
 sky130_fd_sc_hd__buf_1 _16514_ (.A(_12935_),
    .X(_12942_));
 sky130_fd_sc_hd__a22o_1 _16515_ (.A1(\cpuregs[3][3] ),
    .A2(_12941_),
    .B1(_12868_),
    .B2(_12942_),
    .X(_03410_));
 sky130_fd_sc_hd__a22o_1 _16516_ (.A1(\cpuregs[3][2] ),
    .A2(_12941_),
    .B1(_12870_),
    .B2(_12942_),
    .X(_03409_));
 sky130_fd_sc_hd__a22o_1 _16517_ (.A1(\cpuregs[3][1] ),
    .A2(_12941_),
    .B1(_12871_),
    .B2(_12942_),
    .X(_03408_));
 sky130_fd_sc_hd__a22o_1 _16518_ (.A1(\cpuregs[3][0] ),
    .A2(_12941_),
    .B1(_12872_),
    .B2(_12942_),
    .X(_03407_));
 sky130_fd_sc_hd__or2_2 _16519_ (.A(_12561_),
    .B(_12658_),
    .X(_12943_));
 sky130_fd_sc_hd__buf_4 _16520_ (.A(_12943_),
    .X(_12944_));
 sky130_fd_sc_hd__buf_1 _16521_ (.A(_12944_),
    .X(_12945_));
 sky130_fd_sc_hd__clkbuf_2 _16522_ (.A(\cpuregs_wrdata[31] ),
    .X(_12946_));
 sky130_vsdinv _16523_ (.A(_12943_),
    .Y(_12947_));
 sky130_fd_sc_hd__buf_4 _16524_ (.A(_12947_),
    .X(_12948_));
 sky130_fd_sc_hd__buf_1 _16525_ (.A(_12948_),
    .X(_12949_));
 sky130_fd_sc_hd__a22o_1 _16526_ (.A1(\cpuregs[1][31] ),
    .A2(_12945_),
    .B1(_12946_),
    .B2(_12949_),
    .X(_03406_));
 sky130_fd_sc_hd__clkbuf_2 _16527_ (.A(\cpuregs_wrdata[30] ),
    .X(_12950_));
 sky130_fd_sc_hd__a22o_1 _16528_ (.A1(\cpuregs[1][30] ),
    .A2(_12945_),
    .B1(_12950_),
    .B2(_12949_),
    .X(_03405_));
 sky130_fd_sc_hd__clkbuf_2 _16529_ (.A(\cpuregs_wrdata[29] ),
    .X(_12951_));
 sky130_fd_sc_hd__a22o_1 _16530_ (.A1(\cpuregs[1][29] ),
    .A2(_12945_),
    .B1(_12951_),
    .B2(_12949_),
    .X(_03404_));
 sky130_fd_sc_hd__clkbuf_2 _16531_ (.A(\cpuregs_wrdata[28] ),
    .X(_12952_));
 sky130_fd_sc_hd__a22o_1 _16532_ (.A1(\cpuregs[1][28] ),
    .A2(_12945_),
    .B1(_12952_),
    .B2(_12949_),
    .X(_03403_));
 sky130_fd_sc_hd__buf_1 _16533_ (.A(_12944_),
    .X(_12953_));
 sky130_fd_sc_hd__clkbuf_2 _16534_ (.A(\cpuregs_wrdata[27] ),
    .X(_12954_));
 sky130_fd_sc_hd__buf_1 _16535_ (.A(_12948_),
    .X(_12955_));
 sky130_fd_sc_hd__a22o_1 _16536_ (.A1(\cpuregs[1][27] ),
    .A2(_12953_),
    .B1(_12954_),
    .B2(_12955_),
    .X(_03402_));
 sky130_fd_sc_hd__clkbuf_2 _16537_ (.A(\cpuregs_wrdata[26] ),
    .X(_12956_));
 sky130_fd_sc_hd__a22o_1 _16538_ (.A1(\cpuregs[1][26] ),
    .A2(_12953_),
    .B1(_12956_),
    .B2(_12955_),
    .X(_03401_));
 sky130_fd_sc_hd__clkbuf_2 _16539_ (.A(\cpuregs_wrdata[25] ),
    .X(_12957_));
 sky130_fd_sc_hd__a22o_1 _16540_ (.A1(\cpuregs[1][25] ),
    .A2(_12953_),
    .B1(_12957_),
    .B2(_12955_),
    .X(_03400_));
 sky130_fd_sc_hd__clkbuf_2 _16541_ (.A(\cpuregs_wrdata[24] ),
    .X(_12958_));
 sky130_fd_sc_hd__a22o_1 _16542_ (.A1(\cpuregs[1][24] ),
    .A2(_12953_),
    .B1(_12958_),
    .B2(_12955_),
    .X(_03399_));
 sky130_fd_sc_hd__buf_1 _16543_ (.A(_12944_),
    .X(_12959_));
 sky130_fd_sc_hd__clkbuf_2 _16544_ (.A(\cpuregs_wrdata[23] ),
    .X(_12960_));
 sky130_fd_sc_hd__buf_1 _16545_ (.A(_12948_),
    .X(_12961_));
 sky130_fd_sc_hd__a22o_1 _16546_ (.A1(\cpuregs[1][23] ),
    .A2(_12959_),
    .B1(_12960_),
    .B2(_12961_),
    .X(_03398_));
 sky130_fd_sc_hd__clkbuf_2 _16547_ (.A(\cpuregs_wrdata[22] ),
    .X(_12962_));
 sky130_fd_sc_hd__a22o_1 _16548_ (.A1(\cpuregs[1][22] ),
    .A2(_12959_),
    .B1(_12962_),
    .B2(_12961_),
    .X(_03397_));
 sky130_fd_sc_hd__clkbuf_2 _16549_ (.A(\cpuregs_wrdata[21] ),
    .X(_12963_));
 sky130_fd_sc_hd__a22o_1 _16550_ (.A1(\cpuregs[1][21] ),
    .A2(_12959_),
    .B1(_12963_),
    .B2(_12961_),
    .X(_03396_));
 sky130_fd_sc_hd__clkbuf_2 _16551_ (.A(\cpuregs_wrdata[20] ),
    .X(_12964_));
 sky130_fd_sc_hd__a22o_1 _16552_ (.A1(\cpuregs[1][20] ),
    .A2(_12959_),
    .B1(_12964_),
    .B2(_12961_),
    .X(_03395_));
 sky130_fd_sc_hd__buf_1 _16553_ (.A(_12944_),
    .X(_12965_));
 sky130_fd_sc_hd__clkbuf_2 _16554_ (.A(\cpuregs_wrdata[19] ),
    .X(_12966_));
 sky130_fd_sc_hd__buf_1 _16555_ (.A(_12948_),
    .X(_12967_));
 sky130_fd_sc_hd__a22o_1 _16556_ (.A1(\cpuregs[1][19] ),
    .A2(_12965_),
    .B1(_12966_),
    .B2(_12967_),
    .X(_03394_));
 sky130_fd_sc_hd__clkbuf_2 _16557_ (.A(\cpuregs_wrdata[18] ),
    .X(_12968_));
 sky130_fd_sc_hd__a22o_1 _16558_ (.A1(\cpuregs[1][18] ),
    .A2(_12965_),
    .B1(_12968_),
    .B2(_12967_),
    .X(_03393_));
 sky130_fd_sc_hd__clkbuf_2 _16559_ (.A(\cpuregs_wrdata[17] ),
    .X(_12969_));
 sky130_fd_sc_hd__a22o_1 _16560_ (.A1(\cpuregs[1][17] ),
    .A2(_12965_),
    .B1(_12969_),
    .B2(_12967_),
    .X(_03392_));
 sky130_fd_sc_hd__clkbuf_2 _16561_ (.A(\cpuregs_wrdata[16] ),
    .X(_12970_));
 sky130_fd_sc_hd__a22o_1 _16562_ (.A1(\cpuregs[1][16] ),
    .A2(_12965_),
    .B1(_12970_),
    .B2(_12967_),
    .X(_03391_));
 sky130_fd_sc_hd__clkbuf_4 _16563_ (.A(_12943_),
    .X(_12971_));
 sky130_fd_sc_hd__buf_1 _16564_ (.A(_12971_),
    .X(_12972_));
 sky130_fd_sc_hd__clkbuf_2 _16565_ (.A(\cpuregs_wrdata[15] ),
    .X(_12973_));
 sky130_fd_sc_hd__clkbuf_4 _16566_ (.A(_12947_),
    .X(_12974_));
 sky130_fd_sc_hd__buf_1 _16567_ (.A(_12974_),
    .X(_12975_));
 sky130_fd_sc_hd__a22o_1 _16568_ (.A1(\cpuregs[1][15] ),
    .A2(_12972_),
    .B1(_12973_),
    .B2(_12975_),
    .X(_03390_));
 sky130_fd_sc_hd__clkbuf_2 _16569_ (.A(\cpuregs_wrdata[14] ),
    .X(_12976_));
 sky130_fd_sc_hd__a22o_1 _16570_ (.A1(\cpuregs[1][14] ),
    .A2(_12972_),
    .B1(_12976_),
    .B2(_12975_),
    .X(_03389_));
 sky130_fd_sc_hd__buf_1 _16571_ (.A(\cpuregs_wrdata[13] ),
    .X(_12977_));
 sky130_fd_sc_hd__a22o_1 _16572_ (.A1(\cpuregs[1][13] ),
    .A2(_12972_),
    .B1(_12977_),
    .B2(_12975_),
    .X(_03388_));
 sky130_fd_sc_hd__clkbuf_2 _16573_ (.A(\cpuregs_wrdata[12] ),
    .X(_12978_));
 sky130_fd_sc_hd__a22o_1 _16574_ (.A1(\cpuregs[1][12] ),
    .A2(_12972_),
    .B1(_12978_),
    .B2(_12975_),
    .X(_03387_));
 sky130_fd_sc_hd__buf_1 _16575_ (.A(_12971_),
    .X(_12979_));
 sky130_fd_sc_hd__buf_1 _16576_ (.A(\cpuregs_wrdata[11] ),
    .X(_12980_));
 sky130_fd_sc_hd__buf_1 _16577_ (.A(_12974_),
    .X(_12981_));
 sky130_fd_sc_hd__a22o_1 _16578_ (.A1(\cpuregs[1][11] ),
    .A2(_12979_),
    .B1(_12980_),
    .B2(_12981_),
    .X(_03386_));
 sky130_fd_sc_hd__buf_1 _16579_ (.A(\cpuregs_wrdata[10] ),
    .X(_12982_));
 sky130_fd_sc_hd__a22o_1 _16580_ (.A1(\cpuregs[1][10] ),
    .A2(_12979_),
    .B1(_12982_),
    .B2(_12981_),
    .X(_03385_));
 sky130_fd_sc_hd__buf_1 _16581_ (.A(\cpuregs_wrdata[9] ),
    .X(_12983_));
 sky130_fd_sc_hd__a22o_1 _16582_ (.A1(\cpuregs[1][9] ),
    .A2(_12979_),
    .B1(_12983_),
    .B2(_12981_),
    .X(_03384_));
 sky130_fd_sc_hd__buf_1 _16583_ (.A(\cpuregs_wrdata[8] ),
    .X(_12984_));
 sky130_fd_sc_hd__a22o_1 _16584_ (.A1(\cpuregs[1][8] ),
    .A2(_12979_),
    .B1(_12984_),
    .B2(_12981_),
    .X(_03383_));
 sky130_fd_sc_hd__buf_1 _16585_ (.A(_12971_),
    .X(_12985_));
 sky130_fd_sc_hd__clkbuf_2 _16586_ (.A(\cpuregs_wrdata[7] ),
    .X(_12986_));
 sky130_fd_sc_hd__buf_1 _16587_ (.A(_12974_),
    .X(_12987_));
 sky130_fd_sc_hd__a22o_1 _16588_ (.A1(\cpuregs[1][7] ),
    .A2(_12985_),
    .B1(_12986_),
    .B2(_12987_),
    .X(_03382_));
 sky130_fd_sc_hd__buf_1 _16589_ (.A(\cpuregs_wrdata[6] ),
    .X(_12988_));
 sky130_fd_sc_hd__a22o_1 _16590_ (.A1(\cpuregs[1][6] ),
    .A2(_12985_),
    .B1(_12988_),
    .B2(_12987_),
    .X(_03381_));
 sky130_fd_sc_hd__clkbuf_2 _16591_ (.A(\cpuregs_wrdata[5] ),
    .X(_12989_));
 sky130_fd_sc_hd__a22o_1 _16592_ (.A1(\cpuregs[1][5] ),
    .A2(_12985_),
    .B1(_12989_),
    .B2(_12987_),
    .X(_03380_));
 sky130_fd_sc_hd__clkbuf_2 _16593_ (.A(\cpuregs_wrdata[4] ),
    .X(_12990_));
 sky130_fd_sc_hd__a22o_1 _16594_ (.A1(\cpuregs[1][4] ),
    .A2(_12985_),
    .B1(_12990_),
    .B2(_12987_),
    .X(_03379_));
 sky130_fd_sc_hd__buf_1 _16595_ (.A(_12971_),
    .X(_12991_));
 sky130_fd_sc_hd__clkbuf_2 _16596_ (.A(\cpuregs_wrdata[3] ),
    .X(_12992_));
 sky130_fd_sc_hd__buf_1 _16597_ (.A(_12974_),
    .X(_12993_));
 sky130_fd_sc_hd__a22o_1 _16598_ (.A1(\cpuregs[1][3] ),
    .A2(_12991_),
    .B1(_12992_),
    .B2(_12993_),
    .X(_03378_));
 sky130_fd_sc_hd__clkbuf_2 _16599_ (.A(\cpuregs_wrdata[2] ),
    .X(_12994_));
 sky130_fd_sc_hd__a22o_1 _16600_ (.A1(\cpuregs[1][2] ),
    .A2(_12991_),
    .B1(_12994_),
    .B2(_12993_),
    .X(_03377_));
 sky130_fd_sc_hd__clkbuf_2 _16601_ (.A(\cpuregs_wrdata[1] ),
    .X(_12995_));
 sky130_fd_sc_hd__a22o_1 _16602_ (.A1(\cpuregs[1][1] ),
    .A2(_12991_),
    .B1(_12995_),
    .B2(_12993_),
    .X(_03376_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _16603_ (.A(\cpuregs_wrdata[0] ),
    .X(_12996_));
 sky130_fd_sc_hd__a22o_1 _16604_ (.A1(\cpuregs[1][0] ),
    .A2(_12991_),
    .B1(_12996_),
    .B2(_12993_),
    .X(_03375_));
 sky130_fd_sc_hd__or2_1 _16605_ (.A(_12746_),
    .B(_12876_),
    .X(_12997_));
 sky130_fd_sc_hd__buf_4 _16606_ (.A(_12997_),
    .X(_12998_));
 sky130_fd_sc_hd__buf_1 _16607_ (.A(_12998_),
    .X(_12999_));
 sky130_vsdinv _16608_ (.A(_12997_),
    .Y(_13000_));
 sky130_fd_sc_hd__buf_4 _16609_ (.A(_13000_),
    .X(_13001_));
 sky130_fd_sc_hd__buf_1 _16610_ (.A(_13001_),
    .X(_13002_));
 sky130_fd_sc_hd__a22o_1 _16611_ (.A1(\cpuregs[12][31] ),
    .A2(_12999_),
    .B1(_12946_),
    .B2(_13002_),
    .X(_03374_));
 sky130_fd_sc_hd__a22o_1 _16612_ (.A1(\cpuregs[12][30] ),
    .A2(_12999_),
    .B1(_12950_),
    .B2(_13002_),
    .X(_03373_));
 sky130_fd_sc_hd__a22o_1 _16613_ (.A1(\cpuregs[12][29] ),
    .A2(_12999_),
    .B1(_12951_),
    .B2(_13002_),
    .X(_03372_));
 sky130_fd_sc_hd__a22o_1 _16614_ (.A1(\cpuregs[12][28] ),
    .A2(_12999_),
    .B1(_12952_),
    .B2(_13002_),
    .X(_03371_));
 sky130_fd_sc_hd__buf_1 _16615_ (.A(_12998_),
    .X(_13003_));
 sky130_fd_sc_hd__buf_1 _16616_ (.A(_13001_),
    .X(_13004_));
 sky130_fd_sc_hd__a22o_1 _16617_ (.A1(\cpuregs[12][27] ),
    .A2(_13003_),
    .B1(_12954_),
    .B2(_13004_),
    .X(_03370_));
 sky130_fd_sc_hd__a22o_1 _16618_ (.A1(\cpuregs[12][26] ),
    .A2(_13003_),
    .B1(_12956_),
    .B2(_13004_),
    .X(_03369_));
 sky130_fd_sc_hd__a22o_1 _16619_ (.A1(\cpuregs[12][25] ),
    .A2(_13003_),
    .B1(_12957_),
    .B2(_13004_),
    .X(_03368_));
 sky130_fd_sc_hd__a22o_1 _16620_ (.A1(\cpuregs[12][24] ),
    .A2(_13003_),
    .B1(_12958_),
    .B2(_13004_),
    .X(_03367_));
 sky130_fd_sc_hd__buf_1 _16621_ (.A(_12998_),
    .X(_13005_));
 sky130_fd_sc_hd__buf_1 _16622_ (.A(_13001_),
    .X(_13006_));
 sky130_fd_sc_hd__a22o_1 _16623_ (.A1(\cpuregs[12][23] ),
    .A2(_13005_),
    .B1(_12960_),
    .B2(_13006_),
    .X(_03366_));
 sky130_fd_sc_hd__a22o_1 _16624_ (.A1(\cpuregs[12][22] ),
    .A2(_13005_),
    .B1(_12962_),
    .B2(_13006_),
    .X(_03365_));
 sky130_fd_sc_hd__a22o_1 _16625_ (.A1(\cpuregs[12][21] ),
    .A2(_13005_),
    .B1(_12963_),
    .B2(_13006_),
    .X(_03364_));
 sky130_fd_sc_hd__a22o_1 _16626_ (.A1(\cpuregs[12][20] ),
    .A2(_13005_),
    .B1(_12964_),
    .B2(_13006_),
    .X(_03363_));
 sky130_fd_sc_hd__buf_1 _16627_ (.A(_12998_),
    .X(_13007_));
 sky130_fd_sc_hd__buf_1 _16628_ (.A(_13001_),
    .X(_13008_));
 sky130_fd_sc_hd__a22o_1 _16629_ (.A1(\cpuregs[12][19] ),
    .A2(_13007_),
    .B1(_12966_),
    .B2(_13008_),
    .X(_03362_));
 sky130_fd_sc_hd__a22o_1 _16630_ (.A1(\cpuregs[12][18] ),
    .A2(_13007_),
    .B1(_12968_),
    .B2(_13008_),
    .X(_03361_));
 sky130_fd_sc_hd__a22o_1 _16631_ (.A1(\cpuregs[12][17] ),
    .A2(_13007_),
    .B1(_12969_),
    .B2(_13008_),
    .X(_03360_));
 sky130_fd_sc_hd__a22o_1 _16632_ (.A1(\cpuregs[12][16] ),
    .A2(_13007_),
    .B1(_12970_),
    .B2(_13008_),
    .X(_03359_));
 sky130_fd_sc_hd__buf_2 _16633_ (.A(_12997_),
    .X(_13009_));
 sky130_fd_sc_hd__buf_1 _16634_ (.A(_13009_),
    .X(_13010_));
 sky130_fd_sc_hd__buf_2 _16635_ (.A(_13000_),
    .X(_13011_));
 sky130_fd_sc_hd__buf_1 _16636_ (.A(_13011_),
    .X(_13012_));
 sky130_fd_sc_hd__a22o_1 _16637_ (.A1(\cpuregs[12][15] ),
    .A2(_13010_),
    .B1(_12973_),
    .B2(_13012_),
    .X(_03358_));
 sky130_fd_sc_hd__a22o_1 _16638_ (.A1(\cpuregs[12][14] ),
    .A2(_13010_),
    .B1(_12976_),
    .B2(_13012_),
    .X(_03357_));
 sky130_fd_sc_hd__a22o_1 _16639_ (.A1(\cpuregs[12][13] ),
    .A2(_13010_),
    .B1(_12977_),
    .B2(_13012_),
    .X(_03356_));
 sky130_fd_sc_hd__a22o_1 _16640_ (.A1(\cpuregs[12][12] ),
    .A2(_13010_),
    .B1(_12978_),
    .B2(_13012_),
    .X(_03355_));
 sky130_fd_sc_hd__buf_1 _16641_ (.A(_13009_),
    .X(_13013_));
 sky130_fd_sc_hd__buf_1 _16642_ (.A(_13011_),
    .X(_13014_));
 sky130_fd_sc_hd__a22o_1 _16643_ (.A1(\cpuregs[12][11] ),
    .A2(_13013_),
    .B1(_12980_),
    .B2(_13014_),
    .X(_03354_));
 sky130_fd_sc_hd__a22o_1 _16644_ (.A1(\cpuregs[12][10] ),
    .A2(_13013_),
    .B1(_12982_),
    .B2(_13014_),
    .X(_03353_));
 sky130_fd_sc_hd__a22o_1 _16645_ (.A1(\cpuregs[12][9] ),
    .A2(_13013_),
    .B1(_12983_),
    .B2(_13014_),
    .X(_03352_));
 sky130_fd_sc_hd__a22o_1 _16646_ (.A1(\cpuregs[12][8] ),
    .A2(_13013_),
    .B1(_12984_),
    .B2(_13014_),
    .X(_03351_));
 sky130_fd_sc_hd__buf_1 _16647_ (.A(_13009_),
    .X(_13015_));
 sky130_fd_sc_hd__buf_1 _16648_ (.A(_13011_),
    .X(_13016_));
 sky130_fd_sc_hd__a22o_1 _16649_ (.A1(\cpuregs[12][7] ),
    .A2(_13015_),
    .B1(_12986_),
    .B2(_13016_),
    .X(_03350_));
 sky130_fd_sc_hd__a22o_1 _16650_ (.A1(\cpuregs[12][6] ),
    .A2(_13015_),
    .B1(_12988_),
    .B2(_13016_),
    .X(_03349_));
 sky130_fd_sc_hd__a22o_1 _16651_ (.A1(\cpuregs[12][5] ),
    .A2(_13015_),
    .B1(_12989_),
    .B2(_13016_),
    .X(_03348_));
 sky130_fd_sc_hd__a22o_1 _16652_ (.A1(\cpuregs[12][4] ),
    .A2(_13015_),
    .B1(_12990_),
    .B2(_13016_),
    .X(_03347_));
 sky130_fd_sc_hd__buf_1 _16653_ (.A(_13009_),
    .X(_13017_));
 sky130_fd_sc_hd__buf_1 _16654_ (.A(_13011_),
    .X(_13018_));
 sky130_fd_sc_hd__a22o_1 _16655_ (.A1(\cpuregs[12][3] ),
    .A2(_13017_),
    .B1(_12992_),
    .B2(_13018_),
    .X(_03346_));
 sky130_fd_sc_hd__a22o_1 _16656_ (.A1(\cpuregs[12][2] ),
    .A2(_13017_),
    .B1(_12994_),
    .B2(_13018_),
    .X(_03345_));
 sky130_fd_sc_hd__a22o_1 _16657_ (.A1(\cpuregs[12][1] ),
    .A2(_13017_),
    .B1(_12995_),
    .B2(_13018_),
    .X(_03344_));
 sky130_fd_sc_hd__a22o_1 _16658_ (.A1(\cpuregs[12][0] ),
    .A2(_13017_),
    .B1(_12996_),
    .B2(_13018_),
    .X(_03343_));
 sky130_fd_sc_hd__or3_4 _16659_ (.A(_12770_),
    .B(_12771_),
    .C(_12746_),
    .X(_13019_));
 sky130_fd_sc_hd__clkbuf_4 _16660_ (.A(_13019_),
    .X(_13020_));
 sky130_fd_sc_hd__buf_1 _16661_ (.A(_13020_),
    .X(_13021_));
 sky130_vsdinv _16662_ (.A(_13019_),
    .Y(_13022_));
 sky130_fd_sc_hd__clkbuf_4 _16663_ (.A(_13022_),
    .X(_13023_));
 sky130_fd_sc_hd__buf_1 _16664_ (.A(_13023_),
    .X(_13024_));
 sky130_fd_sc_hd__a22o_1 _16665_ (.A1(\cpuregs[16][31] ),
    .A2(_13021_),
    .B1(_12946_),
    .B2(_13024_),
    .X(_03342_));
 sky130_fd_sc_hd__a22o_1 _16666_ (.A1(\cpuregs[16][30] ),
    .A2(_13021_),
    .B1(_12950_),
    .B2(_13024_),
    .X(_03341_));
 sky130_fd_sc_hd__a22o_1 _16667_ (.A1(\cpuregs[16][29] ),
    .A2(_13021_),
    .B1(_12951_),
    .B2(_13024_),
    .X(_03340_));
 sky130_fd_sc_hd__a22o_1 _16668_ (.A1(\cpuregs[16][28] ),
    .A2(_13021_),
    .B1(_12952_),
    .B2(_13024_),
    .X(_03339_));
 sky130_fd_sc_hd__buf_1 _16669_ (.A(_13020_),
    .X(_13025_));
 sky130_fd_sc_hd__buf_1 _16670_ (.A(_13023_),
    .X(_13026_));
 sky130_fd_sc_hd__a22o_1 _16671_ (.A1(\cpuregs[16][27] ),
    .A2(_13025_),
    .B1(_12954_),
    .B2(_13026_),
    .X(_03338_));
 sky130_fd_sc_hd__a22o_1 _16672_ (.A1(\cpuregs[16][26] ),
    .A2(_13025_),
    .B1(_12956_),
    .B2(_13026_),
    .X(_03337_));
 sky130_fd_sc_hd__a22o_1 _16673_ (.A1(\cpuregs[16][25] ),
    .A2(_13025_),
    .B1(_12957_),
    .B2(_13026_),
    .X(_03336_));
 sky130_fd_sc_hd__a22o_1 _16674_ (.A1(\cpuregs[16][24] ),
    .A2(_13025_),
    .B1(_12958_),
    .B2(_13026_),
    .X(_03335_));
 sky130_fd_sc_hd__buf_1 _16675_ (.A(_13020_),
    .X(_13027_));
 sky130_fd_sc_hd__buf_1 _16676_ (.A(_13023_),
    .X(_13028_));
 sky130_fd_sc_hd__a22o_1 _16677_ (.A1(\cpuregs[16][23] ),
    .A2(_13027_),
    .B1(_12960_),
    .B2(_13028_),
    .X(_03334_));
 sky130_fd_sc_hd__a22o_1 _16678_ (.A1(\cpuregs[16][22] ),
    .A2(_13027_),
    .B1(_12962_),
    .B2(_13028_),
    .X(_03333_));
 sky130_fd_sc_hd__a22o_1 _16679_ (.A1(\cpuregs[16][21] ),
    .A2(_13027_),
    .B1(_12963_),
    .B2(_13028_),
    .X(_03332_));
 sky130_fd_sc_hd__a22o_1 _16680_ (.A1(\cpuregs[16][20] ),
    .A2(_13027_),
    .B1(_12964_),
    .B2(_13028_),
    .X(_03331_));
 sky130_fd_sc_hd__buf_1 _16681_ (.A(_13020_),
    .X(_13029_));
 sky130_fd_sc_hd__buf_1 _16682_ (.A(_13023_),
    .X(_13030_));
 sky130_fd_sc_hd__a22o_1 _16683_ (.A1(\cpuregs[16][19] ),
    .A2(_13029_),
    .B1(_12966_),
    .B2(_13030_),
    .X(_03330_));
 sky130_fd_sc_hd__a22o_1 _16684_ (.A1(\cpuregs[16][18] ),
    .A2(_13029_),
    .B1(_12968_),
    .B2(_13030_),
    .X(_03329_));
 sky130_fd_sc_hd__a22o_1 _16685_ (.A1(\cpuregs[16][17] ),
    .A2(_13029_),
    .B1(_12969_),
    .B2(_13030_),
    .X(_03328_));
 sky130_fd_sc_hd__a22o_1 _16686_ (.A1(\cpuregs[16][16] ),
    .A2(_13029_),
    .B1(_12970_),
    .B2(_13030_),
    .X(_03327_));
 sky130_fd_sc_hd__clkbuf_4 _16687_ (.A(_13019_),
    .X(_13031_));
 sky130_fd_sc_hd__buf_1 _16688_ (.A(_13031_),
    .X(_13032_));
 sky130_fd_sc_hd__clkbuf_4 _16689_ (.A(_13022_),
    .X(_13033_));
 sky130_fd_sc_hd__buf_1 _16690_ (.A(_13033_),
    .X(_13034_));
 sky130_fd_sc_hd__a22o_1 _16691_ (.A1(\cpuregs[16][15] ),
    .A2(_13032_),
    .B1(_12973_),
    .B2(_13034_),
    .X(_03326_));
 sky130_fd_sc_hd__a22o_1 _16692_ (.A1(\cpuregs[16][14] ),
    .A2(_13032_),
    .B1(_12976_),
    .B2(_13034_),
    .X(_03325_));
 sky130_fd_sc_hd__a22o_1 _16693_ (.A1(\cpuregs[16][13] ),
    .A2(_13032_),
    .B1(_12977_),
    .B2(_13034_),
    .X(_03324_));
 sky130_fd_sc_hd__a22o_1 _16694_ (.A1(\cpuregs[16][12] ),
    .A2(_13032_),
    .B1(_12978_),
    .B2(_13034_),
    .X(_03323_));
 sky130_fd_sc_hd__buf_1 _16695_ (.A(_13031_),
    .X(_13035_));
 sky130_fd_sc_hd__buf_1 _16696_ (.A(_13033_),
    .X(_13036_));
 sky130_fd_sc_hd__a22o_1 _16697_ (.A1(\cpuregs[16][11] ),
    .A2(_13035_),
    .B1(_12980_),
    .B2(_13036_),
    .X(_03322_));
 sky130_fd_sc_hd__a22o_1 _16698_ (.A1(\cpuregs[16][10] ),
    .A2(_13035_),
    .B1(_12982_),
    .B2(_13036_),
    .X(_03321_));
 sky130_fd_sc_hd__a22o_1 _16699_ (.A1(\cpuregs[16][9] ),
    .A2(_13035_),
    .B1(_12983_),
    .B2(_13036_),
    .X(_03320_));
 sky130_fd_sc_hd__a22o_1 _16700_ (.A1(\cpuregs[16][8] ),
    .A2(_13035_),
    .B1(_12984_),
    .B2(_13036_),
    .X(_03319_));
 sky130_fd_sc_hd__buf_1 _16701_ (.A(_13031_),
    .X(_13037_));
 sky130_fd_sc_hd__buf_1 _16702_ (.A(_13033_),
    .X(_13038_));
 sky130_fd_sc_hd__a22o_1 _16703_ (.A1(\cpuregs[16][7] ),
    .A2(_13037_),
    .B1(_12986_),
    .B2(_13038_),
    .X(_03318_));
 sky130_fd_sc_hd__a22o_1 _16704_ (.A1(\cpuregs[16][6] ),
    .A2(_13037_),
    .B1(_12988_),
    .B2(_13038_),
    .X(_03317_));
 sky130_fd_sc_hd__a22o_1 _16705_ (.A1(\cpuregs[16][5] ),
    .A2(_13037_),
    .B1(_12989_),
    .B2(_13038_),
    .X(_03316_));
 sky130_fd_sc_hd__a22o_1 _16706_ (.A1(\cpuregs[16][4] ),
    .A2(_13037_),
    .B1(_12990_),
    .B2(_13038_),
    .X(_03315_));
 sky130_fd_sc_hd__buf_1 _16707_ (.A(_13031_),
    .X(_13039_));
 sky130_fd_sc_hd__buf_1 _16708_ (.A(_13033_),
    .X(_13040_));
 sky130_fd_sc_hd__a22o_1 _16709_ (.A1(\cpuregs[16][3] ),
    .A2(_13039_),
    .B1(_12992_),
    .B2(_13040_),
    .X(_03314_));
 sky130_fd_sc_hd__a22o_1 _16710_ (.A1(\cpuregs[16][2] ),
    .A2(_13039_),
    .B1(_12994_),
    .B2(_13040_),
    .X(_03313_));
 sky130_fd_sc_hd__a22o_1 _16711_ (.A1(\cpuregs[16][1] ),
    .A2(_13039_),
    .B1(_12995_),
    .B2(_13040_),
    .X(_03312_));
 sky130_fd_sc_hd__a22o_1 _16712_ (.A1(\cpuregs[16][0] ),
    .A2(_13039_),
    .B1(_12996_),
    .B2(_13040_),
    .X(_03311_));
 sky130_fd_sc_hd__or4_4 _16713_ (.A(_12769_),
    .B(_12770_),
    .C(_12771_),
    .D(_12657_),
    .X(_13041_));
 sky130_fd_sc_hd__clkbuf_4 _16714_ (.A(_13041_),
    .X(_13042_));
 sky130_fd_sc_hd__buf_1 _16715_ (.A(_13042_),
    .X(_13043_));
 sky130_vsdinv _16716_ (.A(_13041_),
    .Y(_13044_));
 sky130_fd_sc_hd__clkbuf_4 _16717_ (.A(_13044_),
    .X(_13045_));
 sky130_fd_sc_hd__buf_1 _16718_ (.A(_13045_),
    .X(_13046_));
 sky130_fd_sc_hd__a22o_1 _16719_ (.A1(\cpuregs[17][31] ),
    .A2(_13043_),
    .B1(_12946_),
    .B2(_13046_),
    .X(_03310_));
 sky130_fd_sc_hd__a22o_1 _16720_ (.A1(\cpuregs[17][30] ),
    .A2(_13043_),
    .B1(_12950_),
    .B2(_13046_),
    .X(_03309_));
 sky130_fd_sc_hd__a22o_1 _16721_ (.A1(\cpuregs[17][29] ),
    .A2(_13043_),
    .B1(_12951_),
    .B2(_13046_),
    .X(_03308_));
 sky130_fd_sc_hd__a22o_1 _16722_ (.A1(\cpuregs[17][28] ),
    .A2(_13043_),
    .B1(_12952_),
    .B2(_13046_),
    .X(_03307_));
 sky130_fd_sc_hd__buf_1 _16723_ (.A(_13042_),
    .X(_13047_));
 sky130_fd_sc_hd__buf_1 _16724_ (.A(_13045_),
    .X(_13048_));
 sky130_fd_sc_hd__a22o_1 _16725_ (.A1(\cpuregs[17][27] ),
    .A2(_13047_),
    .B1(_12954_),
    .B2(_13048_),
    .X(_03306_));
 sky130_fd_sc_hd__a22o_1 _16726_ (.A1(\cpuregs[17][26] ),
    .A2(_13047_),
    .B1(_12956_),
    .B2(_13048_),
    .X(_03305_));
 sky130_fd_sc_hd__a22o_1 _16727_ (.A1(\cpuregs[17][25] ),
    .A2(_13047_),
    .B1(_12957_),
    .B2(_13048_),
    .X(_03304_));
 sky130_fd_sc_hd__a22o_1 _16728_ (.A1(\cpuregs[17][24] ),
    .A2(_13047_),
    .B1(_12958_),
    .B2(_13048_),
    .X(_03303_));
 sky130_fd_sc_hd__buf_1 _16729_ (.A(_13042_),
    .X(_13049_));
 sky130_fd_sc_hd__buf_1 _16730_ (.A(_13045_),
    .X(_13050_));
 sky130_fd_sc_hd__a22o_1 _16731_ (.A1(\cpuregs[17][23] ),
    .A2(_13049_),
    .B1(_12960_),
    .B2(_13050_),
    .X(_03302_));
 sky130_fd_sc_hd__a22o_1 _16732_ (.A1(\cpuregs[17][22] ),
    .A2(_13049_),
    .B1(_12962_),
    .B2(_13050_),
    .X(_03301_));
 sky130_fd_sc_hd__a22o_1 _16733_ (.A1(\cpuregs[17][21] ),
    .A2(_13049_),
    .B1(_12963_),
    .B2(_13050_),
    .X(_03300_));
 sky130_fd_sc_hd__a22o_1 _16734_ (.A1(\cpuregs[17][20] ),
    .A2(_13049_),
    .B1(_12964_),
    .B2(_13050_),
    .X(_03299_));
 sky130_fd_sc_hd__buf_1 _16735_ (.A(_13042_),
    .X(_13051_));
 sky130_fd_sc_hd__buf_1 _16736_ (.A(_13045_),
    .X(_13052_));
 sky130_fd_sc_hd__a22o_1 _16737_ (.A1(\cpuregs[17][19] ),
    .A2(_13051_),
    .B1(_12966_),
    .B2(_13052_),
    .X(_03298_));
 sky130_fd_sc_hd__a22o_1 _16738_ (.A1(\cpuregs[17][18] ),
    .A2(_13051_),
    .B1(_12968_),
    .B2(_13052_),
    .X(_03297_));
 sky130_fd_sc_hd__a22o_1 _16739_ (.A1(\cpuregs[17][17] ),
    .A2(_13051_),
    .B1(_12969_),
    .B2(_13052_),
    .X(_03296_));
 sky130_fd_sc_hd__a22o_1 _16740_ (.A1(\cpuregs[17][16] ),
    .A2(_13051_),
    .B1(_12970_),
    .B2(_13052_),
    .X(_03295_));
 sky130_fd_sc_hd__buf_2 _16741_ (.A(_13041_),
    .X(_13053_));
 sky130_fd_sc_hd__buf_1 _16742_ (.A(_13053_),
    .X(_13054_));
 sky130_fd_sc_hd__clkbuf_4 _16743_ (.A(_13044_),
    .X(_13055_));
 sky130_fd_sc_hd__buf_1 _16744_ (.A(_13055_),
    .X(_13056_));
 sky130_fd_sc_hd__a22o_1 _16745_ (.A1(\cpuregs[17][15] ),
    .A2(_13054_),
    .B1(_12973_),
    .B2(_13056_),
    .X(_03294_));
 sky130_fd_sc_hd__a22o_1 _16746_ (.A1(\cpuregs[17][14] ),
    .A2(_13054_),
    .B1(_12976_),
    .B2(_13056_),
    .X(_03293_));
 sky130_fd_sc_hd__a22o_1 _16747_ (.A1(\cpuregs[17][13] ),
    .A2(_13054_),
    .B1(_12977_),
    .B2(_13056_),
    .X(_03292_));
 sky130_fd_sc_hd__a22o_1 _16748_ (.A1(\cpuregs[17][12] ),
    .A2(_13054_),
    .B1(_12978_),
    .B2(_13056_),
    .X(_03291_));
 sky130_fd_sc_hd__buf_1 _16749_ (.A(_13053_),
    .X(_13057_));
 sky130_fd_sc_hd__buf_1 _16750_ (.A(_13055_),
    .X(_13058_));
 sky130_fd_sc_hd__a22o_1 _16751_ (.A1(\cpuregs[17][11] ),
    .A2(_13057_),
    .B1(_12980_),
    .B2(_13058_),
    .X(_03290_));
 sky130_fd_sc_hd__a22o_1 _16752_ (.A1(\cpuregs[17][10] ),
    .A2(_13057_),
    .B1(_12982_),
    .B2(_13058_),
    .X(_03289_));
 sky130_fd_sc_hd__a22o_1 _16753_ (.A1(\cpuregs[17][9] ),
    .A2(_13057_),
    .B1(_12983_),
    .B2(_13058_),
    .X(_03288_));
 sky130_fd_sc_hd__a22o_1 _16754_ (.A1(\cpuregs[17][8] ),
    .A2(_13057_),
    .B1(_12984_),
    .B2(_13058_),
    .X(_03287_));
 sky130_fd_sc_hd__buf_1 _16755_ (.A(_13053_),
    .X(_13059_));
 sky130_fd_sc_hd__buf_1 _16756_ (.A(_13055_),
    .X(_13060_));
 sky130_fd_sc_hd__a22o_1 _16757_ (.A1(\cpuregs[17][7] ),
    .A2(_13059_),
    .B1(_12986_),
    .B2(_13060_),
    .X(_03286_));
 sky130_fd_sc_hd__a22o_1 _16758_ (.A1(\cpuregs[17][6] ),
    .A2(_13059_),
    .B1(_12988_),
    .B2(_13060_),
    .X(_03285_));
 sky130_fd_sc_hd__a22o_1 _16759_ (.A1(\cpuregs[17][5] ),
    .A2(_13059_),
    .B1(_12989_),
    .B2(_13060_),
    .X(_03284_));
 sky130_fd_sc_hd__a22o_1 _16760_ (.A1(\cpuregs[17][4] ),
    .A2(_13059_),
    .B1(_12990_),
    .B2(_13060_),
    .X(_03283_));
 sky130_fd_sc_hd__buf_1 _16761_ (.A(_13053_),
    .X(_13061_));
 sky130_fd_sc_hd__buf_1 _16762_ (.A(_13055_),
    .X(_13062_));
 sky130_fd_sc_hd__a22o_1 _16763_ (.A1(\cpuregs[17][3] ),
    .A2(_13061_),
    .B1(_12992_),
    .B2(_13062_),
    .X(_03282_));
 sky130_fd_sc_hd__a22o_1 _16764_ (.A1(\cpuregs[17][2] ),
    .A2(_13061_),
    .B1(_12994_),
    .B2(_13062_),
    .X(_03281_));
 sky130_fd_sc_hd__a22o_1 _16765_ (.A1(\cpuregs[17][1] ),
    .A2(_13061_),
    .B1(_12995_),
    .B2(_13062_),
    .X(_03280_));
 sky130_fd_sc_hd__a22o_1 _16766_ (.A1(\cpuregs[17][0] ),
    .A2(_13061_),
    .B1(_12996_),
    .B2(_13062_),
    .X(_03279_));
 sky130_fd_sc_hd__clkbuf_4 _16767_ (.A(_11709_),
    .X(_13063_));
 sky130_fd_sc_hd__clkbuf_2 _16768_ (.A(\pcpi_mul.rs2[31] ),
    .X(_13064_));
 sky130_fd_sc_hd__clkbuf_2 _16769_ (.A(_13064_),
    .X(_13065_));
 sky130_fd_sc_hd__buf_1 _16770_ (.A(_13065_),
    .X(_13066_));
 sky130_fd_sc_hd__buf_1 _16771_ (.A(_13066_),
    .X(_13067_));
 sky130_fd_sc_hd__buf_1 _16772_ (.A(_13067_),
    .X(_13068_));
 sky130_fd_sc_hd__buf_1 _16773_ (.A(_11694_),
    .X(_13069_));
 sky130_fd_sc_hd__clkbuf_2 _16774_ (.A(_13069_),
    .X(_13070_));
 sky130_fd_sc_hd__a22o_1 _16775_ (.A1(_11712_),
    .A2(_13063_),
    .B1(_13068_),
    .B2(_13070_),
    .X(_03278_));
 sky130_fd_sc_hd__clkbuf_2 _16776_ (.A(\pcpi_mul.rs2[30] ),
    .X(_13071_));
 sky130_fd_sc_hd__a22o_1 _16777_ (.A1(_13071_),
    .A2(_13070_),
    .B1(_12686_),
    .B2(_03728_),
    .X(_03277_));
 sky130_fd_sc_hd__buf_1 _16778_ (.A(\pcpi_mul.rs2[29] ),
    .X(_13072_));
 sky130_fd_sc_hd__buf_1 _16779_ (.A(_13072_),
    .X(_13073_));
 sky130_fd_sc_hd__buf_2 _16780_ (.A(_13073_),
    .X(_13074_));
 sky130_fd_sc_hd__buf_1 _16781_ (.A(_13074_),
    .X(_13075_));
 sky130_fd_sc_hd__buf_1 _16782_ (.A(_13075_),
    .X(_13076_));
 sky130_fd_sc_hd__clkbuf_2 _16783_ (.A(_13076_),
    .X(_13077_));
 sky130_fd_sc_hd__a22o_1 _16784_ (.A1(_13077_),
    .A2(_13070_),
    .B1(_12687_),
    .B2(_03728_),
    .X(_03276_));
 sky130_fd_sc_hd__buf_1 _16785_ (.A(\pcpi_mul.rs2[28] ),
    .X(_13078_));
 sky130_fd_sc_hd__clkbuf_2 _16786_ (.A(_13078_),
    .X(_13079_));
 sky130_fd_sc_hd__clkbuf_2 _16787_ (.A(_13079_),
    .X(_13080_));
 sky130_fd_sc_hd__buf_1 _16788_ (.A(_13080_),
    .X(_13081_));
 sky130_fd_sc_hd__buf_1 _16789_ (.A(_13081_),
    .X(_13082_));
 sky130_fd_sc_hd__buf_1 _16790_ (.A(_13082_),
    .X(_13083_));
 sky130_fd_sc_hd__buf_1 _16791_ (.A(_13069_),
    .X(_13084_));
 sky130_fd_sc_hd__a22o_1 _16792_ (.A1(_13083_),
    .A2(_13084_),
    .B1(_12688_),
    .B2(_03728_),
    .X(_03275_));
 sky130_fd_sc_hd__buf_1 _16793_ (.A(_11708_),
    .X(_13085_));
 sky130_fd_sc_hd__buf_1 _16794_ (.A(_13085_),
    .X(_13086_));
 sky130_fd_sc_hd__a22o_1 _16795_ (.A1(\pcpi_mul.rs2[27] ),
    .A2(_13084_),
    .B1(_12691_),
    .B2(_13086_),
    .X(_03274_));
 sky130_fd_sc_hd__buf_1 _16796_ (.A(\pcpi_mul.rs2[26] ),
    .X(_13087_));
 sky130_fd_sc_hd__buf_2 _16797_ (.A(_13087_),
    .X(_13088_));
 sky130_fd_sc_hd__buf_1 _16798_ (.A(_13088_),
    .X(_13089_));
 sky130_fd_sc_hd__buf_2 _16799_ (.A(_13089_),
    .X(_13090_));
 sky130_fd_sc_hd__a22o_1 _16800_ (.A1(_13090_),
    .A2(_13084_),
    .B1(_12693_),
    .B2(_13086_),
    .X(_03273_));
 sky130_fd_sc_hd__clkbuf_2 _16801_ (.A(\pcpi_mul.rs2[25] ),
    .X(_13091_));
 sky130_fd_sc_hd__buf_2 _16802_ (.A(_13091_),
    .X(_13092_));
 sky130_fd_sc_hd__buf_1 _16803_ (.A(_13092_),
    .X(_13093_));
 sky130_fd_sc_hd__clkbuf_2 _16804_ (.A(_13093_),
    .X(_13094_));
 sky130_fd_sc_hd__a22o_1 _16805_ (.A1(_13094_),
    .A2(_13084_),
    .B1(_12694_),
    .B2(_13086_),
    .X(_03272_));
 sky130_fd_sc_hd__buf_1 _16806_ (.A(_13069_),
    .X(_13095_));
 sky130_fd_sc_hd__a22o_1 _16807_ (.A1(\pcpi_mul.rs2[24] ),
    .A2(_13095_),
    .B1(_12695_),
    .B2(_13086_),
    .X(_03271_));
 sky130_fd_sc_hd__clkbuf_2 _16808_ (.A(\pcpi_mul.rs2[23] ),
    .X(_13096_));
 sky130_fd_sc_hd__buf_1 _16809_ (.A(_13096_),
    .X(_13097_));
 sky130_fd_sc_hd__buf_2 _16810_ (.A(_13097_),
    .X(_13098_));
 sky130_fd_sc_hd__buf_2 _16811_ (.A(_13098_),
    .X(_13099_));
 sky130_fd_sc_hd__buf_1 _16812_ (.A(_13085_),
    .X(_13100_));
 sky130_fd_sc_hd__a22o_1 _16813_ (.A1(_13099_),
    .A2(_13095_),
    .B1(_12697_),
    .B2(_13100_),
    .X(_03270_));
 sky130_fd_sc_hd__clkbuf_2 _16814_ (.A(\pcpi_mul.rs2[22] ),
    .X(_13101_));
 sky130_fd_sc_hd__buf_1 _16815_ (.A(_13101_),
    .X(_13102_));
 sky130_fd_sc_hd__buf_2 _16816_ (.A(_13102_),
    .X(_13103_));
 sky130_fd_sc_hd__clkbuf_2 _16817_ (.A(_13103_),
    .X(_13104_));
 sky130_fd_sc_hd__a22o_1 _16818_ (.A1(_13104_),
    .A2(_13095_),
    .B1(_12699_),
    .B2(_13100_),
    .X(_03269_));
 sky130_fd_sc_hd__a22o_1 _16819_ (.A1(\pcpi_mul.rs2[21] ),
    .A2(_13095_),
    .B1(_12700_),
    .B2(_13100_),
    .X(_03268_));
 sky130_fd_sc_hd__buf_2 _16820_ (.A(\pcpi_mul.rs2[20] ),
    .X(_13105_));
 sky130_fd_sc_hd__clkbuf_2 _16821_ (.A(_13105_),
    .X(_13106_));
 sky130_fd_sc_hd__buf_1 _16822_ (.A(_13106_),
    .X(_13107_));
 sky130_fd_sc_hd__buf_2 _16823_ (.A(_13107_),
    .X(_13108_));
 sky130_fd_sc_hd__clkbuf_2 _16824_ (.A(_13069_),
    .X(_13109_));
 sky130_fd_sc_hd__a22o_1 _16825_ (.A1(_13108_),
    .A2(_13109_),
    .B1(_12701_),
    .B2(_13100_),
    .X(_03267_));
 sky130_fd_sc_hd__buf_1 _16826_ (.A(\pcpi_mul.rs2[19] ),
    .X(_13110_));
 sky130_fd_sc_hd__clkbuf_2 _16827_ (.A(_13110_),
    .X(_13111_));
 sky130_fd_sc_hd__buf_2 _16828_ (.A(_13111_),
    .X(_13112_));
 sky130_fd_sc_hd__buf_1 _16829_ (.A(_13112_),
    .X(_13113_));
 sky130_fd_sc_hd__buf_2 _16830_ (.A(_13113_),
    .X(_13114_));
 sky130_fd_sc_hd__buf_1 _16831_ (.A(_13085_),
    .X(_13115_));
 sky130_fd_sc_hd__a22o_1 _16832_ (.A1(_13114_),
    .A2(_13109_),
    .B1(_12703_),
    .B2(_13115_),
    .X(_03266_));
 sky130_fd_sc_hd__a22o_1 _16833_ (.A1(\pcpi_mul.rs2[18] ),
    .A2(_13109_),
    .B1(_12705_),
    .B2(_13115_),
    .X(_03265_));
 sky130_fd_sc_hd__clkbuf_2 _16834_ (.A(\pcpi_mul.rs2[17] ),
    .X(_13116_));
 sky130_fd_sc_hd__clkbuf_2 _16835_ (.A(_13116_),
    .X(_13117_));
 sky130_fd_sc_hd__buf_2 _16836_ (.A(_13117_),
    .X(_13118_));
 sky130_fd_sc_hd__buf_2 _16837_ (.A(_13118_),
    .X(_13119_));
 sky130_fd_sc_hd__a22o_1 _16838_ (.A1(_13119_),
    .A2(_13109_),
    .B1(_12706_),
    .B2(_13115_),
    .X(_03264_));
 sky130_fd_sc_hd__clkbuf_2 _16839_ (.A(\pcpi_mul.rs2[16] ),
    .X(_13120_));
 sky130_fd_sc_hd__clkbuf_2 _16840_ (.A(_13120_),
    .X(_13121_));
 sky130_fd_sc_hd__buf_2 _16841_ (.A(_13121_),
    .X(_13122_));
 sky130_fd_sc_hd__buf_2 _16842_ (.A(_13122_),
    .X(_13123_));
 sky130_fd_sc_hd__clkbuf_2 _16843_ (.A(_11694_),
    .X(_13124_));
 sky130_fd_sc_hd__buf_1 _16844_ (.A(_13124_),
    .X(_13125_));
 sky130_fd_sc_hd__a22o_1 _16845_ (.A1(_13123_),
    .A2(_13125_),
    .B1(_12707_),
    .B2(_13115_),
    .X(_03263_));
 sky130_fd_sc_hd__clkbuf_4 _16846_ (.A(\pcpi_mul.rs2[15] ),
    .X(_13126_));
 sky130_fd_sc_hd__buf_1 _16847_ (.A(_13085_),
    .X(_13127_));
 sky130_fd_sc_hd__a22o_1 _16848_ (.A1(_13126_),
    .A2(_13125_),
    .B1(_12711_),
    .B2(_13127_),
    .X(_03262_));
 sky130_fd_sc_hd__buf_1 _16849_ (.A(\pcpi_mul.rs2[14] ),
    .X(_13128_));
 sky130_fd_sc_hd__clkbuf_2 _16850_ (.A(_13128_),
    .X(_13129_));
 sky130_fd_sc_hd__clkbuf_2 _16851_ (.A(_13129_),
    .X(_13130_));
 sky130_fd_sc_hd__a22o_1 _16852_ (.A1(_13130_),
    .A2(_13125_),
    .B1(_12714_),
    .B2(_13127_),
    .X(_03261_));
 sky130_fd_sc_hd__buf_1 _16853_ (.A(\pcpi_mul.rs2[13] ),
    .X(_13131_));
 sky130_fd_sc_hd__clkbuf_2 _16854_ (.A(_13131_),
    .X(_13132_));
 sky130_fd_sc_hd__clkbuf_2 _16855_ (.A(_13132_),
    .X(_13133_));
 sky130_fd_sc_hd__a22o_1 _16856_ (.A1(_13133_),
    .A2(_13125_),
    .B1(_12716_),
    .B2(_13127_),
    .X(_03260_));
 sky130_fd_sc_hd__buf_1 _16857_ (.A(_13124_),
    .X(_13134_));
 sky130_fd_sc_hd__a22o_1 _16858_ (.A1(\pcpi_mul.rs2[12] ),
    .A2(_13134_),
    .B1(_12717_),
    .B2(_13127_),
    .X(_03259_));
 sky130_fd_sc_hd__clkbuf_4 _16859_ (.A(\pcpi_mul.rs2[11] ),
    .X(_13135_));
 sky130_fd_sc_hd__clkbuf_2 _16860_ (.A(_13135_),
    .X(_13136_));
 sky130_fd_sc_hd__clkbuf_2 _16861_ (.A(_13136_),
    .X(_13137_));
 sky130_fd_sc_hd__buf_2 _16862_ (.A(_13137_),
    .X(_13138_));
 sky130_fd_sc_hd__clkbuf_2 _16863_ (.A(_11708_),
    .X(_13139_));
 sky130_fd_sc_hd__buf_1 _16864_ (.A(_13139_),
    .X(_13140_));
 sky130_fd_sc_hd__a22o_1 _16865_ (.A1(_13138_),
    .A2(_13134_),
    .B1(_12720_),
    .B2(_13140_),
    .X(_03258_));
 sky130_fd_sc_hd__clkbuf_2 _16866_ (.A(\pcpi_mul.rs2[10] ),
    .X(_13141_));
 sky130_fd_sc_hd__clkbuf_2 _16867_ (.A(_13141_),
    .X(_13142_));
 sky130_fd_sc_hd__clkbuf_2 _16868_ (.A(_13142_),
    .X(_13143_));
 sky130_fd_sc_hd__clkbuf_2 _16869_ (.A(_13143_),
    .X(_13144_));
 sky130_fd_sc_hd__a22o_1 _16870_ (.A1(_13144_),
    .A2(_13134_),
    .B1(_12722_),
    .B2(_13140_),
    .X(_03257_));
 sky130_fd_sc_hd__a22o_1 _16871_ (.A1(\pcpi_mul.rs2[9] ),
    .A2(_13134_),
    .B1(_12724_),
    .B2(_13140_),
    .X(_03256_));
 sky130_fd_sc_hd__buf_1 _16872_ (.A(\pcpi_mul.rs2[8] ),
    .X(_13145_));
 sky130_fd_sc_hd__clkbuf_4 _16873_ (.A(_13145_),
    .X(_13146_));
 sky130_fd_sc_hd__buf_1 _16874_ (.A(_13146_),
    .X(_13147_));
 sky130_fd_sc_hd__buf_2 _16875_ (.A(_13147_),
    .X(_13148_));
 sky130_fd_sc_hd__buf_2 _16876_ (.A(_13148_),
    .X(_13149_));
 sky130_fd_sc_hd__buf_1 _16877_ (.A(_13124_),
    .X(_13150_));
 sky130_fd_sc_hd__a22o_1 _16878_ (.A1(_13149_),
    .A2(_13150_),
    .B1(_12725_),
    .B2(_13140_),
    .X(_03255_));
 sky130_fd_sc_hd__buf_1 _16879_ (.A(\pcpi_mul.rs2[7] ),
    .X(_13151_));
 sky130_fd_sc_hd__clkbuf_2 _16880_ (.A(_13151_),
    .X(_13152_));
 sky130_fd_sc_hd__buf_1 _16881_ (.A(_13152_),
    .X(_13153_));
 sky130_fd_sc_hd__buf_2 _16882_ (.A(_13153_),
    .X(_13154_));
 sky130_fd_sc_hd__buf_2 _16883_ (.A(_13154_),
    .X(_13155_));
 sky130_fd_sc_hd__buf_1 _16884_ (.A(_13139_),
    .X(_13156_));
 sky130_fd_sc_hd__a22o_1 _16885_ (.A1(_13155_),
    .A2(_13150_),
    .B1(_12728_),
    .B2(_13156_),
    .X(_03254_));
 sky130_fd_sc_hd__a22o_1 _16886_ (.A1(\pcpi_mul.rs2[6] ),
    .A2(_13150_),
    .B1(_12731_),
    .B2(_13156_),
    .X(_03253_));
 sky130_fd_sc_hd__buf_1 _16887_ (.A(\pcpi_mul.rs2[5] ),
    .X(_13157_));
 sky130_fd_sc_hd__buf_1 _16888_ (.A(_13157_),
    .X(_13158_));
 sky130_fd_sc_hd__clkbuf_2 _16889_ (.A(_13158_),
    .X(_13159_));
 sky130_fd_sc_hd__buf_1 _16890_ (.A(_13159_),
    .X(_13160_));
 sky130_fd_sc_hd__clkbuf_2 _16891_ (.A(_13160_),
    .X(_13161_));
 sky130_fd_sc_hd__buf_2 _16892_ (.A(_13161_),
    .X(_13162_));
 sky130_fd_sc_hd__a22o_1 _16893_ (.A1(_13162_),
    .A2(_13150_),
    .B1(_12733_),
    .B2(_13156_),
    .X(_03252_));
 sky130_fd_sc_hd__buf_1 _16894_ (.A(\pcpi_mul.rs2[4] ),
    .X(_13163_));
 sky130_fd_sc_hd__buf_1 _16895_ (.A(_13163_),
    .X(_13164_));
 sky130_fd_sc_hd__clkbuf_2 _16896_ (.A(_13164_),
    .X(_13165_));
 sky130_fd_sc_hd__buf_1 _16897_ (.A(_13165_),
    .X(_13166_));
 sky130_fd_sc_hd__clkbuf_2 _16898_ (.A(_13166_),
    .X(_13167_));
 sky130_fd_sc_hd__buf_2 _16899_ (.A(_13167_),
    .X(_13168_));
 sky130_fd_sc_hd__buf_1 _16900_ (.A(_13124_),
    .X(_13169_));
 sky130_fd_sc_hd__a22o_1 _16901_ (.A1(_13168_),
    .A2(_13169_),
    .B1(_12735_),
    .B2(_13156_),
    .X(_03251_));
 sky130_fd_sc_hd__buf_1 _16902_ (.A(_13139_),
    .X(_13170_));
 sky130_fd_sc_hd__a22o_1 _16903_ (.A1(\pcpi_mul.rs2[3] ),
    .A2(_13169_),
    .B1(_12738_),
    .B2(_13170_),
    .X(_03250_));
 sky130_fd_sc_hd__buf_1 _16904_ (.A(\pcpi_mul.rs2[2] ),
    .X(_13171_));
 sky130_fd_sc_hd__buf_1 _16905_ (.A(_13171_),
    .X(_13172_));
 sky130_fd_sc_hd__clkbuf_2 _16906_ (.A(_13172_),
    .X(_13173_));
 sky130_fd_sc_hd__clkbuf_2 _16907_ (.A(_13173_),
    .X(_13174_));
 sky130_fd_sc_hd__buf_2 _16908_ (.A(_13174_),
    .X(_13175_));
 sky130_fd_sc_hd__a22o_1 _16909_ (.A1(_13175_),
    .A2(_13169_),
    .B1(_12741_),
    .B2(_13170_),
    .X(_03249_));
 sky130_fd_sc_hd__buf_1 _16910_ (.A(\pcpi_mul.rs2[1] ),
    .X(_13176_));
 sky130_fd_sc_hd__buf_1 _16911_ (.A(_13176_),
    .X(_13177_));
 sky130_fd_sc_hd__clkbuf_2 _16912_ (.A(_13177_),
    .X(_13178_));
 sky130_fd_sc_hd__clkbuf_2 _16913_ (.A(_13178_),
    .X(_13179_));
 sky130_fd_sc_hd__buf_2 _16914_ (.A(_13179_),
    .X(_13180_));
 sky130_fd_sc_hd__a22o_1 _16915_ (.A1(_13180_),
    .A2(_13169_),
    .B1(_12743_),
    .B2(_13170_),
    .X(_03248_));
 sky130_fd_sc_hd__clkbuf_2 _16916_ (.A(_11693_),
    .X(_13181_));
 sky130_fd_sc_hd__clkbuf_2 _16917_ (.A(_13181_),
    .X(_13182_));
 sky130_fd_sc_hd__a22o_1 _16918_ (.A1(\pcpi_mul.rs2[0] ),
    .A2(_13182_),
    .B1(_12745_),
    .B2(_13170_),
    .X(_03247_));
 sky130_fd_sc_hd__buf_1 _16919_ (.A(_11583_),
    .X(_13183_));
 sky130_fd_sc_hd__buf_1 _16920_ (.A(_11584_),
    .X(_13184_));
 sky130_fd_sc_hd__a22o_1 _16921_ (.A1(net273),
    .A2(_13183_),
    .B1(_02541_),
    .B2(_13184_),
    .X(_03246_));
 sky130_fd_sc_hd__a22o_1 _16922_ (.A1(net272),
    .A2(_13183_),
    .B1(_02540_),
    .B2(_13184_),
    .X(_03245_));
 sky130_fd_sc_hd__a22o_1 _16923_ (.A1(net271),
    .A2(_13183_),
    .B1(_02539_),
    .B2(_13184_),
    .X(_03244_));
 sky130_fd_sc_hd__a22o_1 _16924_ (.A1(net270),
    .A2(_11583_),
    .B1(_02538_),
    .B2(_11584_),
    .X(_03243_));
 sky130_vsdinv _16925_ (.A(_00328_),
    .Y(_13185_));
 sky130_fd_sc_hd__or4_4 _16926_ (.A(_00327_),
    .B(_11607_),
    .C(_00330_),
    .D(_11598_),
    .X(_13186_));
 sky130_fd_sc_hd__o32a_1 _16927_ (.A1(_11888_),
    .A2(_13185_),
    .A3(_13186_),
    .B1(_11918_),
    .B2(_11614_),
    .X(_13187_));
 sky130_vsdinv _16928_ (.A(_13187_),
    .Y(_03242_));
 sky130_fd_sc_hd__buf_1 _16929_ (.A(_11600_),
    .X(_13188_));
 sky130_fd_sc_hd__o32a_1 _16930_ (.A1(_11887_),
    .A2(_13185_),
    .A3(_13186_),
    .B1(_11961_),
    .B2(_13188_),
    .X(_13189_));
 sky130_vsdinv _16931_ (.A(_13189_),
    .Y(_03241_));
 sky130_fd_sc_hd__or2_1 _16932_ (.A(_12658_),
    .B(_12876_),
    .X(_13190_));
 sky130_fd_sc_hd__clkbuf_4 _16933_ (.A(_13190_),
    .X(_13191_));
 sky130_fd_sc_hd__buf_1 _16934_ (.A(_13191_),
    .X(_13192_));
 sky130_fd_sc_hd__clkbuf_2 _16935_ (.A(\cpuregs_wrdata[31] ),
    .X(_13193_));
 sky130_vsdinv _16936_ (.A(_13190_),
    .Y(_13194_));
 sky130_fd_sc_hd__buf_4 _16937_ (.A(_13194_),
    .X(_13195_));
 sky130_fd_sc_hd__buf_1 _16938_ (.A(_13195_),
    .X(_13196_));
 sky130_fd_sc_hd__a22o_1 _16939_ (.A1(\cpuregs[13][31] ),
    .A2(_13192_),
    .B1(_13193_),
    .B2(_13196_),
    .X(_03240_));
 sky130_fd_sc_hd__clkbuf_2 _16940_ (.A(\cpuregs_wrdata[30] ),
    .X(_13197_));
 sky130_fd_sc_hd__a22o_1 _16941_ (.A1(\cpuregs[13][30] ),
    .A2(_13192_),
    .B1(_13197_),
    .B2(_13196_),
    .X(_03239_));
 sky130_fd_sc_hd__clkbuf_2 _16942_ (.A(\cpuregs_wrdata[29] ),
    .X(_13198_));
 sky130_fd_sc_hd__a22o_1 _16943_ (.A1(\cpuregs[13][29] ),
    .A2(_13192_),
    .B1(_13198_),
    .B2(_13196_),
    .X(_03238_));
 sky130_fd_sc_hd__clkbuf_2 _16944_ (.A(\cpuregs_wrdata[28] ),
    .X(_13199_));
 sky130_fd_sc_hd__a22o_1 _16945_ (.A1(\cpuregs[13][28] ),
    .A2(_13192_),
    .B1(_13199_),
    .B2(_13196_),
    .X(_03237_));
 sky130_fd_sc_hd__buf_1 _16946_ (.A(_13191_),
    .X(_13200_));
 sky130_fd_sc_hd__clkbuf_2 _16947_ (.A(\cpuregs_wrdata[27] ),
    .X(_13201_));
 sky130_fd_sc_hd__buf_1 _16948_ (.A(_13195_),
    .X(_13202_));
 sky130_fd_sc_hd__a22o_1 _16949_ (.A1(\cpuregs[13][27] ),
    .A2(_13200_),
    .B1(_13201_),
    .B2(_13202_),
    .X(_03236_));
 sky130_fd_sc_hd__clkbuf_2 _16950_ (.A(\cpuregs_wrdata[26] ),
    .X(_13203_));
 sky130_fd_sc_hd__a22o_1 _16951_ (.A1(\cpuregs[13][26] ),
    .A2(_13200_),
    .B1(_13203_),
    .B2(_13202_),
    .X(_03235_));
 sky130_fd_sc_hd__clkbuf_2 _16952_ (.A(\cpuregs_wrdata[25] ),
    .X(_13204_));
 sky130_fd_sc_hd__a22o_1 _16953_ (.A1(\cpuregs[13][25] ),
    .A2(_13200_),
    .B1(_13204_),
    .B2(_13202_),
    .X(_03234_));
 sky130_fd_sc_hd__clkbuf_2 _16954_ (.A(\cpuregs_wrdata[24] ),
    .X(_13205_));
 sky130_fd_sc_hd__a22o_1 _16955_ (.A1(\cpuregs[13][24] ),
    .A2(_13200_),
    .B1(_13205_),
    .B2(_13202_),
    .X(_03233_));
 sky130_fd_sc_hd__buf_1 _16956_ (.A(_13191_),
    .X(_13206_));
 sky130_fd_sc_hd__clkbuf_2 _16957_ (.A(\cpuregs_wrdata[23] ),
    .X(_13207_));
 sky130_fd_sc_hd__buf_1 _16958_ (.A(_13195_),
    .X(_13208_));
 sky130_fd_sc_hd__a22o_1 _16959_ (.A1(\cpuregs[13][23] ),
    .A2(_13206_),
    .B1(_13207_),
    .B2(_13208_),
    .X(_03232_));
 sky130_fd_sc_hd__clkbuf_2 _16960_ (.A(\cpuregs_wrdata[22] ),
    .X(_13209_));
 sky130_fd_sc_hd__a22o_1 _16961_ (.A1(\cpuregs[13][22] ),
    .A2(_13206_),
    .B1(_13209_),
    .B2(_13208_),
    .X(_03231_));
 sky130_fd_sc_hd__clkbuf_2 _16962_ (.A(\cpuregs_wrdata[21] ),
    .X(_13210_));
 sky130_fd_sc_hd__a22o_1 _16963_ (.A1(\cpuregs[13][21] ),
    .A2(_13206_),
    .B1(_13210_),
    .B2(_13208_),
    .X(_03230_));
 sky130_fd_sc_hd__clkbuf_2 _16964_ (.A(\cpuregs_wrdata[20] ),
    .X(_13211_));
 sky130_fd_sc_hd__a22o_1 _16965_ (.A1(\cpuregs[13][20] ),
    .A2(_13206_),
    .B1(_13211_),
    .B2(_13208_),
    .X(_03229_));
 sky130_fd_sc_hd__buf_1 _16966_ (.A(_13191_),
    .X(_13212_));
 sky130_fd_sc_hd__clkbuf_2 _16967_ (.A(\cpuregs_wrdata[19] ),
    .X(_13213_));
 sky130_fd_sc_hd__buf_1 _16968_ (.A(_13195_),
    .X(_13214_));
 sky130_fd_sc_hd__a22o_1 _16969_ (.A1(\cpuregs[13][19] ),
    .A2(_13212_),
    .B1(_13213_),
    .B2(_13214_),
    .X(_03228_));
 sky130_fd_sc_hd__clkbuf_2 _16970_ (.A(\cpuregs_wrdata[18] ),
    .X(_13215_));
 sky130_fd_sc_hd__a22o_1 _16971_ (.A1(\cpuregs[13][18] ),
    .A2(_13212_),
    .B1(_13215_),
    .B2(_13214_),
    .X(_03227_));
 sky130_fd_sc_hd__clkbuf_2 _16972_ (.A(\cpuregs_wrdata[17] ),
    .X(_13216_));
 sky130_fd_sc_hd__a22o_1 _16973_ (.A1(\cpuregs[13][17] ),
    .A2(_13212_),
    .B1(_13216_),
    .B2(_13214_),
    .X(_03226_));
 sky130_fd_sc_hd__clkbuf_2 _16974_ (.A(\cpuregs_wrdata[16] ),
    .X(_13217_));
 sky130_fd_sc_hd__a22o_1 _16975_ (.A1(\cpuregs[13][16] ),
    .A2(_13212_),
    .B1(_13217_),
    .B2(_13214_),
    .X(_03225_));
 sky130_fd_sc_hd__buf_2 _16976_ (.A(_13190_),
    .X(_13218_));
 sky130_fd_sc_hd__buf_1 _16977_ (.A(_13218_),
    .X(_13219_));
 sky130_fd_sc_hd__clkbuf_2 _16978_ (.A(\cpuregs_wrdata[15] ),
    .X(_13220_));
 sky130_fd_sc_hd__buf_2 _16979_ (.A(_13194_),
    .X(_13221_));
 sky130_fd_sc_hd__buf_1 _16980_ (.A(_13221_),
    .X(_13222_));
 sky130_fd_sc_hd__a22o_1 _16981_ (.A1(\cpuregs[13][15] ),
    .A2(_13219_),
    .B1(_13220_),
    .B2(_13222_),
    .X(_03224_));
 sky130_fd_sc_hd__clkbuf_2 _16982_ (.A(\cpuregs_wrdata[14] ),
    .X(_13223_));
 sky130_fd_sc_hd__a22o_1 _16983_ (.A1(\cpuregs[13][14] ),
    .A2(_13219_),
    .B1(_13223_),
    .B2(_13222_),
    .X(_03223_));
 sky130_fd_sc_hd__clkbuf_2 _16984_ (.A(\cpuregs_wrdata[13] ),
    .X(_13224_));
 sky130_fd_sc_hd__a22o_1 _16985_ (.A1(\cpuregs[13][13] ),
    .A2(_13219_),
    .B1(_13224_),
    .B2(_13222_),
    .X(_03222_));
 sky130_fd_sc_hd__clkbuf_2 _16986_ (.A(\cpuregs_wrdata[12] ),
    .X(_13225_));
 sky130_fd_sc_hd__a22o_1 _16987_ (.A1(\cpuregs[13][12] ),
    .A2(_13219_),
    .B1(_13225_),
    .B2(_13222_),
    .X(_03221_));
 sky130_fd_sc_hd__buf_1 _16988_ (.A(_13218_),
    .X(_13226_));
 sky130_fd_sc_hd__clkbuf_2 _16989_ (.A(\cpuregs_wrdata[11] ),
    .X(_13227_));
 sky130_fd_sc_hd__buf_1 _16990_ (.A(_13221_),
    .X(_13228_));
 sky130_fd_sc_hd__a22o_1 _16991_ (.A1(\cpuregs[13][11] ),
    .A2(_13226_),
    .B1(_13227_),
    .B2(_13228_),
    .X(_03220_));
 sky130_fd_sc_hd__clkbuf_2 _16992_ (.A(\cpuregs_wrdata[10] ),
    .X(_13229_));
 sky130_fd_sc_hd__a22o_1 _16993_ (.A1(\cpuregs[13][10] ),
    .A2(_13226_),
    .B1(_13229_),
    .B2(_13228_),
    .X(_03219_));
 sky130_fd_sc_hd__clkbuf_2 _16994_ (.A(\cpuregs_wrdata[9] ),
    .X(_13230_));
 sky130_fd_sc_hd__a22o_1 _16995_ (.A1(\cpuregs[13][9] ),
    .A2(_13226_),
    .B1(_13230_),
    .B2(_13228_),
    .X(_03218_));
 sky130_fd_sc_hd__clkbuf_2 _16996_ (.A(\cpuregs_wrdata[8] ),
    .X(_13231_));
 sky130_fd_sc_hd__a22o_1 _16997_ (.A1(\cpuregs[13][8] ),
    .A2(_13226_),
    .B1(_13231_),
    .B2(_13228_),
    .X(_03217_));
 sky130_fd_sc_hd__buf_1 _16998_ (.A(_13218_),
    .X(_13232_));
 sky130_fd_sc_hd__clkbuf_2 _16999_ (.A(\cpuregs_wrdata[7] ),
    .X(_13233_));
 sky130_fd_sc_hd__buf_1 _17000_ (.A(_13221_),
    .X(_13234_));
 sky130_fd_sc_hd__a22o_1 _17001_ (.A1(\cpuregs[13][7] ),
    .A2(_13232_),
    .B1(_13233_),
    .B2(_13234_),
    .X(_03216_));
 sky130_fd_sc_hd__clkbuf_2 _17002_ (.A(\cpuregs_wrdata[6] ),
    .X(_13235_));
 sky130_fd_sc_hd__a22o_1 _17003_ (.A1(\cpuregs[13][6] ),
    .A2(_13232_),
    .B1(_13235_),
    .B2(_13234_),
    .X(_03215_));
 sky130_fd_sc_hd__clkbuf_2 _17004_ (.A(\cpuregs_wrdata[5] ),
    .X(_13236_));
 sky130_fd_sc_hd__a22o_1 _17005_ (.A1(\cpuregs[13][5] ),
    .A2(_13232_),
    .B1(_13236_),
    .B2(_13234_),
    .X(_03214_));
 sky130_fd_sc_hd__clkbuf_2 _17006_ (.A(\cpuregs_wrdata[4] ),
    .X(_13237_));
 sky130_fd_sc_hd__a22o_1 _17007_ (.A1(\cpuregs[13][4] ),
    .A2(_13232_),
    .B1(_13237_),
    .B2(_13234_),
    .X(_03213_));
 sky130_fd_sc_hd__buf_1 _17008_ (.A(_13218_),
    .X(_13238_));
 sky130_fd_sc_hd__clkbuf_2 _17009_ (.A(\cpuregs_wrdata[3] ),
    .X(_13239_));
 sky130_fd_sc_hd__buf_1 _17010_ (.A(_13221_),
    .X(_13240_));
 sky130_fd_sc_hd__a22o_1 _17011_ (.A1(\cpuregs[13][3] ),
    .A2(_13238_),
    .B1(_13239_),
    .B2(_13240_),
    .X(_03212_));
 sky130_fd_sc_hd__clkbuf_2 _17012_ (.A(\cpuregs_wrdata[2] ),
    .X(_13241_));
 sky130_fd_sc_hd__a22o_1 _17013_ (.A1(\cpuregs[13][2] ),
    .A2(_13238_),
    .B1(_13241_),
    .B2(_13240_),
    .X(_03211_));
 sky130_fd_sc_hd__clkbuf_2 _17014_ (.A(\cpuregs_wrdata[1] ),
    .X(_13242_));
 sky130_fd_sc_hd__a22o_1 _17015_ (.A1(\cpuregs[13][1] ),
    .A2(_13238_),
    .B1(_13242_),
    .B2(_13240_),
    .X(_03210_));
 sky130_fd_sc_hd__clkbuf_2 _17016_ (.A(\cpuregs_wrdata[0] ),
    .X(_13243_));
 sky130_fd_sc_hd__a22o_1 _17017_ (.A1(\cpuregs[13][0] ),
    .A2(_13238_),
    .B1(_13243_),
    .B2(_13240_),
    .X(_03209_));
 sky130_fd_sc_hd__buf_1 _17018_ (.A(_00328_),
    .X(_13244_));
 sky130_fd_sc_hd__o32a_1 _17019_ (.A1(_11888_),
    .A2(_13244_),
    .A3(_13186_),
    .B1(_11801_),
    .B2(_13188_),
    .X(_13245_));
 sky130_vsdinv _17020_ (.A(_13245_),
    .Y(_03208_));
 sky130_fd_sc_hd__clkbuf_2 _17021_ (.A(_11922_),
    .X(_13246_));
 sky130_fd_sc_hd__buf_2 _17022_ (.A(_13246_),
    .X(_13247_));
 sky130_fd_sc_hd__a31oi_2 _17023_ (.A1(_00335_),
    .A2(_11940_),
    .A3(_11944_),
    .B1(_11961_),
    .Y(_13248_));
 sky130_fd_sc_hd__buf_2 _17024_ (.A(_11931_),
    .X(_13249_));
 sky130_fd_sc_hd__clkbuf_4 _17025_ (.A(_13249_),
    .X(_13250_));
 sky130_fd_sc_hd__o32a_1 _17026_ (.A1(_11812_),
    .A2(_13247_),
    .A3(_13248_),
    .B1(is_jalr_addi_slti_sltiu_xori_ori_andi),
    .B2(_13250_),
    .X(_03207_));
 sky130_fd_sc_hd__buf_2 _17027_ (.A(is_slli_srli_srai),
    .X(_13251_));
 sky130_fd_sc_hd__buf_2 _17028_ (.A(_13251_),
    .X(_13252_));
 sky130_fd_sc_hd__buf_2 _17029_ (.A(_13246_),
    .X(_13253_));
 sky130_fd_sc_hd__buf_2 _17030_ (.A(_13253_),
    .X(_13254_));
 sky130_fd_sc_hd__clkbuf_2 _17031_ (.A(_11921_),
    .X(_13255_));
 sky130_fd_sc_hd__o31a_1 _17032_ (.A1(_13255_),
    .A2(_00334_),
    .A3(_11927_),
    .B1(_11910_),
    .X(_13256_));
 sky130_fd_sc_hd__or4_4 _17033_ (.A(_11947_),
    .B(_11905_),
    .C(_11960_),
    .D(_13246_),
    .X(_13257_));
 sky130_fd_sc_hd__o2bb2ai_1 _17034_ (.A1_N(_13252_),
    .A2_N(_13254_),
    .B1(_13256_),
    .B2(_13257_),
    .Y(_03206_));
 sky130_fd_sc_hd__o32a_1 _17035_ (.A1(_11887_),
    .A2(_13244_),
    .A3(_13186_),
    .B1(_11797_),
    .B2(_13188_),
    .X(_13258_));
 sky130_vsdinv _17036_ (.A(_13258_),
    .Y(_03205_));
 sky130_fd_sc_hd__buf_1 _17037_ (.A(\decoded_imm_uj[20] ),
    .X(_13259_));
 sky130_fd_sc_hd__buf_1 _17038_ (.A(_13259_),
    .X(_13260_));
 sky130_fd_sc_hd__buf_1 _17039_ (.A(_13260_),
    .X(_13261_));
 sky130_fd_sc_hd__clkbuf_2 _17040_ (.A(_13261_),
    .X(_13262_));
 sky130_fd_sc_hd__clkbuf_4 _17041_ (.A(_13262_),
    .X(_13263_));
 sky130_fd_sc_hd__clkbuf_2 _17042_ (.A(_11895_),
    .X(_13264_));
 sky130_fd_sc_hd__a22o_2 _17043_ (.A1(_13263_),
    .A2(_13264_),
    .B1(\mem_rdata_latched[31] ),
    .B2(_14286_),
    .X(_03204_));
 sky130_fd_sc_hd__buf_1 _17044_ (.A(_11601_),
    .X(_13265_));
 sky130_fd_sc_hd__a22o_1 _17045_ (.A1(\decoded_imm_uj[19] ),
    .A2(_13264_),
    .B1(\mem_rdata_latched[19] ),
    .B2(_13265_),
    .X(_03203_));
 sky130_fd_sc_hd__buf_1 _17046_ (.A(_11892_),
    .X(_13266_));
 sky130_fd_sc_hd__clkbuf_2 _17047_ (.A(_11602_),
    .X(_13267_));
 sky130_fd_sc_hd__a22o_1 _17048_ (.A1(\mem_rdata_latched[18] ),
    .A2(_13266_),
    .B1(\decoded_imm_uj[18] ),
    .B2(_13267_),
    .X(_03202_));
 sky130_fd_sc_hd__buf_1 _17049_ (.A(_11892_),
    .X(_13268_));
 sky130_fd_sc_hd__a22o_1 _17050_ (.A1(\mem_rdata_latched[17] ),
    .A2(_13268_),
    .B1(\decoded_imm_uj[17] ),
    .B2(_13267_),
    .X(_03201_));
 sky130_fd_sc_hd__a22o_1 _17051_ (.A1(\mem_rdata_latched[16] ),
    .A2(_13268_),
    .B1(\decoded_imm_uj[16] ),
    .B2(_13267_),
    .X(_03200_));
 sky130_fd_sc_hd__a22o_1 _17052_ (.A1(\mem_rdata_latched[15] ),
    .A2(_13268_),
    .B1(\decoded_imm_uj[15] ),
    .B2(_13264_),
    .X(_03199_));
 sky130_fd_sc_hd__buf_1 _17053_ (.A(_11895_),
    .X(_13269_));
 sky130_fd_sc_hd__a22o_1 _17054_ (.A1(\decoded_imm_uj[14] ),
    .A2(_13269_),
    .B1(\mem_rdata_latched[14] ),
    .B2(_13265_),
    .X(_03198_));
 sky130_fd_sc_hd__a22o_1 _17055_ (.A1(\decoded_imm_uj[13] ),
    .A2(_13269_),
    .B1(\mem_rdata_latched[13] ),
    .B2(_13265_),
    .X(_03197_));
 sky130_fd_sc_hd__a22o_1 _17056_ (.A1(\decoded_imm_uj[12] ),
    .A2(_13269_),
    .B1(\mem_rdata_latched[12] ),
    .B2(_13265_),
    .X(_03196_));
 sky130_fd_sc_hd__buf_1 _17057_ (.A(_11601_),
    .X(_13270_));
 sky130_fd_sc_hd__a22o_1 _17058_ (.A1(\decoded_imm_uj[11] ),
    .A2(_13269_),
    .B1(\mem_rdata_latched[20] ),
    .B2(_13270_),
    .X(_03195_));
 sky130_fd_sc_hd__buf_1 _17059_ (.A(_11895_),
    .X(_13271_));
 sky130_fd_sc_hd__a22o_1 _17060_ (.A1(\decoded_imm_uj[10] ),
    .A2(_13271_),
    .B1(\mem_rdata_latched[30] ),
    .B2(_13270_),
    .X(_03194_));
 sky130_fd_sc_hd__a22o_1 _17061_ (.A1(\decoded_imm_uj[9] ),
    .A2(_13271_),
    .B1(\mem_rdata_latched[29] ),
    .B2(_13270_),
    .X(_03193_));
 sky130_fd_sc_hd__a22o_1 _17062_ (.A1(\decoded_imm_uj[8] ),
    .A2(_13271_),
    .B1(\mem_rdata_latched[28] ),
    .B2(_13270_),
    .X(_03192_));
 sky130_fd_sc_hd__a22o_1 _17063_ (.A1(\mem_rdata_latched[27] ),
    .A2(_13268_),
    .B1(\decoded_imm_uj[7] ),
    .B2(_13264_),
    .X(_03191_));
 sky130_fd_sc_hd__buf_1 _17064_ (.A(\decoded_imm_uj[6] ),
    .X(_13272_));
 sky130_fd_sc_hd__buf_1 _17065_ (.A(_11601_),
    .X(_13273_));
 sky130_fd_sc_hd__a22o_1 _17066_ (.A1(_13272_),
    .A2(_13271_),
    .B1(\mem_rdata_latched[26] ),
    .B2(_13273_),
    .X(_03190_));
 sky130_fd_sc_hd__buf_1 _17067_ (.A(_11885_),
    .X(_13274_));
 sky130_fd_sc_hd__a22o_1 _17068_ (.A1(\decoded_imm_uj[5] ),
    .A2(_13274_),
    .B1(\mem_rdata_latched[25] ),
    .B2(_13273_),
    .X(_03189_));
 sky130_fd_sc_hd__a22o_1 _17069_ (.A1(\decoded_imm_uj[4] ),
    .A2(_13274_),
    .B1(\mem_rdata_latched[24] ),
    .B2(_13273_),
    .X(_03188_));
 sky130_fd_sc_hd__a22o_1 _17070_ (.A1(\decoded_imm_uj[3] ),
    .A2(_13274_),
    .B1(\mem_rdata_latched[23] ),
    .B2(_13273_),
    .X(_03187_));
 sky130_fd_sc_hd__buf_1 _17071_ (.A(_11892_),
    .X(_13275_));
 sky130_fd_sc_hd__a22o_1 _17072_ (.A1(\decoded_imm_uj[2] ),
    .A2(_13274_),
    .B1(\mem_rdata_latched[22] ),
    .B2(_13275_),
    .X(_03186_));
 sky130_fd_sc_hd__buf_1 _17073_ (.A(_11885_),
    .X(_13276_));
 sky130_fd_sc_hd__a22o_1 _17074_ (.A1(\decoded_imm_uj[1] ),
    .A2(_13276_),
    .B1(\mem_rdata_latched[21] ),
    .B2(_13275_),
    .X(_03185_));
 sky130_vsdinv _17075_ (.A(\decoded_imm[0] ),
    .Y(_13277_));
 sky130_fd_sc_hd__clkbuf_2 _17076_ (.A(_13277_),
    .X(_13278_));
 sky130_fd_sc_hd__buf_1 _17077_ (.A(_11955_),
    .X(_13279_));
 sky130_fd_sc_hd__buf_2 _17078_ (.A(_13279_),
    .X(_13280_));
 sky130_vsdinv _17079_ (.A(\mem_rdata_q[7] ),
    .Y(_13281_));
 sky130_vsdinv _17080_ (.A(\mem_rdata_q[20] ),
    .Y(_13282_));
 sky130_fd_sc_hd__or3_4 _17081_ (.A(is_alu_reg_imm),
    .B(is_lb_lh_lw_lbu_lhu),
    .C(_11812_),
    .X(_13283_));
 sky130_vsdinv _17082_ (.A(_13283_),
    .Y(_13284_));
 sky130_fd_sc_hd__buf_1 _17083_ (.A(_13284_),
    .X(_13285_));
 sky130_fd_sc_hd__o22a_1 _17084_ (.A1(_11801_),
    .A2(_13281_),
    .B1(_13282_),
    .B2(_13285_),
    .X(_13286_));
 sky130_fd_sc_hd__o22ai_1 _17085_ (.A1(_13278_),
    .A2(_13280_),
    .B1(_13254_),
    .B2(_13286_),
    .Y(_03184_));
 sky130_fd_sc_hd__a22o_1 _17086_ (.A1(\decoded_rd[4] ),
    .A2(_13276_),
    .B1(\mem_rdata_latched[11] ),
    .B2(_13275_),
    .X(_03183_));
 sky130_fd_sc_hd__a22o_1 _17087_ (.A1(\decoded_rd[3] ),
    .A2(_13276_),
    .B1(\mem_rdata_latched[10] ),
    .B2(_13275_),
    .X(_03182_));
 sky130_fd_sc_hd__a22o_1 _17088_ (.A1(\decoded_rd[2] ),
    .A2(_13276_),
    .B1(\mem_rdata_latched[9] ),
    .B2(_13266_),
    .X(_03181_));
 sky130_fd_sc_hd__a22o_1 _17089_ (.A1(\decoded_rd[1] ),
    .A2(_11886_),
    .B1(\mem_rdata_latched[8] ),
    .B2(_13266_),
    .X(_03180_));
 sky130_fd_sc_hd__a22o_1 _17090_ (.A1(\decoded_rd[0] ),
    .A2(_11886_),
    .B1(\mem_rdata_latched[7] ),
    .B2(_13266_),
    .X(_03179_));
 sky130_vsdinv _17091_ (.A(\mem_rdata_q[27] ),
    .Y(_13287_));
 sky130_fd_sc_hd__or2_1 _17092_ (.A(_13287_),
    .B(_11922_),
    .X(_13288_));
 sky130_vsdinv _17093_ (.A(\mem_rdata_q[1] ),
    .Y(_13289_));
 sky130_vsdinv _17094_ (.A(\mem_rdata_q[0] ),
    .Y(_13290_));
 sky130_fd_sc_hd__or4_4 _17095_ (.A(_13289_),
    .B(_13290_),
    .C(\mem_rdata_q[6] ),
    .D(\mem_rdata_q[5] ),
    .X(_13291_));
 sky130_fd_sc_hd__or4b_4 _17096_ (.A(\mem_rdata_q[4] ),
    .B(_13291_),
    .C(\mem_rdata_q[2] ),
    .D_N(\mem_rdata_q[3] ),
    .X(_13292_));
 sky130_fd_sc_hd__buf_1 _17097_ (.A(\mem_rdata_q[28] ),
    .X(_13293_));
 sky130_fd_sc_hd__buf_2 _17098_ (.A(_13293_),
    .X(_13294_));
 sky130_fd_sc_hd__clkbuf_2 _17099_ (.A(\mem_rdata_q[26] ),
    .X(_13295_));
 sky130_vsdinv _17100_ (.A(\mem_rdata_q[25] ),
    .Y(_13296_));
 sky130_fd_sc_hd__or4_4 _17101_ (.A(\mem_rdata_q[31] ),
    .B(_11924_),
    .C(_11921_),
    .D(_13296_),
    .X(_13297_));
 sky130_fd_sc_hd__or3_1 _17102_ (.A(_13294_),
    .B(_13295_),
    .C(_13297_),
    .X(_13298_));
 sky130_vsdinv _17103_ (.A(instr_timer),
    .Y(_13299_));
 sky130_fd_sc_hd__buf_2 _17104_ (.A(_13299_),
    .X(_13300_));
 sky130_fd_sc_hd__clkbuf_4 _17105_ (.A(_11931_),
    .X(_13301_));
 sky130_fd_sc_hd__o32a_1 _17106_ (.A1(_13288_),
    .A2(_13292_),
    .A3(_13298_),
    .B1(_13300_),
    .B2(_13301_),
    .X(_13302_));
 sky130_vsdinv _17107_ (.A(_13302_),
    .Y(_03178_));
 sky130_fd_sc_hd__nor2_1 _17108_ (.A(_11608_),
    .B(_11611_),
    .Y(_13303_));
 sky130_fd_sc_hd__a32o_1 _17109_ (.A1(\mem_rdata_latched[27] ),
    .A2(_11614_),
    .A3(_13303_),
    .B1(instr_waitirq),
    .B2(_11897_),
    .X(_03177_));
 sky130_vsdinv _17110_ (.A(\mem_rdata_q[26] ),
    .Y(_13304_));
 sky130_fd_sc_hd__clkbuf_2 _17111_ (.A(\mem_rdata_q[27] ),
    .X(_13305_));
 sky130_fd_sc_hd__or4_4 _17112_ (.A(_13304_),
    .B(_11922_),
    .C(_13293_),
    .D(_13305_),
    .X(_13306_));
 sky130_fd_sc_hd__buf_2 _17113_ (.A(_11815_),
    .X(_13307_));
 sky130_fd_sc_hd__o32a_1 _17114_ (.A1(_13297_),
    .A2(_13306_),
    .A3(_13292_),
    .B1(_13307_),
    .B2(_13301_),
    .X(_13308_));
 sky130_vsdinv _17115_ (.A(_13308_),
    .Y(_03176_));
 sky130_fd_sc_hd__a2bb2o_1 _17116_ (.A1_N(_00337_),
    .A2_N(_11894_),
    .B1(_11568_),
    .B2(_00337_),
    .X(_03175_));
 sky130_fd_sc_hd__buf_2 _17117_ (.A(_13249_),
    .X(_13309_));
 sky130_fd_sc_hd__or4_4 _17118_ (.A(_13305_),
    .B(_11997_),
    .C(_13292_),
    .D(_13298_),
    .X(_13310_));
 sky130_fd_sc_hd__o21ai_1 _17119_ (.A1(_12873_),
    .A2(_13309_),
    .B1(_13310_),
    .Y(_03174_));
 sky130_fd_sc_hd__buf_1 _17120_ (.A(_11900_),
    .X(_13311_));
 sky130_fd_sc_hd__buf_2 _17121_ (.A(_13311_),
    .X(_13312_));
 sky130_vsdinv _17122_ (.A(_11911_),
    .Y(_13313_));
 sky130_vsdinv _17123_ (.A(_13292_),
    .Y(_13314_));
 sky130_fd_sc_hd__a22o_1 _17124_ (.A1(instr_getq),
    .A2(_13312_),
    .B1(_13313_),
    .B2(_13314_),
    .X(_03173_));
 sky130_fd_sc_hd__clkbuf_2 _17125_ (.A(\mem_rdata_q[21] ),
    .X(_13315_));
 sky130_fd_sc_hd__or2_1 _17126_ (.A(\mem_rdata_q[23] ),
    .B(\mem_rdata_q[22] ),
    .X(_13316_));
 sky130_fd_sc_hd__or4_4 _17127_ (.A(\mem_rdata_q[11] ),
    .B(\mem_rdata_q[10] ),
    .C(\mem_rdata_q[8] ),
    .D(\mem_rdata_q[7] ),
    .X(_13317_));
 sky130_fd_sc_hd__or4_4 _17128_ (.A(\mem_rdata_q[24] ),
    .B(_13315_),
    .C(_13316_),
    .D(_13317_),
    .X(_13318_));
 sky130_fd_sc_hd__or4_4 _17129_ (.A(\mem_rdata_q[9] ),
    .B(_13246_),
    .C(_11950_),
    .D(_13318_),
    .X(_13319_));
 sky130_fd_sc_hd__or2_1 _17130_ (.A(\mem_rdata_q[19] ),
    .B(\mem_rdata_q[18] ),
    .X(_13320_));
 sky130_fd_sc_hd__or4_4 _17131_ (.A(\mem_rdata_q[17] ),
    .B(\mem_rdata_q[16] ),
    .C(\mem_rdata_q[15] ),
    .D(_13320_),
    .X(_13321_));
 sky130_fd_sc_hd__or4bb_4 _17132_ (.A(_13289_),
    .B(_13290_),
    .C_N(\mem_rdata_q[6] ),
    .D_N(\mem_rdata_q[5] ),
    .X(_13322_));
 sky130_fd_sc_hd__or4b_4 _17133_ (.A(_13322_),
    .B(\mem_rdata_q[3] ),
    .C(\mem_rdata_q[2] ),
    .D_N(\mem_rdata_q[4] ),
    .X(_13323_));
 sky130_fd_sc_hd__or3_1 _17134_ (.A(_11910_),
    .B(_13321_),
    .C(_13323_),
    .X(_13324_));
 sky130_fd_sc_hd__o2bb2ai_1 _17135_ (.A1_N(instr_ecall_ebreak),
    .A2_N(_13254_),
    .B1(_13319_),
    .B2(_13324_),
    .Y(_03172_));
 sky130_vsdinv _17136_ (.A(\mem_rdata_q[21] ),
    .Y(_13325_));
 sky130_fd_sc_hd__or2_1 _17137_ (.A(_13325_),
    .B(_13316_),
    .X(_13326_));
 sky130_fd_sc_hd__or4_4 _17138_ (.A(\mem_rdata_q[20] ),
    .B(_11899_),
    .C(_13326_),
    .D(_13323_),
    .X(_13327_));
 sky130_vsdinv _17139_ (.A(\mem_rdata_q[31] ),
    .Y(_13328_));
 sky130_fd_sc_hd__or4_4 _17140_ (.A(_13328_),
    .B(_11925_),
    .C(_11921_),
    .D(_13293_),
    .X(_13329_));
 sky130_fd_sc_hd__buf_1 _17141_ (.A(\mem_rdata_q[25] ),
    .X(_13330_));
 sky130_fd_sc_hd__or2_1 _17142_ (.A(_13330_),
    .B(\mem_rdata_q[24] ),
    .X(_13331_));
 sky130_fd_sc_hd__or4_4 _17143_ (.A(_13329_),
    .B(_13331_),
    .C(_13287_),
    .D(\mem_rdata_q[26] ),
    .X(_13332_));
 sky130_fd_sc_hd__or2_2 _17144_ (.A(_11943_),
    .B(_13321_),
    .X(_13333_));
 sky130_fd_sc_hd__buf_2 _17145_ (.A(_11741_),
    .X(_13334_));
 sky130_fd_sc_hd__clkbuf_2 _17146_ (.A(_11931_),
    .X(_13335_));
 sky130_fd_sc_hd__o32a_1 _17147_ (.A1(_13327_),
    .A2(_13332_),
    .A3(_13333_),
    .B1(_13334_),
    .B2(_13335_),
    .X(_13336_));
 sky130_vsdinv _17148_ (.A(_13336_),
    .Y(_03171_));
 sky130_fd_sc_hd__clkbuf_2 _17149_ (.A(_11742_),
    .X(_13337_));
 sky130_fd_sc_hd__clkbuf_2 _17150_ (.A(\mem_rdata_q[24] ),
    .X(_13338_));
 sky130_fd_sc_hd__clkbuf_4 _17151_ (.A(_13328_),
    .X(_13339_));
 sky130_fd_sc_hd__or3_2 _17152_ (.A(\mem_rdata_q[29] ),
    .B(_13293_),
    .C(_13330_),
    .X(_13340_));
 sky130_fd_sc_hd__or4_4 _17153_ (.A(_13339_),
    .B(_11926_),
    .C(_13340_),
    .D(\mem_rdata_q[27] ),
    .X(_13341_));
 sky130_fd_sc_hd__or4_4 _17154_ (.A(_13295_),
    .B(_13338_),
    .C(_13333_),
    .D(_13341_),
    .X(_13342_));
 sky130_fd_sc_hd__o22ai_1 _17155_ (.A1(_13337_),
    .A2(_13280_),
    .B1(_13327_),
    .B2(_13342_),
    .Y(_03170_));
 sky130_fd_sc_hd__or4_4 _17156_ (.A(_13315_),
    .B(_11899_),
    .C(_13316_),
    .D(_13323_),
    .X(_13343_));
 sky130_fd_sc_hd__clkbuf_2 _17157_ (.A(_11743_),
    .X(_13344_));
 sky130_fd_sc_hd__o32a_1 _17158_ (.A1(_13332_),
    .A2(_13343_),
    .A3(_13333_),
    .B1(_13344_),
    .B2(_13335_),
    .X(_13345_));
 sky130_vsdinv _17159_ (.A(_13345_),
    .Y(_03169_));
 sky130_fd_sc_hd__buf_2 _17160_ (.A(_11999_),
    .X(_13346_));
 sky130_fd_sc_hd__o22ai_1 _17161_ (.A1(_11740_),
    .A2(_13346_),
    .B1(_13342_),
    .B2(_13343_),
    .Y(_03168_));
 sky130_vsdinv _17162_ (.A(_11920_),
    .Y(_13347_));
 sky130_vsdinv _17163_ (.A(_11928_),
    .Y(_13348_));
 sky130_fd_sc_hd__buf_1 _17164_ (.A(_11942_),
    .X(_13349_));
 sky130_fd_sc_hd__a32o_1 _17165_ (.A1(_11959_),
    .A2(_13347_),
    .A3(_13348_),
    .B1(instr_srai),
    .B2(_13349_),
    .X(_03167_));
 sky130_fd_sc_hd__a32o_1 _17166_ (.A1(_11959_),
    .A2(_13347_),
    .A3(_13313_),
    .B1(instr_srli),
    .B2(_13349_),
    .X(_03166_));
 sky130_vsdinv _17167_ (.A(_11948_),
    .Y(_13350_));
 sky130_fd_sc_hd__a32o_1 _17168_ (.A1(_11959_),
    .A2(_13350_),
    .A3(_13313_),
    .B1(instr_slli),
    .B2(_13349_),
    .X(_03165_));
 sky130_vsdinv _17169_ (.A(instr_sw),
    .Y(_13351_));
 sky130_fd_sc_hd__o32a_1 _17170_ (.A1(_11801_),
    .A2(_11997_),
    .A3(_11944_),
    .B1(_13351_),
    .B2(_13335_),
    .X(_13352_));
 sky130_vsdinv _17171_ (.A(_13352_),
    .Y(_03164_));
 sky130_fd_sc_hd__clkbuf_2 _17172_ (.A(is_sb_sh_sw),
    .X(_13353_));
 sky130_fd_sc_hd__buf_2 _17173_ (.A(_11955_),
    .X(_13354_));
 sky130_fd_sc_hd__buf_1 _17174_ (.A(_13354_),
    .X(_13355_));
 sky130_fd_sc_hd__a32o_1 _17175_ (.A1(_13353_),
    .A2(_13355_),
    .A3(_13350_),
    .B1(instr_sh),
    .B2(_13349_),
    .X(_03163_));
 sky130_vsdinv _17176_ (.A(_11951_),
    .Y(_13356_));
 sky130_fd_sc_hd__buf_1 _17177_ (.A(_13311_),
    .X(_13357_));
 sky130_fd_sc_hd__a32o_1 _17178_ (.A1(_13353_),
    .A2(_13355_),
    .A3(_13356_),
    .B1(instr_sb),
    .B2(_13357_),
    .X(_03162_));
 sky130_fd_sc_hd__buf_1 _17179_ (.A(is_lb_lh_lw_lbu_lhu),
    .X(_13358_));
 sky130_fd_sc_hd__a32o_1 _17180_ (.A1(_13358_),
    .A2(_13355_),
    .A3(_13347_),
    .B1(instr_lhu),
    .B2(_13357_),
    .X(_03161_));
 sky130_vsdinv _17181_ (.A(_11937_),
    .Y(_13359_));
 sky130_fd_sc_hd__a32o_1 _17182_ (.A1(_13358_),
    .A2(_13355_),
    .A3(_13359_),
    .B1(instr_lbu),
    .B2(_13357_),
    .X(_03160_));
 sky130_vsdinv _17183_ (.A(instr_lw),
    .Y(_13360_));
 sky130_fd_sc_hd__o32a_1 _17184_ (.A1(_11797_),
    .A2(_11997_),
    .A3(_11943_),
    .B1(_13360_),
    .B2(_13335_),
    .X(_13361_));
 sky130_vsdinv _17185_ (.A(_13361_),
    .Y(_03159_));
 sky130_fd_sc_hd__buf_2 _17186_ (.A(_13354_),
    .X(_13362_));
 sky130_fd_sc_hd__a32o_1 _17187_ (.A1(_13358_),
    .A2(_13362_),
    .A3(_13350_),
    .B1(instr_lh),
    .B2(_13357_),
    .X(_03158_));
 sky130_fd_sc_hd__clkbuf_2 _17188_ (.A(_13311_),
    .X(_13363_));
 sky130_fd_sc_hd__a32o_1 _17189_ (.A1(_13358_),
    .A2(_13362_),
    .A3(_13356_),
    .B1(instr_lb),
    .B2(_13363_),
    .X(_03157_));
 sky130_fd_sc_hd__or3b_1 _17190_ (.A(_11605_),
    .B(_11606_),
    .C_N(_00326_),
    .X(_13364_));
 sky130_fd_sc_hd__or2_2 _17191_ (.A(_00327_),
    .B(_13364_),
    .X(_13365_));
 sky130_fd_sc_hd__or4_4 _17192_ (.A(\mem_rdata_latched[14] ),
    .B(\mem_rdata_latched[13] ),
    .C(\mem_rdata_latched[12] ),
    .D(_11889_),
    .X(_13366_));
 sky130_vsdinv _17193_ (.A(_11812_),
    .Y(_02063_));
 sky130_fd_sc_hd__o32a_1 _17194_ (.A1(_13365_),
    .A2(_13366_),
    .A3(_11885_),
    .B1(_02063_),
    .B2(_13188_),
    .X(_13367_));
 sky130_vsdinv _17195_ (.A(_13367_),
    .Y(_03156_));
 sky130_vsdinv _17196_ (.A(instr_jal),
    .Y(_13368_));
 sky130_fd_sc_hd__buf_2 _17197_ (.A(_13368_),
    .X(_13369_));
 sky130_fd_sc_hd__clkbuf_2 _17198_ (.A(_13369_),
    .X(_13370_));
 sky130_fd_sc_hd__clkbuf_2 _17199_ (.A(_13370_),
    .X(_00323_));
 sky130_fd_sc_hd__or3_1 _17200_ (.A(_11603_),
    .B(_11889_),
    .C(_13364_),
    .X(_13371_));
 sky130_fd_sc_hd__o22ai_1 _17201_ (.A1(_00323_),
    .A2(_14286_),
    .B1(_11896_),
    .B2(_13371_),
    .Y(_03155_));
 sky130_fd_sc_hd__nor3_4 _17202_ (.A(_00330_),
    .B(_11886_),
    .C(_13365_),
    .Y(_13372_));
 sky130_fd_sc_hd__a32o_1 _17203_ (.A1(_11888_),
    .A2(_13244_),
    .A3(_13372_),
    .B1(instr_auipc),
    .B2(_11897_),
    .X(_03154_));
 sky130_fd_sc_hd__buf_2 _17204_ (.A(instr_lui),
    .X(_13373_));
 sky130_fd_sc_hd__a32o_1 _17205_ (.A1(_11887_),
    .A2(_13244_),
    .A3(_13372_),
    .B1(_13373_),
    .B2(_13267_),
    .X(_03153_));
 sky130_fd_sc_hd__clkbuf_2 _17206_ (.A(_13311_),
    .X(_13374_));
 sky130_fd_sc_hd__buf_1 _17207_ (.A(_11955_),
    .X(_13375_));
 sky130_fd_sc_hd__buf_2 _17208_ (.A(_13375_),
    .X(_13376_));
 sky130_fd_sc_hd__a22o_1 _17209_ (.A1(net298),
    .A2(_13374_),
    .B1(_11923_),
    .B2(_13376_),
    .X(_03152_));
 sky130_fd_sc_hd__a22o_1 _17210_ (.A1(net297),
    .A2(_13374_),
    .B1(_11924_),
    .B2(_13376_),
    .X(_03151_));
 sky130_fd_sc_hd__o22a_1 _17211_ (.A1(_13255_),
    .A2(_13363_),
    .B1(net295),
    .B2(_13309_),
    .X(_03150_));
 sky130_fd_sc_hd__a22o_1 _17212_ (.A1(net294),
    .A2(_13374_),
    .B1(_13294_),
    .B2(_13376_),
    .X(_03149_));
 sky130_fd_sc_hd__o22a_1 _17213_ (.A1(_13305_),
    .A2(_13363_),
    .B1(net293),
    .B2(_13309_),
    .X(_03148_));
 sky130_fd_sc_hd__clkbuf_2 _17214_ (.A(_13375_),
    .X(_13377_));
 sky130_fd_sc_hd__a22o_1 _17215_ (.A1(_13295_),
    .A2(_13377_),
    .B1(net292),
    .B2(_13363_),
    .X(_03147_));
 sky130_fd_sc_hd__clkbuf_2 _17216_ (.A(_13279_),
    .X(_13378_));
 sky130_fd_sc_hd__a22o_1 _17217_ (.A1(net291),
    .A2(_13374_),
    .B1(_13330_),
    .B2(_13378_),
    .X(_03146_));
 sky130_fd_sc_hd__clkbuf_2 _17218_ (.A(_11900_),
    .X(_13379_));
 sky130_fd_sc_hd__buf_1 _17219_ (.A(_13379_),
    .X(_13380_));
 sky130_fd_sc_hd__a22o_1 _17220_ (.A1(net290),
    .A2(_13380_),
    .B1(_13338_),
    .B2(_13378_),
    .X(_03145_));
 sky130_fd_sc_hd__a22o_1 _17221_ (.A1(net289),
    .A2(_13380_),
    .B1(\mem_rdata_q[23] ),
    .B2(_13378_),
    .X(_03144_));
 sky130_fd_sc_hd__a22o_1 _17222_ (.A1(net288),
    .A2(_13380_),
    .B1(\mem_rdata_q[22] ),
    .B2(_13378_),
    .X(_03143_));
 sky130_fd_sc_hd__o22a_1 _17223_ (.A1(_13315_),
    .A2(_13312_),
    .B1(net287),
    .B2(_13309_),
    .X(_03142_));
 sky130_fd_sc_hd__o22a_1 _17224_ (.A1(\mem_rdata_q[20] ),
    .A2(_13312_),
    .B1(net286),
    .B2(_13250_),
    .X(_03141_));
 sky130_fd_sc_hd__clkbuf_2 _17225_ (.A(_13279_),
    .X(_13381_));
 sky130_fd_sc_hd__a22o_1 _17226_ (.A1(net284),
    .A2(_13380_),
    .B1(\mem_rdata_q[19] ),
    .B2(_13381_),
    .X(_03140_));
 sky130_fd_sc_hd__buf_1 _17227_ (.A(_13379_),
    .X(_13382_));
 sky130_fd_sc_hd__a22o_1 _17228_ (.A1(net283),
    .A2(_13382_),
    .B1(\mem_rdata_q[18] ),
    .B2(_13381_),
    .X(_03139_));
 sky130_fd_sc_hd__a22o_1 _17229_ (.A1(net282),
    .A2(_13382_),
    .B1(\mem_rdata_q[17] ),
    .B2(_13381_),
    .X(_03138_));
 sky130_fd_sc_hd__a22o_1 _17230_ (.A1(net281),
    .A2(_13382_),
    .B1(\mem_rdata_q[16] ),
    .B2(_13381_),
    .X(_03137_));
 sky130_fd_sc_hd__clkbuf_2 _17231_ (.A(_13279_),
    .X(_13383_));
 sky130_fd_sc_hd__a22o_1 _17232_ (.A1(net280),
    .A2(_13382_),
    .B1(\mem_rdata_q[15] ),
    .B2(_13383_),
    .X(_03136_));
 sky130_fd_sc_hd__buf_1 _17233_ (.A(_13379_),
    .X(_13384_));
 sky130_fd_sc_hd__a22o_1 _17234_ (.A1(net279),
    .A2(_13384_),
    .B1(_11939_),
    .B2(_13383_),
    .X(_03135_));
 sky130_fd_sc_hd__a22o_1 _17235_ (.A1(net278),
    .A2(_13384_),
    .B1(_11947_),
    .B2(_13383_),
    .X(_03134_));
 sky130_fd_sc_hd__a22o_1 _17236_ (.A1(net277),
    .A2(_13384_),
    .B1(_11915_),
    .B2(_13383_),
    .X(_03133_));
 sky130_fd_sc_hd__buf_1 _17237_ (.A(_13375_),
    .X(_13385_));
 sky130_fd_sc_hd__a22o_1 _17238_ (.A1(net276),
    .A2(_13384_),
    .B1(\mem_rdata_q[11] ),
    .B2(_13385_),
    .X(_03132_));
 sky130_fd_sc_hd__buf_1 _17239_ (.A(_13379_),
    .X(_13386_));
 sky130_fd_sc_hd__a22o_1 _17240_ (.A1(net275),
    .A2(_13386_),
    .B1(\mem_rdata_q[10] ),
    .B2(_13385_),
    .X(_03131_));
 sky130_fd_sc_hd__o22a_1 _17241_ (.A1(\mem_rdata_q[9] ),
    .A2(_13312_),
    .B1(net305),
    .B2(_13250_),
    .X(_03130_));
 sky130_fd_sc_hd__a22o_1 _17242_ (.A1(net304),
    .A2(_13386_),
    .B1(\mem_rdata_q[8] ),
    .B2(_13385_),
    .X(_03129_));
 sky130_fd_sc_hd__a22o_1 _17243_ (.A1(net303),
    .A2(_13386_),
    .B1(\mem_rdata_q[7] ),
    .B2(_13385_),
    .X(_03128_));
 sky130_fd_sc_hd__buf_1 _17244_ (.A(_13375_),
    .X(_13387_));
 sky130_fd_sc_hd__a22o_1 _17245_ (.A1(net302),
    .A2(_13386_),
    .B1(\mem_rdata_q[6] ),
    .B2(_13387_),
    .X(_03127_));
 sky130_fd_sc_hd__clkbuf_2 _17246_ (.A(_11963_),
    .X(_13388_));
 sky130_fd_sc_hd__a22o_1 _17247_ (.A1(net301),
    .A2(_13388_),
    .B1(\mem_rdata_q[5] ),
    .B2(_13387_),
    .X(_03126_));
 sky130_fd_sc_hd__a22o_1 _17248_ (.A1(net300),
    .A2(_13388_),
    .B1(\mem_rdata_q[4] ),
    .B2(_13387_),
    .X(_03125_));
 sky130_fd_sc_hd__a22o_1 _17249_ (.A1(net299),
    .A2(_13388_),
    .B1(\mem_rdata_q[3] ),
    .B2(_13387_),
    .X(_03124_));
 sky130_fd_sc_hd__a22o_1 _17250_ (.A1(net296),
    .A2(_13388_),
    .B1(\mem_rdata_q[2] ),
    .B2(_13377_),
    .X(_03123_));
 sky130_fd_sc_hd__a22o_1 _17251_ (.A1(net285),
    .A2(_13247_),
    .B1(\mem_rdata_q[1] ),
    .B2(_13377_),
    .X(_03122_));
 sky130_fd_sc_hd__a22o_1 _17252_ (.A1(net274),
    .A2(_13247_),
    .B1(\mem_rdata_q[0] ),
    .B2(_13377_),
    .X(_03121_));
 sky130_vsdinv _17253_ (.A(\cpu_state[5] ),
    .Y(_13389_));
 sky130_fd_sc_hd__and3_1 _17254_ (.A(_11569_),
    .B(_11559_),
    .C(_13389_),
    .X(_13390_));
 sky130_fd_sc_hd__or4_4 _17255_ (.A(_11580_),
    .B(_00318_),
    .C(_00320_),
    .D(_13390_),
    .X(_13391_));
 sky130_fd_sc_hd__buf_2 _17256_ (.A(_13391_),
    .X(_13392_));
 sky130_fd_sc_hd__buf_1 _17257_ (.A(_13392_),
    .X(_13393_));
 sky130_fd_sc_hd__buf_2 _17258_ (.A(_11682_),
    .X(_13394_));
 sky130_vsdinv _17259_ (.A(_13391_),
    .Y(_13395_));
 sky130_fd_sc_hd__buf_2 _17260_ (.A(_13395_),
    .X(_13396_));
 sky130_fd_sc_hd__buf_1 _17261_ (.A(_13396_),
    .X(_13397_));
 sky130_fd_sc_hd__o22a_1 _17262_ (.A1(_02499_),
    .A2(_13393_),
    .B1(_13394_),
    .B2(_13397_),
    .X(_03120_));
 sky130_fd_sc_hd__buf_1 _17263_ (.A(net329),
    .X(_13398_));
 sky130_fd_sc_hd__buf_2 _17264_ (.A(_13398_),
    .X(_13399_));
 sky130_fd_sc_hd__o22a_1 _17265_ (.A1(_02498_),
    .A2(_13393_),
    .B1(_13399_),
    .B2(_13397_),
    .X(_03119_));
 sky130_fd_sc_hd__clkbuf_2 _17266_ (.A(net327),
    .X(_13400_));
 sky130_fd_sc_hd__buf_1 _17267_ (.A(_13400_),
    .X(_13401_));
 sky130_fd_sc_hd__buf_2 _17268_ (.A(_13401_),
    .X(_13402_));
 sky130_fd_sc_hd__o22a_1 _17269_ (.A1(_02496_),
    .A2(_13393_),
    .B1(_13402_),
    .B2(_13397_),
    .X(_03118_));
 sky130_fd_sc_hd__clkbuf_2 _17270_ (.A(net326),
    .X(_13403_));
 sky130_fd_sc_hd__buf_1 _17271_ (.A(_13403_),
    .X(_13404_));
 sky130_fd_sc_hd__buf_2 _17272_ (.A(_13404_),
    .X(_13405_));
 sky130_fd_sc_hd__o22a_1 _17273_ (.A1(_02495_),
    .A2(_13393_),
    .B1(_13405_),
    .B2(_13397_),
    .X(_03117_));
 sky130_fd_sc_hd__buf_1 _17274_ (.A(_13392_),
    .X(_13406_));
 sky130_fd_sc_hd__clkbuf_2 _17275_ (.A(net325),
    .X(_13407_));
 sky130_fd_sc_hd__clkbuf_4 _17276_ (.A(_13407_),
    .X(_13408_));
 sky130_fd_sc_hd__buf_1 _17277_ (.A(_13396_),
    .X(_13409_));
 sky130_fd_sc_hd__o22a_1 _17278_ (.A1(_02494_),
    .A2(_13406_),
    .B1(_13408_),
    .B2(_13409_),
    .X(_03116_));
 sky130_fd_sc_hd__buf_1 _17279_ (.A(net324),
    .X(_13410_));
 sky130_fd_sc_hd__buf_1 _17280_ (.A(_13410_),
    .X(_13411_));
 sky130_fd_sc_hd__clkbuf_4 _17281_ (.A(_13411_),
    .X(_13412_));
 sky130_fd_sc_hd__o22a_1 _17282_ (.A1(_02493_),
    .A2(_13406_),
    .B1(_13412_),
    .B2(_13409_),
    .X(_03115_));
 sky130_fd_sc_hd__buf_1 _17283_ (.A(net323),
    .X(_13413_));
 sky130_fd_sc_hd__clkbuf_4 _17284_ (.A(_13413_),
    .X(_13414_));
 sky130_fd_sc_hd__o22a_1 _17285_ (.A1(_02492_),
    .A2(_13406_),
    .B1(_13414_),
    .B2(_13409_),
    .X(_03114_));
 sky130_fd_sc_hd__buf_1 _17286_ (.A(net322),
    .X(_13415_));
 sky130_fd_sc_hd__clkbuf_2 _17287_ (.A(_13415_),
    .X(_13416_));
 sky130_fd_sc_hd__clkbuf_4 _17288_ (.A(_13416_),
    .X(_13417_));
 sky130_fd_sc_hd__o22a_1 _17289_ (.A1(_02491_),
    .A2(_13406_),
    .B1(_13417_),
    .B2(_13409_),
    .X(_03113_));
 sky130_fd_sc_hd__buf_1 _17290_ (.A(_13392_),
    .X(_13418_));
 sky130_fd_sc_hd__clkbuf_2 _17291_ (.A(net321),
    .X(_13419_));
 sky130_fd_sc_hd__buf_4 _17292_ (.A(_13419_),
    .X(_13420_));
 sky130_fd_sc_hd__buf_1 _17293_ (.A(_13396_),
    .X(_13421_));
 sky130_fd_sc_hd__o22a_1 _17294_ (.A1(_02490_),
    .A2(_13418_),
    .B1(_13420_),
    .B2(_13421_),
    .X(_03112_));
 sky130_fd_sc_hd__clkbuf_2 _17295_ (.A(net320),
    .X(_13422_));
 sky130_fd_sc_hd__buf_4 _17296_ (.A(_13422_),
    .X(_13423_));
 sky130_fd_sc_hd__o22a_1 _17297_ (.A1(_02489_),
    .A2(_13418_),
    .B1(_13423_),
    .B2(_13421_),
    .X(_03111_));
 sky130_fd_sc_hd__clkbuf_2 _17298_ (.A(net319),
    .X(_13424_));
 sky130_fd_sc_hd__buf_4 _17299_ (.A(_13424_),
    .X(_13425_));
 sky130_fd_sc_hd__o22a_1 _17300_ (.A1(_02488_),
    .A2(_13418_),
    .B1(_13425_),
    .B2(_13421_),
    .X(_03110_));
 sky130_fd_sc_hd__clkbuf_2 _17301_ (.A(net318),
    .X(_13426_));
 sky130_fd_sc_hd__buf_4 _17302_ (.A(_13426_),
    .X(_13427_));
 sky130_fd_sc_hd__o22a_1 _17303_ (.A1(_02487_),
    .A2(_13418_),
    .B1(_13427_),
    .B2(_13421_),
    .X(_03109_));
 sky130_fd_sc_hd__buf_1 _17304_ (.A(_13392_),
    .X(_13428_));
 sky130_fd_sc_hd__clkbuf_2 _17305_ (.A(net316),
    .X(_13429_));
 sky130_fd_sc_hd__buf_4 _17306_ (.A(_13429_),
    .X(_13430_));
 sky130_fd_sc_hd__buf_1 _17307_ (.A(_13396_),
    .X(_13431_));
 sky130_fd_sc_hd__o22a_1 _17308_ (.A1(_02485_),
    .A2(_13428_),
    .B1(_13430_),
    .B2(_13431_),
    .X(_03108_));
 sky130_fd_sc_hd__buf_1 _17309_ (.A(net315),
    .X(_13432_));
 sky130_fd_sc_hd__buf_4 _17310_ (.A(_13432_),
    .X(_13433_));
 sky130_fd_sc_hd__o22a_1 _17311_ (.A1(_02484_),
    .A2(_13428_),
    .B1(_13433_),
    .B2(_13431_),
    .X(_03107_));
 sky130_fd_sc_hd__buf_1 _17312_ (.A(net314),
    .X(_13434_));
 sky130_fd_sc_hd__clkbuf_4 _17313_ (.A(_13434_),
    .X(_13435_));
 sky130_fd_sc_hd__o22a_1 _17314_ (.A1(_02483_),
    .A2(_13428_),
    .B1(_13435_),
    .B2(_13431_),
    .X(_03106_));
 sky130_fd_sc_hd__buf_1 _17315_ (.A(net313),
    .X(_13436_));
 sky130_fd_sc_hd__buf_1 _17316_ (.A(_13436_),
    .X(_13437_));
 sky130_fd_sc_hd__clkbuf_4 _17317_ (.A(_13437_),
    .X(_13438_));
 sky130_fd_sc_hd__o22a_1 _17318_ (.A1(_02482_),
    .A2(_13428_),
    .B1(_13438_),
    .B2(_13431_),
    .X(_03105_));
 sky130_fd_sc_hd__clkbuf_2 _17319_ (.A(_13391_),
    .X(_13439_));
 sky130_fd_sc_hd__clkbuf_2 _17320_ (.A(_13439_),
    .X(_13440_));
 sky130_fd_sc_hd__clkbuf_2 _17321_ (.A(net312),
    .X(_13441_));
 sky130_fd_sc_hd__buf_4 _17322_ (.A(_13441_),
    .X(_13442_));
 sky130_fd_sc_hd__buf_2 _17323_ (.A(_13395_),
    .X(_13443_));
 sky130_fd_sc_hd__buf_1 _17324_ (.A(_13443_),
    .X(_13444_));
 sky130_fd_sc_hd__o22a_1 _17325_ (.A1(_02481_),
    .A2(_13440_),
    .B1(_13442_),
    .B2(_13444_),
    .X(_03104_));
 sky130_fd_sc_hd__clkbuf_2 _17326_ (.A(net311),
    .X(_13445_));
 sky130_fd_sc_hd__buf_4 _17327_ (.A(_13445_),
    .X(_13446_));
 sky130_fd_sc_hd__o22a_1 _17328_ (.A1(_02480_),
    .A2(_13440_),
    .B1(_13446_),
    .B2(_13444_),
    .X(_03103_));
 sky130_fd_sc_hd__clkbuf_2 _17329_ (.A(net310),
    .X(_13447_));
 sky130_fd_sc_hd__clkbuf_4 _17330_ (.A(_13447_),
    .X(_13448_));
 sky130_fd_sc_hd__o22a_1 _17331_ (.A1(_02479_),
    .A2(_13440_),
    .B1(_13448_),
    .B2(_13444_),
    .X(_03102_));
 sky130_fd_sc_hd__buf_1 _17332_ (.A(net309),
    .X(_13449_));
 sky130_fd_sc_hd__clkbuf_4 _17333_ (.A(_13449_),
    .X(_13450_));
 sky130_fd_sc_hd__o22a_1 _17334_ (.A1(_02478_),
    .A2(_13440_),
    .B1(_13450_),
    .B2(_13444_),
    .X(_03101_));
 sky130_fd_sc_hd__buf_1 _17335_ (.A(_13439_),
    .X(_13451_));
 sky130_fd_sc_hd__buf_1 _17336_ (.A(net308),
    .X(_13452_));
 sky130_fd_sc_hd__clkbuf_4 _17337_ (.A(_13452_),
    .X(_13453_));
 sky130_fd_sc_hd__buf_1 _17338_ (.A(_13443_),
    .X(_13454_));
 sky130_fd_sc_hd__o22a_1 _17339_ (.A1(_02477_),
    .A2(_13451_),
    .B1(_13453_),
    .B2(_13454_),
    .X(_03100_));
 sky130_fd_sc_hd__clkbuf_2 _17340_ (.A(net307),
    .X(_13455_));
 sky130_fd_sc_hd__clkbuf_4 _17341_ (.A(_13455_),
    .X(_13456_));
 sky130_fd_sc_hd__o22a_1 _17342_ (.A1(_02476_),
    .A2(_13451_),
    .B1(_13456_),
    .B2(_13454_),
    .X(_03099_));
 sky130_fd_sc_hd__buf_1 _17343_ (.A(net337),
    .X(_13457_));
 sky130_fd_sc_hd__clkbuf_4 _17344_ (.A(_13457_),
    .X(_13458_));
 sky130_fd_sc_hd__o22a_1 _17345_ (.A1(_02506_),
    .A2(_13451_),
    .B1(_13458_),
    .B2(_13454_),
    .X(_03098_));
 sky130_fd_sc_hd__buf_1 _17346_ (.A(net336),
    .X(_13459_));
 sky130_fd_sc_hd__buf_1 _17347_ (.A(_13459_),
    .X(_13460_));
 sky130_fd_sc_hd__buf_2 _17348_ (.A(_13460_),
    .X(_13461_));
 sky130_fd_sc_hd__o22a_1 _17349_ (.A1(_02505_),
    .A2(_13451_),
    .B1(_13461_),
    .B2(_13454_),
    .X(_03097_));
 sky130_fd_sc_hd__buf_1 _17350_ (.A(_13439_),
    .X(_13462_));
 sky130_fd_sc_hd__clkbuf_2 _17351_ (.A(net335),
    .X(_13463_));
 sky130_fd_sc_hd__clkbuf_2 _17352_ (.A(_13463_),
    .X(_13464_));
 sky130_fd_sc_hd__clkbuf_4 _17353_ (.A(_13464_),
    .X(_13465_));
 sky130_fd_sc_hd__buf_1 _17354_ (.A(_13443_),
    .X(_13466_));
 sky130_fd_sc_hd__o22a_1 _17355_ (.A1(_02504_),
    .A2(_13462_),
    .B1(_13465_),
    .B2(_13466_),
    .X(_03096_));
 sky130_fd_sc_hd__buf_1 _17356_ (.A(net334),
    .X(_13467_));
 sky130_fd_sc_hd__clkbuf_2 _17357_ (.A(_13467_),
    .X(_13468_));
 sky130_fd_sc_hd__buf_2 _17358_ (.A(_13468_),
    .X(_13469_));
 sky130_fd_sc_hd__o22a_1 _17359_ (.A1(_02503_),
    .A2(_13462_),
    .B1(_13469_),
    .B2(_13466_),
    .X(_03095_));
 sky130_fd_sc_hd__clkbuf_2 _17360_ (.A(net333),
    .X(_13470_));
 sky130_fd_sc_hd__clkbuf_2 _17361_ (.A(_13470_),
    .X(_13471_));
 sky130_fd_sc_hd__buf_2 _17362_ (.A(_13471_),
    .X(_13472_));
 sky130_fd_sc_hd__o22a_1 _17363_ (.A1(_02502_),
    .A2(_13462_),
    .B1(_13472_),
    .B2(_13466_),
    .X(_03094_));
 sky130_fd_sc_hd__clkbuf_2 _17364_ (.A(net332),
    .X(_13473_));
 sky130_fd_sc_hd__buf_1 _17365_ (.A(_13473_),
    .X(_13474_));
 sky130_fd_sc_hd__buf_2 _17366_ (.A(_13474_),
    .X(_13475_));
 sky130_fd_sc_hd__o22a_1 _17367_ (.A1(_02501_),
    .A2(_13462_),
    .B1(_13475_),
    .B2(_13466_),
    .X(_03093_));
 sky130_fd_sc_hd__buf_1 _17368_ (.A(_13439_),
    .X(_13476_));
 sky130_fd_sc_hd__clkbuf_2 _17369_ (.A(net331),
    .X(_13477_));
 sky130_fd_sc_hd__buf_1 _17370_ (.A(_13477_),
    .X(_13478_));
 sky130_fd_sc_hd__buf_2 _17371_ (.A(_13478_),
    .X(_13479_));
 sky130_fd_sc_hd__buf_1 _17372_ (.A(_13443_),
    .X(_13480_));
 sky130_fd_sc_hd__o22a_1 _17373_ (.A1(_02500_),
    .A2(_13476_),
    .B1(_13479_),
    .B2(_13480_),
    .X(_03092_));
 sky130_fd_sc_hd__buf_1 _17374_ (.A(net328),
    .X(_13481_));
 sky130_fd_sc_hd__clkbuf_2 _17375_ (.A(_13481_),
    .X(_13482_));
 sky130_fd_sc_hd__buf_2 _17376_ (.A(_13482_),
    .X(_13483_));
 sky130_fd_sc_hd__o22a_1 _17377_ (.A1(_02497_),
    .A2(_13476_),
    .B1(_13483_),
    .B2(_13480_),
    .X(_03091_));
 sky130_fd_sc_hd__clkbuf_2 _17378_ (.A(net317),
    .X(_13484_));
 sky130_fd_sc_hd__buf_4 _17379_ (.A(_13484_),
    .X(_13485_));
 sky130_fd_sc_hd__clkbuf_4 _17380_ (.A(_13485_),
    .X(_13486_));
 sky130_fd_sc_hd__o22a_1 _17381_ (.A1(_02486_),
    .A2(_13476_),
    .B1(_13486_),
    .B2(_13480_),
    .X(_03090_));
 sky130_fd_sc_hd__buf_2 _17382_ (.A(net306),
    .X(_13487_));
 sky130_fd_sc_hd__buf_2 _17383_ (.A(_13487_),
    .X(_13488_));
 sky130_fd_sc_hd__o22a_1 _17384_ (.A1(_02475_),
    .A2(_13476_),
    .B1(_13488_),
    .B2(_13480_),
    .X(_03089_));
 sky130_fd_sc_hd__buf_6 _17385_ (.A(_11882_),
    .X(_13489_));
 sky130_fd_sc_hd__a22o_1 _17386_ (.A1(net158),
    .A2(_11884_),
    .B1(net191),
    .B2(_13489_),
    .X(_03088_));
 sky130_fd_sc_hd__a22o_1 _17387_ (.A1(net157),
    .A2(_11884_),
    .B1(net190),
    .B2(_13489_),
    .X(_03087_));
 sky130_fd_sc_hd__a22o_1 _17388_ (.A1(net155),
    .A2(_11884_),
    .B1(net188),
    .B2(_13489_),
    .X(_03086_));
 sky130_fd_sc_hd__buf_2 _17389_ (.A(_11883_),
    .X(_13490_));
 sky130_fd_sc_hd__clkbuf_2 _17390_ (.A(_13490_),
    .X(_13491_));
 sky130_fd_sc_hd__a22o_1 _17391_ (.A1(net154),
    .A2(_13491_),
    .B1(net187),
    .B2(_13489_),
    .X(_03085_));
 sky130_fd_sc_hd__buf_1 _17392_ (.A(_11881_),
    .X(_13492_));
 sky130_fd_sc_hd__buf_2 _17393_ (.A(_13492_),
    .X(_13493_));
 sky130_fd_sc_hd__a22o_1 _17394_ (.A1(net153),
    .A2(_13491_),
    .B1(net186),
    .B2(_13493_),
    .X(_03084_));
 sky130_fd_sc_hd__a22o_1 _17395_ (.A1(net152),
    .A2(_13491_),
    .B1(net185),
    .B2(_13493_),
    .X(_03083_));
 sky130_fd_sc_hd__a22o_1 _17396_ (.A1(net151),
    .A2(_13491_),
    .B1(net184),
    .B2(_13493_),
    .X(_03082_));
 sky130_fd_sc_hd__clkbuf_2 _17397_ (.A(_11883_),
    .X(_13494_));
 sky130_fd_sc_hd__buf_1 _17398_ (.A(_13494_),
    .X(_13495_));
 sky130_fd_sc_hd__a22o_1 _17399_ (.A1(net150),
    .A2(_13495_),
    .B1(net183),
    .B2(_13493_),
    .X(_03081_));
 sky130_fd_sc_hd__buf_1 _17400_ (.A(_13492_),
    .X(_13496_));
 sky130_fd_sc_hd__a22o_1 _17401_ (.A1(net149),
    .A2(_13495_),
    .B1(net182),
    .B2(_13496_),
    .X(_03080_));
 sky130_fd_sc_hd__a22o_1 _17402_ (.A1(net148),
    .A2(_13495_),
    .B1(net181),
    .B2(_13496_),
    .X(_03079_));
 sky130_fd_sc_hd__a22o_1 _17403_ (.A1(net147),
    .A2(_13495_),
    .B1(net180),
    .B2(_13496_),
    .X(_03078_));
 sky130_fd_sc_hd__clkbuf_2 _17404_ (.A(_13494_),
    .X(_13497_));
 sky130_fd_sc_hd__a22o_1 _17405_ (.A1(net146),
    .A2(_13497_),
    .B1(net179),
    .B2(_13496_),
    .X(_03077_));
 sky130_fd_sc_hd__clkbuf_2 _17406_ (.A(_13492_),
    .X(_13498_));
 sky130_fd_sc_hd__a22o_1 _17407_ (.A1(net144),
    .A2(_13497_),
    .B1(net177),
    .B2(_13498_),
    .X(_03076_));
 sky130_fd_sc_hd__a22o_1 _17408_ (.A1(net143),
    .A2(_13497_),
    .B1(net176),
    .B2(_13498_),
    .X(_03075_));
 sky130_fd_sc_hd__a22o_1 _17409_ (.A1(net142),
    .A2(_13497_),
    .B1(net175),
    .B2(_13498_),
    .X(_03074_));
 sky130_fd_sc_hd__clkbuf_4 _17410_ (.A(_13494_),
    .X(_13499_));
 sky130_fd_sc_hd__a22o_1 _17411_ (.A1(net141),
    .A2(_13499_),
    .B1(net174),
    .B2(_13498_),
    .X(_03073_));
 sky130_fd_sc_hd__clkbuf_4 _17412_ (.A(_13492_),
    .X(_13500_));
 sky130_fd_sc_hd__a22o_1 _17413_ (.A1(net140),
    .A2(_13499_),
    .B1(net173),
    .B2(_13500_),
    .X(_03072_));
 sky130_fd_sc_hd__a22o_1 _17414_ (.A1(net139),
    .A2(_13499_),
    .B1(net172),
    .B2(_13500_),
    .X(_03071_));
 sky130_fd_sc_hd__a22o_1 _17415_ (.A1(net138),
    .A2(_13499_),
    .B1(net171),
    .B2(_13500_),
    .X(_03070_));
 sky130_fd_sc_hd__buf_4 _17416_ (.A(_13494_),
    .X(_13501_));
 sky130_fd_sc_hd__a22o_1 _17417_ (.A1(net137),
    .A2(_13501_),
    .B1(net170),
    .B2(_13500_),
    .X(_03069_));
 sky130_fd_sc_hd__buf_6 _17418_ (.A(_11881_),
    .X(_13502_));
 sky130_fd_sc_hd__a22o_1 _17419_ (.A1(net136),
    .A2(_13501_),
    .B1(net169),
    .B2(_13502_),
    .X(_03068_));
 sky130_fd_sc_hd__a22o_1 _17420_ (.A1(net135),
    .A2(_13501_),
    .B1(net168),
    .B2(_13502_),
    .X(_03067_));
 sky130_fd_sc_hd__a22o_1 _17421_ (.A1(net165),
    .A2(_13501_),
    .B1(net198),
    .B2(_13502_),
    .X(_03066_));
 sky130_fd_sc_hd__clkbuf_4 _17422_ (.A(_11883_),
    .X(_13503_));
 sky130_fd_sc_hd__a22o_1 _17423_ (.A1(net164),
    .A2(_13503_),
    .B1(net197),
    .B2(_13502_),
    .X(_03065_));
 sky130_fd_sc_hd__buf_2 _17424_ (.A(_11881_),
    .X(_13504_));
 sky130_fd_sc_hd__a22o_1 _17425_ (.A1(net163),
    .A2(_13503_),
    .B1(net196),
    .B2(_13504_),
    .X(_03064_));
 sky130_fd_sc_hd__a22o_1 _17426_ (.A1(net162),
    .A2(_13503_),
    .B1(net195),
    .B2(_13504_),
    .X(_03063_));
 sky130_fd_sc_hd__a22o_1 _17427_ (.A1(net161),
    .A2(_13503_),
    .B1(net194),
    .B2(_13504_),
    .X(_03062_));
 sky130_fd_sc_hd__a22o_1 _17428_ (.A1(net160),
    .A2(_13490_),
    .B1(net193),
    .B2(_13504_),
    .X(_03061_));
 sky130_fd_sc_hd__a22o_1 _17429_ (.A1(net159),
    .A2(_13490_),
    .B1(net192),
    .B2(_11882_),
    .X(_03060_));
 sky130_fd_sc_hd__a22o_1 _17430_ (.A1(net156),
    .A2(_13490_),
    .B1(net189),
    .B2(_11882_),
    .X(_03059_));
 sky130_fd_sc_hd__buf_1 _17431_ (.A(\pcpi_mul.rs1[31] ),
    .X(_13505_));
 sky130_fd_sc_hd__buf_1 _17432_ (.A(_13505_),
    .X(_13506_));
 sky130_fd_sc_hd__clkbuf_2 _17433_ (.A(_13506_),
    .X(_13507_));
 sky130_fd_sc_hd__clkbuf_2 _17434_ (.A(_13507_),
    .X(_13508_));
 sky130_fd_sc_hd__a22o_1 _17435_ (.A1(_13394_),
    .A2(_11710_),
    .B1(_13508_),
    .B2(_13070_),
    .X(_03058_));
 sky130_fd_sc_hd__buf_1 _17436_ (.A(\pcpi_mul.rs1[30] ),
    .X(_13509_));
 sky130_fd_sc_hd__buf_1 _17437_ (.A(_13509_),
    .X(_13510_));
 sky130_fd_sc_hd__clkbuf_2 _17438_ (.A(_13510_),
    .X(_13511_));
 sky130_fd_sc_hd__clkbuf_2 _17439_ (.A(_13511_),
    .X(_13512_));
 sky130_fd_sc_hd__buf_1 _17440_ (.A(_13512_),
    .X(_13513_));
 sky130_fd_sc_hd__buf_1 _17441_ (.A(_13139_),
    .X(_13514_));
 sky130_fd_sc_hd__a22o_1 _17442_ (.A1(_13513_),
    .A2(_13182_),
    .B1(_13399_),
    .B2(_13514_),
    .X(_03057_));
 sky130_fd_sc_hd__buf_1 _17443_ (.A(\pcpi_mul.rs1[29] ),
    .X(_13515_));
 sky130_fd_sc_hd__clkbuf_2 _17444_ (.A(_13515_),
    .X(_13516_));
 sky130_fd_sc_hd__clkbuf_2 _17445_ (.A(_13516_),
    .X(_13517_));
 sky130_fd_sc_hd__buf_1 _17446_ (.A(_13517_),
    .X(_13518_));
 sky130_fd_sc_hd__a22o_1 _17447_ (.A1(_13518_),
    .A2(_13182_),
    .B1(_13402_),
    .B2(_13514_),
    .X(_03056_));
 sky130_fd_sc_hd__buf_1 _17448_ (.A(\pcpi_mul.rs1[28] ),
    .X(_13519_));
 sky130_fd_sc_hd__clkbuf_2 _17449_ (.A(_13519_),
    .X(_13520_));
 sky130_fd_sc_hd__clkbuf_2 _17450_ (.A(_13520_),
    .X(_13521_));
 sky130_fd_sc_hd__buf_1 _17451_ (.A(_13521_),
    .X(_13522_));
 sky130_fd_sc_hd__a22o_1 _17452_ (.A1(_13522_),
    .A2(_13182_),
    .B1(_13405_),
    .B2(_13514_),
    .X(_03055_));
 sky130_fd_sc_hd__buf_1 _17453_ (.A(\pcpi_mul.rs1[27] ),
    .X(_13523_));
 sky130_fd_sc_hd__buf_1 _17454_ (.A(_13523_),
    .X(_13524_));
 sky130_fd_sc_hd__buf_1 _17455_ (.A(_13524_),
    .X(_13525_));
 sky130_fd_sc_hd__buf_1 _17456_ (.A(_13525_),
    .X(_13526_));
 sky130_fd_sc_hd__buf_1 _17457_ (.A(_13181_),
    .X(_13527_));
 sky130_fd_sc_hd__a22o_1 _17458_ (.A1(_13526_),
    .A2(_13527_),
    .B1(_13408_),
    .B2(_13514_),
    .X(_03054_));
 sky130_fd_sc_hd__buf_1 _17459_ (.A(\pcpi_mul.rs1[26] ),
    .X(_13528_));
 sky130_fd_sc_hd__buf_1 _17460_ (.A(_13528_),
    .X(_13529_));
 sky130_fd_sc_hd__buf_1 _17461_ (.A(_13529_),
    .X(_13530_));
 sky130_fd_sc_hd__buf_1 _17462_ (.A(_13530_),
    .X(_13531_));
 sky130_fd_sc_hd__clkbuf_2 _17463_ (.A(_11708_),
    .X(_13532_));
 sky130_fd_sc_hd__clkbuf_2 _17464_ (.A(_13532_),
    .X(_13533_));
 sky130_fd_sc_hd__a22o_1 _17465_ (.A1(_13531_),
    .A2(_13527_),
    .B1(_13412_),
    .B2(_13533_),
    .X(_03053_));
 sky130_fd_sc_hd__buf_1 _17466_ (.A(\pcpi_mul.rs1[25] ),
    .X(_13534_));
 sky130_fd_sc_hd__clkbuf_2 _17467_ (.A(_13534_),
    .X(_13535_));
 sky130_fd_sc_hd__buf_1 _17468_ (.A(_13535_),
    .X(_13536_));
 sky130_fd_sc_hd__buf_1 _17469_ (.A(_13536_),
    .X(_13537_));
 sky130_fd_sc_hd__a22o_1 _17470_ (.A1(_13537_),
    .A2(_13527_),
    .B1(_13414_),
    .B2(_13533_),
    .X(_03052_));
 sky130_fd_sc_hd__buf_1 _17471_ (.A(\pcpi_mul.rs1[24] ),
    .X(_13538_));
 sky130_fd_sc_hd__clkbuf_2 _17472_ (.A(_13538_),
    .X(_13539_));
 sky130_fd_sc_hd__buf_1 _17473_ (.A(_13539_),
    .X(_13540_));
 sky130_fd_sc_hd__a22o_1 _17474_ (.A1(_13540_),
    .A2(_13527_),
    .B1(_13417_),
    .B2(_13533_),
    .X(_03051_));
 sky130_fd_sc_hd__buf_1 _17475_ (.A(\pcpi_mul.rs1[23] ),
    .X(_13541_));
 sky130_fd_sc_hd__clkbuf_2 _17476_ (.A(_13541_),
    .X(_13542_));
 sky130_fd_sc_hd__clkbuf_2 _17477_ (.A(_13542_),
    .X(_13543_));
 sky130_fd_sc_hd__buf_1 _17478_ (.A(_13181_),
    .X(_13544_));
 sky130_fd_sc_hd__a22o_1 _17479_ (.A1(_13543_),
    .A2(_13544_),
    .B1(_13420_),
    .B2(_13533_),
    .X(_03050_));
 sky130_fd_sc_hd__buf_1 _17480_ (.A(\pcpi_mul.rs1[22] ),
    .X(_13545_));
 sky130_fd_sc_hd__clkbuf_2 _17481_ (.A(_13545_),
    .X(_13546_));
 sky130_fd_sc_hd__clkbuf_2 _17482_ (.A(_13546_),
    .X(_13547_));
 sky130_fd_sc_hd__buf_1 _17483_ (.A(_13532_),
    .X(_13548_));
 sky130_fd_sc_hd__a22o_1 _17484_ (.A1(_13547_),
    .A2(_13544_),
    .B1(_13423_),
    .B2(_13548_),
    .X(_03049_));
 sky130_fd_sc_hd__buf_1 _17485_ (.A(\pcpi_mul.rs1[21] ),
    .X(_13549_));
 sky130_fd_sc_hd__buf_1 _17486_ (.A(_13549_),
    .X(_13550_));
 sky130_fd_sc_hd__buf_2 _17487_ (.A(_13550_),
    .X(_13551_));
 sky130_fd_sc_hd__a22o_1 _17488_ (.A1(_13551_),
    .A2(_13544_),
    .B1(_13425_),
    .B2(_13548_),
    .X(_03048_));
 sky130_fd_sc_hd__buf_1 _17489_ (.A(\pcpi_mul.rs1[20] ),
    .X(_13552_));
 sky130_fd_sc_hd__buf_1 _17490_ (.A(_13552_),
    .X(_13553_));
 sky130_fd_sc_hd__clkbuf_2 _17491_ (.A(_13553_),
    .X(_13554_));
 sky130_fd_sc_hd__a22o_1 _17492_ (.A1(_13554_),
    .A2(_13544_),
    .B1(_13427_),
    .B2(_13548_),
    .X(_03047_));
 sky130_fd_sc_hd__buf_1 _17493_ (.A(\pcpi_mul.rs1[19] ),
    .X(_13555_));
 sky130_fd_sc_hd__clkbuf_2 _17494_ (.A(_13555_),
    .X(_13556_));
 sky130_fd_sc_hd__clkbuf_2 _17495_ (.A(_13556_),
    .X(_13557_));
 sky130_fd_sc_hd__clkbuf_2 _17496_ (.A(_13181_),
    .X(_13558_));
 sky130_fd_sc_hd__a22o_1 _17497_ (.A1(_13557_),
    .A2(_13558_),
    .B1(_13430_),
    .B2(_13548_),
    .X(_03046_));
 sky130_fd_sc_hd__buf_1 _17498_ (.A(\pcpi_mul.rs1[18] ),
    .X(_13559_));
 sky130_fd_sc_hd__buf_1 _17499_ (.A(_13559_),
    .X(_13560_));
 sky130_fd_sc_hd__clkbuf_2 _17500_ (.A(_13560_),
    .X(_13561_));
 sky130_fd_sc_hd__clkbuf_2 _17501_ (.A(_13532_),
    .X(_13562_));
 sky130_fd_sc_hd__a22o_1 _17502_ (.A1(_13561_),
    .A2(_13558_),
    .B1(_13433_),
    .B2(_13562_),
    .X(_03045_));
 sky130_fd_sc_hd__buf_1 _17503_ (.A(\pcpi_mul.rs1[17] ),
    .X(_13563_));
 sky130_fd_sc_hd__buf_1 _17504_ (.A(_13563_),
    .X(_13564_));
 sky130_fd_sc_hd__buf_2 _17505_ (.A(_13564_),
    .X(_13565_));
 sky130_fd_sc_hd__a22o_1 _17506_ (.A1(_13565_),
    .A2(_13558_),
    .B1(_13435_),
    .B2(_13562_),
    .X(_03044_));
 sky130_fd_sc_hd__buf_1 _17507_ (.A(\pcpi_mul.rs1[16] ),
    .X(_13566_));
 sky130_fd_sc_hd__buf_1 _17508_ (.A(_13566_),
    .X(_13567_));
 sky130_fd_sc_hd__buf_2 _17509_ (.A(_13567_),
    .X(_13568_));
 sky130_fd_sc_hd__a22o_1 _17510_ (.A1(_13568_),
    .A2(_13558_),
    .B1(_13438_),
    .B2(_13562_),
    .X(_03043_));
 sky130_fd_sc_hd__buf_1 _17511_ (.A(\pcpi_mul.rs1[15] ),
    .X(_13569_));
 sky130_fd_sc_hd__buf_1 _17512_ (.A(_13569_),
    .X(_13570_));
 sky130_fd_sc_hd__clkbuf_2 _17513_ (.A(_13570_),
    .X(_13571_));
 sky130_fd_sc_hd__clkbuf_2 _17514_ (.A(_11693_),
    .X(_13572_));
 sky130_fd_sc_hd__buf_1 _17515_ (.A(_13572_),
    .X(_13573_));
 sky130_fd_sc_hd__a22o_1 _17516_ (.A1(_13571_),
    .A2(_13573_),
    .B1(_13442_),
    .B2(_13562_),
    .X(_03042_));
 sky130_fd_sc_hd__buf_1 _17517_ (.A(\pcpi_mul.rs1[14] ),
    .X(_13574_));
 sky130_fd_sc_hd__buf_1 _17518_ (.A(_13574_),
    .X(_13575_));
 sky130_fd_sc_hd__clkbuf_2 _17519_ (.A(_13575_),
    .X(_13576_));
 sky130_fd_sc_hd__clkbuf_2 _17520_ (.A(_13532_),
    .X(_13577_));
 sky130_fd_sc_hd__a22o_1 _17521_ (.A1(_13576_),
    .A2(_13573_),
    .B1(_13446_),
    .B2(_13577_),
    .X(_03041_));
 sky130_fd_sc_hd__buf_1 _17522_ (.A(\pcpi_mul.rs1[13] ),
    .X(_13578_));
 sky130_fd_sc_hd__buf_1 _17523_ (.A(_13578_),
    .X(_13579_));
 sky130_fd_sc_hd__clkbuf_2 _17524_ (.A(_13579_),
    .X(_13580_));
 sky130_fd_sc_hd__a22o_1 _17525_ (.A1(_13580_),
    .A2(_13573_),
    .B1(_13448_),
    .B2(_13577_),
    .X(_03040_));
 sky130_fd_sc_hd__buf_1 _17526_ (.A(\pcpi_mul.rs1[12] ),
    .X(_13581_));
 sky130_fd_sc_hd__buf_1 _17527_ (.A(_13581_),
    .X(_13582_));
 sky130_fd_sc_hd__clkbuf_2 _17528_ (.A(_13582_),
    .X(_13583_));
 sky130_fd_sc_hd__a22o_1 _17529_ (.A1(_13583_),
    .A2(_13573_),
    .B1(_13450_),
    .B2(_13577_),
    .X(_03039_));
 sky130_fd_sc_hd__buf_1 _17530_ (.A(\pcpi_mul.rs1[11] ),
    .X(_13584_));
 sky130_fd_sc_hd__clkbuf_4 _17531_ (.A(_13584_),
    .X(_13585_));
 sky130_fd_sc_hd__buf_1 _17532_ (.A(_13572_),
    .X(_13586_));
 sky130_fd_sc_hd__a22o_1 _17533_ (.A1(_13585_),
    .A2(_13586_),
    .B1(_13453_),
    .B2(_13577_),
    .X(_03038_));
 sky130_fd_sc_hd__clkbuf_2 _17534_ (.A(\pcpi_mul.rs1[10] ),
    .X(_13587_));
 sky130_fd_sc_hd__buf_2 _17535_ (.A(_13587_),
    .X(_13588_));
 sky130_fd_sc_hd__buf_1 _17536_ (.A(_11709_),
    .X(_13589_));
 sky130_fd_sc_hd__a22o_1 _17537_ (.A1(_13588_),
    .A2(_13586_),
    .B1(_13456_),
    .B2(_13589_),
    .X(_03037_));
 sky130_fd_sc_hd__clkbuf_2 _17538_ (.A(\pcpi_mul.rs1[9] ),
    .X(_13590_));
 sky130_fd_sc_hd__clkbuf_2 _17539_ (.A(_13590_),
    .X(_13591_));
 sky130_fd_sc_hd__buf_2 _17540_ (.A(_13591_),
    .X(_13592_));
 sky130_fd_sc_hd__a22o_1 _17541_ (.A1(_13592_),
    .A2(_13586_),
    .B1(_13458_),
    .B2(_13589_),
    .X(_03036_));
 sky130_fd_sc_hd__clkbuf_2 _17542_ (.A(\pcpi_mul.rs1[8] ),
    .X(_13593_));
 sky130_fd_sc_hd__buf_1 _17543_ (.A(_13593_),
    .X(_13594_));
 sky130_fd_sc_hd__buf_2 _17544_ (.A(_13594_),
    .X(_13595_));
 sky130_fd_sc_hd__a22o_1 _17545_ (.A1(_13595_),
    .A2(_13586_),
    .B1(_13461_),
    .B2(_13589_),
    .X(_03035_));
 sky130_fd_sc_hd__clkbuf_2 _17546_ (.A(\pcpi_mul.rs1[7] ),
    .X(_13596_));
 sky130_fd_sc_hd__buf_1 _17547_ (.A(_13596_),
    .X(_13597_));
 sky130_fd_sc_hd__clkbuf_2 _17548_ (.A(_13597_),
    .X(_13598_));
 sky130_fd_sc_hd__buf_2 _17549_ (.A(_13598_),
    .X(_13599_));
 sky130_fd_sc_hd__buf_1 _17550_ (.A(_13572_),
    .X(_13600_));
 sky130_fd_sc_hd__a22o_1 _17551_ (.A1(_13599_),
    .A2(_13600_),
    .B1(_13465_),
    .B2(_13589_),
    .X(_03034_));
 sky130_fd_sc_hd__buf_1 _17552_ (.A(\pcpi_mul.rs1[6] ),
    .X(_13601_));
 sky130_fd_sc_hd__clkbuf_2 _17553_ (.A(_13601_),
    .X(_13602_));
 sky130_fd_sc_hd__buf_1 _17554_ (.A(_13602_),
    .X(_13603_));
 sky130_fd_sc_hd__buf_2 _17555_ (.A(_13603_),
    .X(_13604_));
 sky130_fd_sc_hd__buf_1 _17556_ (.A(_11709_),
    .X(_13605_));
 sky130_fd_sc_hd__a22o_1 _17557_ (.A1(_13604_),
    .A2(_13600_),
    .B1(_13469_),
    .B2(_13605_),
    .X(_03033_));
 sky130_fd_sc_hd__buf_1 _17558_ (.A(\pcpi_mul.rs1[5] ),
    .X(_13606_));
 sky130_fd_sc_hd__clkbuf_2 _17559_ (.A(_13606_),
    .X(_13607_));
 sky130_fd_sc_hd__clkbuf_2 _17560_ (.A(_13607_),
    .X(_13608_));
 sky130_fd_sc_hd__buf_2 _17561_ (.A(_13608_),
    .X(_13609_));
 sky130_fd_sc_hd__a22o_1 _17562_ (.A1(_13609_),
    .A2(_13600_),
    .B1(_13472_),
    .B2(_13605_),
    .X(_03032_));
 sky130_fd_sc_hd__buf_1 _17563_ (.A(\pcpi_mul.rs1[4] ),
    .X(_13610_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _17564_ (.A(_13610_),
    .X(_13611_));
 sky130_fd_sc_hd__buf_1 _17565_ (.A(_13611_),
    .X(_13612_));
 sky130_fd_sc_hd__buf_2 _17566_ (.A(_13612_),
    .X(_13613_));
 sky130_fd_sc_hd__a22o_1 _17567_ (.A1(_13613_),
    .A2(_13600_),
    .B1(_13475_),
    .B2(_13605_),
    .X(_03031_));
 sky130_fd_sc_hd__buf_1 _17568_ (.A(\pcpi_mul.rs1[3] ),
    .X(_13614_));
 sky130_fd_sc_hd__buf_1 _17569_ (.A(_13614_),
    .X(_13615_));
 sky130_fd_sc_hd__buf_2 _17570_ (.A(_13615_),
    .X(_13616_));
 sky130_fd_sc_hd__buf_1 _17571_ (.A(_13572_),
    .X(_13617_));
 sky130_fd_sc_hd__a22o_1 _17572_ (.A1(_13616_),
    .A2(_13617_),
    .B1(_13479_),
    .B2(_13605_),
    .X(_03030_));
 sky130_fd_sc_hd__buf_1 _17573_ (.A(\pcpi_mul.rs1[2] ),
    .X(_13618_));
 sky130_fd_sc_hd__buf_1 _17574_ (.A(_13618_),
    .X(_13619_));
 sky130_fd_sc_hd__buf_2 _17575_ (.A(_13619_),
    .X(_13620_));
 sky130_fd_sc_hd__a22o_1 _17576_ (.A1(_13620_),
    .A2(_13617_),
    .B1(_13483_),
    .B2(_13063_),
    .X(_03029_));
 sky130_fd_sc_hd__buf_1 _17577_ (.A(\pcpi_mul.rs1[1] ),
    .X(_13621_));
 sky130_fd_sc_hd__buf_1 _17578_ (.A(_13621_),
    .X(_13622_));
 sky130_fd_sc_hd__buf_1 _17579_ (.A(_13622_),
    .X(_13623_));
 sky130_fd_sc_hd__buf_2 _17580_ (.A(_13623_),
    .X(_13624_));
 sky130_fd_sc_hd__a22o_1 _17581_ (.A1(_13624_),
    .A2(_13617_),
    .B1(_13486_),
    .B2(_13063_),
    .X(_03028_));
 sky130_fd_sc_hd__buf_1 _17582_ (.A(\pcpi_mul.rs1[0] ),
    .X(_13625_));
 sky130_fd_sc_hd__buf_2 _17583_ (.A(_13625_),
    .X(_13626_));
 sky130_fd_sc_hd__a22o_1 _17584_ (.A1(_13626_),
    .A2(_13617_),
    .B1(_13488_),
    .B2(_13063_),
    .X(_03027_));
 sky130_fd_sc_hd__or2_2 _17585_ (.A(_12556_),
    .B(_12658_),
    .X(_13627_));
 sky130_fd_sc_hd__buf_4 _17586_ (.A(_13627_),
    .X(_13628_));
 sky130_fd_sc_hd__buf_1 _17587_ (.A(_13628_),
    .X(_13629_));
 sky130_vsdinv _17588_ (.A(_13627_),
    .Y(_13630_));
 sky130_fd_sc_hd__clkbuf_4 _17589_ (.A(_13630_),
    .X(_13631_));
 sky130_fd_sc_hd__buf_1 _17590_ (.A(_13631_),
    .X(_13632_));
 sky130_fd_sc_hd__a22o_1 _17591_ (.A1(\cpuregs[5][31] ),
    .A2(_13629_),
    .B1(_13193_),
    .B2(_13632_),
    .X(_03026_));
 sky130_fd_sc_hd__a22o_1 _17592_ (.A1(\cpuregs[5][30] ),
    .A2(_13629_),
    .B1(_13197_),
    .B2(_13632_),
    .X(_03025_));
 sky130_fd_sc_hd__a22o_1 _17593_ (.A1(\cpuregs[5][29] ),
    .A2(_13629_),
    .B1(_13198_),
    .B2(_13632_),
    .X(_03024_));
 sky130_fd_sc_hd__a22o_1 _17594_ (.A1(\cpuregs[5][28] ),
    .A2(_13629_),
    .B1(_13199_),
    .B2(_13632_),
    .X(_03023_));
 sky130_fd_sc_hd__buf_1 _17595_ (.A(_13628_),
    .X(_13633_));
 sky130_fd_sc_hd__buf_1 _17596_ (.A(_13631_),
    .X(_13634_));
 sky130_fd_sc_hd__a22o_1 _17597_ (.A1(\cpuregs[5][27] ),
    .A2(_13633_),
    .B1(_13201_),
    .B2(_13634_),
    .X(_03022_));
 sky130_fd_sc_hd__a22o_1 _17598_ (.A1(\cpuregs[5][26] ),
    .A2(_13633_),
    .B1(_13203_),
    .B2(_13634_),
    .X(_03021_));
 sky130_fd_sc_hd__a22o_1 _17599_ (.A1(\cpuregs[5][25] ),
    .A2(_13633_),
    .B1(_13204_),
    .B2(_13634_),
    .X(_03020_));
 sky130_fd_sc_hd__a22o_1 _17600_ (.A1(\cpuregs[5][24] ),
    .A2(_13633_),
    .B1(_13205_),
    .B2(_13634_),
    .X(_03019_));
 sky130_fd_sc_hd__buf_1 _17601_ (.A(_13628_),
    .X(_13635_));
 sky130_fd_sc_hd__buf_1 _17602_ (.A(_13631_),
    .X(_13636_));
 sky130_fd_sc_hd__a22o_1 _17603_ (.A1(\cpuregs[5][23] ),
    .A2(_13635_),
    .B1(_13207_),
    .B2(_13636_),
    .X(_03018_));
 sky130_fd_sc_hd__a22o_1 _17604_ (.A1(\cpuregs[5][22] ),
    .A2(_13635_),
    .B1(_13209_),
    .B2(_13636_),
    .X(_03017_));
 sky130_fd_sc_hd__a22o_1 _17605_ (.A1(\cpuregs[5][21] ),
    .A2(_13635_),
    .B1(_13210_),
    .B2(_13636_),
    .X(_03016_));
 sky130_fd_sc_hd__a22o_1 _17606_ (.A1(\cpuregs[5][20] ),
    .A2(_13635_),
    .B1(_13211_),
    .B2(_13636_),
    .X(_03015_));
 sky130_fd_sc_hd__buf_1 _17607_ (.A(_13628_),
    .X(_13637_));
 sky130_fd_sc_hd__buf_1 _17608_ (.A(_13631_),
    .X(_13638_));
 sky130_fd_sc_hd__a22o_1 _17609_ (.A1(\cpuregs[5][19] ),
    .A2(_13637_),
    .B1(_13213_),
    .B2(_13638_),
    .X(_03014_));
 sky130_fd_sc_hd__a22o_1 _17610_ (.A1(\cpuregs[5][18] ),
    .A2(_13637_),
    .B1(_13215_),
    .B2(_13638_),
    .X(_03013_));
 sky130_fd_sc_hd__a22o_1 _17611_ (.A1(\cpuregs[5][17] ),
    .A2(_13637_),
    .B1(_13216_),
    .B2(_13638_),
    .X(_03012_));
 sky130_fd_sc_hd__a22o_1 _17612_ (.A1(\cpuregs[5][16] ),
    .A2(_13637_),
    .B1(_13217_),
    .B2(_13638_),
    .X(_03011_));
 sky130_fd_sc_hd__buf_2 _17613_ (.A(_13627_),
    .X(_13639_));
 sky130_fd_sc_hd__buf_1 _17614_ (.A(_13639_),
    .X(_13640_));
 sky130_fd_sc_hd__buf_2 _17615_ (.A(_13630_),
    .X(_13641_));
 sky130_fd_sc_hd__buf_1 _17616_ (.A(_13641_),
    .X(_13642_));
 sky130_fd_sc_hd__a22o_1 _17617_ (.A1(\cpuregs[5][15] ),
    .A2(_13640_),
    .B1(_13220_),
    .B2(_13642_),
    .X(_03010_));
 sky130_fd_sc_hd__a22o_1 _17618_ (.A1(\cpuregs[5][14] ),
    .A2(_13640_),
    .B1(_13223_),
    .B2(_13642_),
    .X(_03009_));
 sky130_fd_sc_hd__a22o_1 _17619_ (.A1(\cpuregs[5][13] ),
    .A2(_13640_),
    .B1(_13224_),
    .B2(_13642_),
    .X(_03008_));
 sky130_fd_sc_hd__a22o_1 _17620_ (.A1(\cpuregs[5][12] ),
    .A2(_13640_),
    .B1(_13225_),
    .B2(_13642_),
    .X(_03007_));
 sky130_fd_sc_hd__buf_1 _17621_ (.A(_13639_),
    .X(_13643_));
 sky130_fd_sc_hd__buf_1 _17622_ (.A(_13641_),
    .X(_13644_));
 sky130_fd_sc_hd__a22o_1 _17623_ (.A1(\cpuregs[5][11] ),
    .A2(_13643_),
    .B1(_13227_),
    .B2(_13644_),
    .X(_03006_));
 sky130_fd_sc_hd__a22o_1 _17624_ (.A1(\cpuregs[5][10] ),
    .A2(_13643_),
    .B1(_13229_),
    .B2(_13644_),
    .X(_03005_));
 sky130_fd_sc_hd__a22o_1 _17625_ (.A1(\cpuregs[5][9] ),
    .A2(_13643_),
    .B1(_13230_),
    .B2(_13644_),
    .X(_03004_));
 sky130_fd_sc_hd__a22o_1 _17626_ (.A1(\cpuregs[5][8] ),
    .A2(_13643_),
    .B1(_13231_),
    .B2(_13644_),
    .X(_03003_));
 sky130_fd_sc_hd__buf_1 _17627_ (.A(_13639_),
    .X(_13645_));
 sky130_fd_sc_hd__buf_1 _17628_ (.A(_13641_),
    .X(_13646_));
 sky130_fd_sc_hd__a22o_1 _17629_ (.A1(\cpuregs[5][7] ),
    .A2(_13645_),
    .B1(_13233_),
    .B2(_13646_),
    .X(_03002_));
 sky130_fd_sc_hd__a22o_1 _17630_ (.A1(\cpuregs[5][6] ),
    .A2(_13645_),
    .B1(_13235_),
    .B2(_13646_),
    .X(_03001_));
 sky130_fd_sc_hd__a22o_1 _17631_ (.A1(\cpuregs[5][5] ),
    .A2(_13645_),
    .B1(_13236_),
    .B2(_13646_),
    .X(_03000_));
 sky130_fd_sc_hd__a22o_1 _17632_ (.A1(\cpuregs[5][4] ),
    .A2(_13645_),
    .B1(_13237_),
    .B2(_13646_),
    .X(_02999_));
 sky130_fd_sc_hd__buf_1 _17633_ (.A(_13639_),
    .X(_13647_));
 sky130_fd_sc_hd__buf_1 _17634_ (.A(_13641_),
    .X(_13648_));
 sky130_fd_sc_hd__a22o_1 _17635_ (.A1(\cpuregs[5][3] ),
    .A2(_13647_),
    .B1(_13239_),
    .B2(_13648_),
    .X(_02998_));
 sky130_fd_sc_hd__a22o_1 _17636_ (.A1(\cpuregs[5][2] ),
    .A2(_13647_),
    .B1(_13241_),
    .B2(_13648_),
    .X(_02997_));
 sky130_fd_sc_hd__a22o_1 _17637_ (.A1(\cpuregs[5][1] ),
    .A2(_13647_),
    .B1(_13242_),
    .B2(_13648_),
    .X(_02996_));
 sky130_fd_sc_hd__a22o_1 _17638_ (.A1(\cpuregs[5][0] ),
    .A2(_13647_),
    .B1(_13243_),
    .B2(_13648_),
    .X(_02995_));
 sky130_fd_sc_hd__or2_1 _17639_ (.A(_12561_),
    .B(_12567_),
    .X(_13649_));
 sky130_fd_sc_hd__buf_4 _17640_ (.A(_13649_),
    .X(_13650_));
 sky130_fd_sc_hd__buf_1 _17641_ (.A(_13650_),
    .X(_13651_));
 sky130_vsdinv _17642_ (.A(_13649_),
    .Y(_13652_));
 sky130_fd_sc_hd__buf_4 _17643_ (.A(_13652_),
    .X(_13653_));
 sky130_fd_sc_hd__buf_1 _17644_ (.A(_13653_),
    .X(_13654_));
 sky130_fd_sc_hd__a22o_1 _17645_ (.A1(\cpuregs[2][31] ),
    .A2(_13651_),
    .B1(_13193_),
    .B2(_13654_),
    .X(_02994_));
 sky130_fd_sc_hd__a22o_1 _17646_ (.A1(\cpuregs[2][30] ),
    .A2(_13651_),
    .B1(_13197_),
    .B2(_13654_),
    .X(_02993_));
 sky130_fd_sc_hd__a22o_1 _17647_ (.A1(\cpuregs[2][29] ),
    .A2(_13651_),
    .B1(_13198_),
    .B2(_13654_),
    .X(_02992_));
 sky130_fd_sc_hd__a22o_1 _17648_ (.A1(\cpuregs[2][28] ),
    .A2(_13651_),
    .B1(_13199_),
    .B2(_13654_),
    .X(_02991_));
 sky130_fd_sc_hd__buf_1 _17649_ (.A(_13650_),
    .X(_13655_));
 sky130_fd_sc_hd__buf_1 _17650_ (.A(_13653_),
    .X(_13656_));
 sky130_fd_sc_hd__a22o_1 _17651_ (.A1(\cpuregs[2][27] ),
    .A2(_13655_),
    .B1(_13201_),
    .B2(_13656_),
    .X(_02990_));
 sky130_fd_sc_hd__a22o_1 _17652_ (.A1(\cpuregs[2][26] ),
    .A2(_13655_),
    .B1(_13203_),
    .B2(_13656_),
    .X(_02989_));
 sky130_fd_sc_hd__a22o_1 _17653_ (.A1(\cpuregs[2][25] ),
    .A2(_13655_),
    .B1(_13204_),
    .B2(_13656_),
    .X(_02988_));
 sky130_fd_sc_hd__a22o_1 _17654_ (.A1(\cpuregs[2][24] ),
    .A2(_13655_),
    .B1(_13205_),
    .B2(_13656_),
    .X(_02987_));
 sky130_fd_sc_hd__buf_1 _17655_ (.A(_13650_),
    .X(_13657_));
 sky130_fd_sc_hd__buf_1 _17656_ (.A(_13653_),
    .X(_13658_));
 sky130_fd_sc_hd__a22o_1 _17657_ (.A1(\cpuregs[2][23] ),
    .A2(_13657_),
    .B1(_13207_),
    .B2(_13658_),
    .X(_02986_));
 sky130_fd_sc_hd__a22o_1 _17658_ (.A1(\cpuregs[2][22] ),
    .A2(_13657_),
    .B1(_13209_),
    .B2(_13658_),
    .X(_02985_));
 sky130_fd_sc_hd__a22o_1 _17659_ (.A1(\cpuregs[2][21] ),
    .A2(_13657_),
    .B1(_13210_),
    .B2(_13658_),
    .X(_02984_));
 sky130_fd_sc_hd__a22o_1 _17660_ (.A1(\cpuregs[2][20] ),
    .A2(_13657_),
    .B1(_13211_),
    .B2(_13658_),
    .X(_02983_));
 sky130_fd_sc_hd__buf_1 _17661_ (.A(_13650_),
    .X(_13659_));
 sky130_fd_sc_hd__buf_1 _17662_ (.A(_13653_),
    .X(_13660_));
 sky130_fd_sc_hd__a22o_1 _17663_ (.A1(\cpuregs[2][19] ),
    .A2(_13659_),
    .B1(_13213_),
    .B2(_13660_),
    .X(_02982_));
 sky130_fd_sc_hd__a22o_1 _17664_ (.A1(\cpuregs[2][18] ),
    .A2(_13659_),
    .B1(_13215_),
    .B2(_13660_),
    .X(_02981_));
 sky130_fd_sc_hd__a22o_1 _17665_ (.A1(\cpuregs[2][17] ),
    .A2(_13659_),
    .B1(_13216_),
    .B2(_13660_),
    .X(_02980_));
 sky130_fd_sc_hd__a22o_1 _17666_ (.A1(\cpuregs[2][16] ),
    .A2(_13659_),
    .B1(_13217_),
    .B2(_13660_),
    .X(_02979_));
 sky130_fd_sc_hd__clkbuf_4 _17667_ (.A(_13649_),
    .X(_13661_));
 sky130_fd_sc_hd__buf_1 _17668_ (.A(_13661_),
    .X(_13662_));
 sky130_fd_sc_hd__clkbuf_4 _17669_ (.A(_13652_),
    .X(_13663_));
 sky130_fd_sc_hd__buf_1 _17670_ (.A(_13663_),
    .X(_13664_));
 sky130_fd_sc_hd__a22o_1 _17671_ (.A1(\cpuregs[2][15] ),
    .A2(_13662_),
    .B1(_13220_),
    .B2(_13664_),
    .X(_02978_));
 sky130_fd_sc_hd__a22o_1 _17672_ (.A1(\cpuregs[2][14] ),
    .A2(_13662_),
    .B1(_13223_),
    .B2(_13664_),
    .X(_02977_));
 sky130_fd_sc_hd__a22o_1 _17673_ (.A1(\cpuregs[2][13] ),
    .A2(_13662_),
    .B1(_13224_),
    .B2(_13664_),
    .X(_02976_));
 sky130_fd_sc_hd__a22o_1 _17674_ (.A1(\cpuregs[2][12] ),
    .A2(_13662_),
    .B1(_13225_),
    .B2(_13664_),
    .X(_02975_));
 sky130_fd_sc_hd__buf_1 _17675_ (.A(_13661_),
    .X(_13665_));
 sky130_fd_sc_hd__buf_1 _17676_ (.A(_13663_),
    .X(_13666_));
 sky130_fd_sc_hd__a22o_1 _17677_ (.A1(\cpuregs[2][11] ),
    .A2(_13665_),
    .B1(_13227_),
    .B2(_13666_),
    .X(_02974_));
 sky130_fd_sc_hd__a22o_1 _17678_ (.A1(\cpuregs[2][10] ),
    .A2(_13665_),
    .B1(_13229_),
    .B2(_13666_),
    .X(_02973_));
 sky130_fd_sc_hd__a22o_1 _17679_ (.A1(\cpuregs[2][9] ),
    .A2(_13665_),
    .B1(_13230_),
    .B2(_13666_),
    .X(_02972_));
 sky130_fd_sc_hd__a22o_1 _17680_ (.A1(\cpuregs[2][8] ),
    .A2(_13665_),
    .B1(_13231_),
    .B2(_13666_),
    .X(_02971_));
 sky130_fd_sc_hd__buf_1 _17681_ (.A(_13661_),
    .X(_13667_));
 sky130_fd_sc_hd__buf_1 _17682_ (.A(_13663_),
    .X(_13668_));
 sky130_fd_sc_hd__a22o_1 _17683_ (.A1(\cpuregs[2][7] ),
    .A2(_13667_),
    .B1(_13233_),
    .B2(_13668_),
    .X(_02970_));
 sky130_fd_sc_hd__a22o_1 _17684_ (.A1(\cpuregs[2][6] ),
    .A2(_13667_),
    .B1(_13235_),
    .B2(_13668_),
    .X(_02969_));
 sky130_fd_sc_hd__a22o_1 _17685_ (.A1(\cpuregs[2][5] ),
    .A2(_13667_),
    .B1(_13236_),
    .B2(_13668_),
    .X(_02968_));
 sky130_fd_sc_hd__a22o_1 _17686_ (.A1(\cpuregs[2][4] ),
    .A2(_13667_),
    .B1(_13237_),
    .B2(_13668_),
    .X(_02967_));
 sky130_fd_sc_hd__buf_1 _17687_ (.A(_13661_),
    .X(_13669_));
 sky130_fd_sc_hd__buf_1 _17688_ (.A(_13663_),
    .X(_13670_));
 sky130_fd_sc_hd__a22o_1 _17689_ (.A1(\cpuregs[2][3] ),
    .A2(_13669_),
    .B1(_13239_),
    .B2(_13670_),
    .X(_02966_));
 sky130_fd_sc_hd__a22o_1 _17690_ (.A1(\cpuregs[2][2] ),
    .A2(_13669_),
    .B1(_13241_),
    .B2(_13670_),
    .X(_02965_));
 sky130_fd_sc_hd__a22o_1 _17691_ (.A1(\cpuregs[2][1] ),
    .A2(_13669_),
    .B1(_13242_),
    .B2(_13670_),
    .X(_02964_));
 sky130_fd_sc_hd__a22o_1 _17692_ (.A1(\cpuregs[2][0] ),
    .A2(_13669_),
    .B1(_13243_),
    .B2(_13670_),
    .X(_02963_));
 sky130_fd_sc_hd__buf_2 _17693_ (.A(_11547_),
    .X(_13671_));
 sky130_fd_sc_hd__clkbuf_2 _17694_ (.A(_13671_),
    .X(_13672_));
 sky130_fd_sc_hd__buf_8 _17695_ (.A(_13672_),
    .X(mem_xfer));
 sky130_fd_sc_hd__buf_1 _17696_ (.A(_11546_),
    .X(_13673_));
 sky130_fd_sc_hd__buf_1 _17697_ (.A(_13673_),
    .X(_13674_));
 sky130_fd_sc_hd__a22o_1 _17698_ (.A1(_11923_),
    .A2(_13674_),
    .B1(net57),
    .B2(net415),
    .X(_02962_));
 sky130_fd_sc_hd__a22o_1 _17699_ (.A1(_11924_),
    .A2(_13674_),
    .B1(net56),
    .B2(net415),
    .X(_02961_));
 sky130_fd_sc_hd__buf_1 _17700_ (.A(_13672_),
    .X(_13675_));
 sky130_fd_sc_hd__a22o_1 _17701_ (.A1(_13255_),
    .A2(_13674_),
    .B1(net54),
    .B2(_13675_),
    .X(_02960_));
 sky130_fd_sc_hd__a22o_1 _17702_ (.A1(_13294_),
    .A2(_13674_),
    .B1(net53),
    .B2(_13675_),
    .X(_02959_));
 sky130_fd_sc_hd__buf_1 _17703_ (.A(_13673_),
    .X(_13676_));
 sky130_fd_sc_hd__a22o_1 _17704_ (.A1(_13305_),
    .A2(_13676_),
    .B1(net52),
    .B2(_13675_),
    .X(_02958_));
 sky130_fd_sc_hd__a22o_1 _17705_ (.A1(_13295_),
    .A2(_13676_),
    .B1(net51),
    .B2(_13675_),
    .X(_02957_));
 sky130_fd_sc_hd__buf_1 _17706_ (.A(_13671_),
    .X(_13677_));
 sky130_fd_sc_hd__clkbuf_2 _17707_ (.A(_13677_),
    .X(_13678_));
 sky130_fd_sc_hd__a22o_1 _17708_ (.A1(_13330_),
    .A2(_13676_),
    .B1(net50),
    .B2(_13678_),
    .X(_02956_));
 sky130_fd_sc_hd__a22o_1 _17709_ (.A1(_13338_),
    .A2(_13676_),
    .B1(net49),
    .B2(_13678_),
    .X(_02955_));
 sky130_fd_sc_hd__buf_1 _17710_ (.A(_13673_),
    .X(_13679_));
 sky130_fd_sc_hd__a22o_1 _17711_ (.A1(\mem_rdata_q[23] ),
    .A2(_13679_),
    .B1(net48),
    .B2(_13678_),
    .X(_02954_));
 sky130_fd_sc_hd__a22o_1 _17712_ (.A1(\mem_rdata_q[22] ),
    .A2(_13679_),
    .B1(net47),
    .B2(_13678_),
    .X(_02953_));
 sky130_fd_sc_hd__buf_1 _17713_ (.A(_13677_),
    .X(_13680_));
 sky130_fd_sc_hd__a22o_1 _17714_ (.A1(_13315_),
    .A2(_13679_),
    .B1(net46),
    .B2(_13680_),
    .X(_02952_));
 sky130_fd_sc_hd__a22o_1 _17715_ (.A1(\mem_rdata_q[20] ),
    .A2(_13679_),
    .B1(net464),
    .B2(_13680_),
    .X(_02951_));
 sky130_fd_sc_hd__buf_1 _17716_ (.A(_13673_),
    .X(_13681_));
 sky130_fd_sc_hd__a22o_1 _17717_ (.A1(\mem_rdata_q[19] ),
    .A2(_13681_),
    .B1(net43),
    .B2(_13680_),
    .X(_02950_));
 sky130_fd_sc_hd__a22o_1 _17718_ (.A1(\mem_rdata_q[18] ),
    .A2(_13681_),
    .B1(net42),
    .B2(_13680_),
    .X(_02949_));
 sky130_fd_sc_hd__clkbuf_2 _17719_ (.A(_13677_),
    .X(_13682_));
 sky130_fd_sc_hd__a22o_1 _17720_ (.A1(\mem_rdata_q[17] ),
    .A2(_13681_),
    .B1(net41),
    .B2(_13682_),
    .X(_02948_));
 sky130_fd_sc_hd__a22o_1 _17721_ (.A1(\mem_rdata_q[16] ),
    .A2(_13681_),
    .B1(net40),
    .B2(_13682_),
    .X(_02947_));
 sky130_fd_sc_hd__buf_1 _17722_ (.A(_11546_),
    .X(_13683_));
 sky130_fd_sc_hd__clkbuf_2 _17723_ (.A(_13683_),
    .X(_13684_));
 sky130_fd_sc_hd__a22o_1 _17724_ (.A1(\mem_rdata_q[15] ),
    .A2(_13684_),
    .B1(net39),
    .B2(_13682_),
    .X(_02946_));
 sky130_fd_sc_hd__a22o_1 _17725_ (.A1(_11939_),
    .A2(_13684_),
    .B1(net38),
    .B2(_13682_),
    .X(_02945_));
 sky130_fd_sc_hd__buf_1 _17726_ (.A(_13677_),
    .X(_13685_));
 sky130_fd_sc_hd__a22o_1 _17727_ (.A1(_11947_),
    .A2(_13684_),
    .B1(net37),
    .B2(_13685_),
    .X(_02944_));
 sky130_fd_sc_hd__a22o_1 _17728_ (.A1(_11915_),
    .A2(_13684_),
    .B1(net36),
    .B2(_13685_),
    .X(_02943_));
 sky130_fd_sc_hd__buf_1 _17729_ (.A(_13683_),
    .X(_13686_));
 sky130_fd_sc_hd__a22o_1 _17730_ (.A1(\mem_rdata_q[11] ),
    .A2(_13686_),
    .B1(net35),
    .B2(_13685_),
    .X(_02942_));
 sky130_fd_sc_hd__a22o_1 _17731_ (.A1(\mem_rdata_q[10] ),
    .A2(_13686_),
    .B1(net34),
    .B2(_13685_),
    .X(_02941_));
 sky130_fd_sc_hd__buf_1 _17732_ (.A(_13671_),
    .X(_13687_));
 sky130_fd_sc_hd__a22o_1 _17733_ (.A1(\mem_rdata_q[9] ),
    .A2(_13686_),
    .B1(net64),
    .B2(_13687_),
    .X(_02940_));
 sky130_fd_sc_hd__a22o_1 _17734_ (.A1(\mem_rdata_q[8] ),
    .A2(_13686_),
    .B1(net63),
    .B2(_13687_),
    .X(_02939_));
 sky130_fd_sc_hd__buf_1 _17735_ (.A(_13683_),
    .X(_13688_));
 sky130_fd_sc_hd__a22o_1 _17736_ (.A1(\mem_rdata_q[7] ),
    .A2(_13688_),
    .B1(net62),
    .B2(_13687_),
    .X(_02938_));
 sky130_fd_sc_hd__a22o_1 _17737_ (.A1(\mem_rdata_q[6] ),
    .A2(_13688_),
    .B1(net61),
    .B2(_13687_),
    .X(_02937_));
 sky130_fd_sc_hd__buf_1 _17738_ (.A(_13671_),
    .X(_13689_));
 sky130_fd_sc_hd__a22o_1 _17739_ (.A1(\mem_rdata_q[5] ),
    .A2(_13688_),
    .B1(net60),
    .B2(_13689_),
    .X(_02936_));
 sky130_fd_sc_hd__a22o_1 _17740_ (.A1(\mem_rdata_q[4] ),
    .A2(_13688_),
    .B1(net59),
    .B2(_13689_),
    .X(_02935_));
 sky130_fd_sc_hd__buf_1 _17741_ (.A(_13683_),
    .X(_13690_));
 sky130_fd_sc_hd__a22o_1 _17742_ (.A1(\mem_rdata_q[3] ),
    .A2(_13690_),
    .B1(net58),
    .B2(_13689_),
    .X(_02934_));
 sky130_fd_sc_hd__a22o_1 _17743_ (.A1(\mem_rdata_q[2] ),
    .A2(_13690_),
    .B1(net55),
    .B2(_13689_),
    .X(_02933_));
 sky130_fd_sc_hd__a22o_1 _17744_ (.A1(\mem_rdata_q[1] ),
    .A2(_13690_),
    .B1(net44),
    .B2(_13672_),
    .X(_02932_));
 sky130_fd_sc_hd__a22o_1 _17745_ (.A1(\mem_rdata_q[0] ),
    .A2(_13690_),
    .B1(net33),
    .B2(_13672_),
    .X(_02931_));
 sky130_fd_sc_hd__or4_4 _17746_ (.A(_12769_),
    .B(_12554_),
    .C(_12553_),
    .D(_12566_),
    .X(_13691_));
 sky130_fd_sc_hd__clkbuf_4 _17747_ (.A(_13691_),
    .X(_13692_));
 sky130_fd_sc_hd__buf_1 _17748_ (.A(_13692_),
    .X(_13693_));
 sky130_vsdinv _17749_ (.A(_13691_),
    .Y(_13694_));
 sky130_fd_sc_hd__clkbuf_4 _17750_ (.A(_13694_),
    .X(_13695_));
 sky130_fd_sc_hd__buf_1 _17751_ (.A(_13695_),
    .X(_13696_));
 sky130_fd_sc_hd__a22o_1 _17752_ (.A1(\cpuregs[18][31] ),
    .A2(_13693_),
    .B1(_13193_),
    .B2(_13696_),
    .X(_02930_));
 sky130_fd_sc_hd__a22o_1 _17753_ (.A1(\cpuregs[18][30] ),
    .A2(_13693_),
    .B1(_13197_),
    .B2(_13696_),
    .X(_02929_));
 sky130_fd_sc_hd__a22o_1 _17754_ (.A1(\cpuregs[18][29] ),
    .A2(_13693_),
    .B1(_13198_),
    .B2(_13696_),
    .X(_02928_));
 sky130_fd_sc_hd__a22o_1 _17755_ (.A1(\cpuregs[18][28] ),
    .A2(_13693_),
    .B1(_13199_),
    .B2(_13696_),
    .X(_02927_));
 sky130_fd_sc_hd__clkbuf_2 _17756_ (.A(_13692_),
    .X(_13697_));
 sky130_fd_sc_hd__clkbuf_2 _17757_ (.A(_13695_),
    .X(_13698_));
 sky130_fd_sc_hd__a22o_1 _17758_ (.A1(\cpuregs[18][27] ),
    .A2(_13697_),
    .B1(_13201_),
    .B2(_13698_),
    .X(_02926_));
 sky130_fd_sc_hd__a22o_1 _17759_ (.A1(\cpuregs[18][26] ),
    .A2(_13697_),
    .B1(_13203_),
    .B2(_13698_),
    .X(_02925_));
 sky130_fd_sc_hd__a22o_1 _17760_ (.A1(\cpuregs[18][25] ),
    .A2(_13697_),
    .B1(_13204_),
    .B2(_13698_),
    .X(_02924_));
 sky130_fd_sc_hd__a22o_1 _17761_ (.A1(\cpuregs[18][24] ),
    .A2(_13697_),
    .B1(_13205_),
    .B2(_13698_),
    .X(_02923_));
 sky130_fd_sc_hd__buf_1 _17762_ (.A(_13692_),
    .X(_13699_));
 sky130_fd_sc_hd__buf_1 _17763_ (.A(_13695_),
    .X(_13700_));
 sky130_fd_sc_hd__a22o_1 _17764_ (.A1(\cpuregs[18][23] ),
    .A2(_13699_),
    .B1(_13207_),
    .B2(_13700_),
    .X(_02922_));
 sky130_fd_sc_hd__a22o_1 _17765_ (.A1(\cpuregs[18][22] ),
    .A2(_13699_),
    .B1(_13209_),
    .B2(_13700_),
    .X(_02921_));
 sky130_fd_sc_hd__a22o_1 _17766_ (.A1(\cpuregs[18][21] ),
    .A2(_13699_),
    .B1(_13210_),
    .B2(_13700_),
    .X(_02920_));
 sky130_fd_sc_hd__a22o_1 _17767_ (.A1(\cpuregs[18][20] ),
    .A2(_13699_),
    .B1(_13211_),
    .B2(_13700_),
    .X(_02919_));
 sky130_fd_sc_hd__buf_1 _17768_ (.A(_13692_),
    .X(_13701_));
 sky130_fd_sc_hd__buf_1 _17769_ (.A(_13695_),
    .X(_13702_));
 sky130_fd_sc_hd__a22o_1 _17770_ (.A1(\cpuregs[18][19] ),
    .A2(_13701_),
    .B1(_13213_),
    .B2(_13702_),
    .X(_02918_));
 sky130_fd_sc_hd__a22o_1 _17771_ (.A1(\cpuregs[18][18] ),
    .A2(_13701_),
    .B1(_13215_),
    .B2(_13702_),
    .X(_02917_));
 sky130_fd_sc_hd__a22o_1 _17772_ (.A1(\cpuregs[18][17] ),
    .A2(_13701_),
    .B1(_13216_),
    .B2(_13702_),
    .X(_02916_));
 sky130_fd_sc_hd__a22o_1 _17773_ (.A1(\cpuregs[18][16] ),
    .A2(_13701_),
    .B1(_13217_),
    .B2(_13702_),
    .X(_02915_));
 sky130_fd_sc_hd__buf_2 _17774_ (.A(_13691_),
    .X(_13703_));
 sky130_fd_sc_hd__buf_1 _17775_ (.A(_13703_),
    .X(_13704_));
 sky130_fd_sc_hd__clkbuf_4 _17776_ (.A(_13694_),
    .X(_13705_));
 sky130_fd_sc_hd__buf_1 _17777_ (.A(_13705_),
    .X(_13706_));
 sky130_fd_sc_hd__a22o_1 _17778_ (.A1(\cpuregs[18][15] ),
    .A2(_13704_),
    .B1(_13220_),
    .B2(_13706_),
    .X(_02914_));
 sky130_fd_sc_hd__a22o_1 _17779_ (.A1(\cpuregs[18][14] ),
    .A2(_13704_),
    .B1(_13223_),
    .B2(_13706_),
    .X(_02913_));
 sky130_fd_sc_hd__a22o_1 _17780_ (.A1(\cpuregs[18][13] ),
    .A2(_13704_),
    .B1(_13224_),
    .B2(_13706_),
    .X(_02912_));
 sky130_fd_sc_hd__a22o_1 _17781_ (.A1(\cpuregs[18][12] ),
    .A2(_13704_),
    .B1(_13225_),
    .B2(_13706_),
    .X(_02911_));
 sky130_fd_sc_hd__buf_1 _17782_ (.A(_13703_),
    .X(_13707_));
 sky130_fd_sc_hd__buf_1 _17783_ (.A(_13705_),
    .X(_13708_));
 sky130_fd_sc_hd__a22o_1 _17784_ (.A1(\cpuregs[18][11] ),
    .A2(_13707_),
    .B1(_13227_),
    .B2(_13708_),
    .X(_02910_));
 sky130_fd_sc_hd__a22o_1 _17785_ (.A1(\cpuregs[18][10] ),
    .A2(_13707_),
    .B1(_13229_),
    .B2(_13708_),
    .X(_02909_));
 sky130_fd_sc_hd__a22o_1 _17786_ (.A1(\cpuregs[18][9] ),
    .A2(_13707_),
    .B1(_13230_),
    .B2(_13708_),
    .X(_02908_));
 sky130_fd_sc_hd__a22o_1 _17787_ (.A1(\cpuregs[18][8] ),
    .A2(_13707_),
    .B1(_13231_),
    .B2(_13708_),
    .X(_02907_));
 sky130_fd_sc_hd__buf_1 _17788_ (.A(_13703_),
    .X(_13709_));
 sky130_fd_sc_hd__buf_1 _17789_ (.A(_13705_),
    .X(_13710_));
 sky130_fd_sc_hd__a22o_1 _17790_ (.A1(\cpuregs[18][7] ),
    .A2(_13709_),
    .B1(_13233_),
    .B2(_13710_),
    .X(_02906_));
 sky130_fd_sc_hd__a22o_1 _17791_ (.A1(\cpuregs[18][6] ),
    .A2(_13709_),
    .B1(_13235_),
    .B2(_13710_),
    .X(_02905_));
 sky130_fd_sc_hd__a22o_1 _17792_ (.A1(\cpuregs[18][5] ),
    .A2(_13709_),
    .B1(_13236_),
    .B2(_13710_),
    .X(_02904_));
 sky130_fd_sc_hd__a22o_1 _17793_ (.A1(\cpuregs[18][4] ),
    .A2(_13709_),
    .B1(_13237_),
    .B2(_13710_),
    .X(_02903_));
 sky130_fd_sc_hd__buf_1 _17794_ (.A(_13703_),
    .X(_13711_));
 sky130_fd_sc_hd__buf_1 _17795_ (.A(_13705_),
    .X(_13712_));
 sky130_fd_sc_hd__a22o_1 _17796_ (.A1(\cpuregs[18][3] ),
    .A2(_13711_),
    .B1(_13239_),
    .B2(_13712_),
    .X(_02902_));
 sky130_fd_sc_hd__a22o_1 _17797_ (.A1(\cpuregs[18][2] ),
    .A2(_13711_),
    .B1(_13241_),
    .B2(_13712_),
    .X(_02901_));
 sky130_fd_sc_hd__a22o_1 _17798_ (.A1(\cpuregs[18][1] ),
    .A2(_13711_),
    .B1(_13242_),
    .B2(_13712_),
    .X(_02900_));
 sky130_fd_sc_hd__a22o_1 _17799_ (.A1(\cpuregs[18][0] ),
    .A2(_13711_),
    .B1(_13243_),
    .B2(_13712_),
    .X(_02899_));
 sky130_fd_sc_hd__or2_2 _17800_ (.A(_12567_),
    .B(_12655_),
    .X(_13713_));
 sky130_fd_sc_hd__clkbuf_4 _17801_ (.A(_13713_),
    .X(_13714_));
 sky130_fd_sc_hd__buf_1 _17802_ (.A(_13714_),
    .X(_13715_));
 sky130_vsdinv _17803_ (.A(_13713_),
    .Y(_13716_));
 sky130_fd_sc_hd__clkbuf_4 _17804_ (.A(_13716_),
    .X(_13717_));
 sky130_fd_sc_hd__buf_1 _17805_ (.A(_13717_),
    .X(_13718_));
 sky130_fd_sc_hd__a22o_1 _17806_ (.A1(\cpuregs[10][31] ),
    .A2(_13715_),
    .B1(_12571_),
    .B2(_13718_),
    .X(_02898_));
 sky130_fd_sc_hd__a22o_1 _17807_ (.A1(\cpuregs[10][30] ),
    .A2(_13715_),
    .B1(_12576_),
    .B2(_13718_),
    .X(_02897_));
 sky130_fd_sc_hd__a22o_1 _17808_ (.A1(\cpuregs[10][29] ),
    .A2(_13715_),
    .B1(_12578_),
    .B2(_13718_),
    .X(_02896_));
 sky130_fd_sc_hd__a22o_1 _17809_ (.A1(\cpuregs[10][28] ),
    .A2(_13715_),
    .B1(_12580_),
    .B2(_13718_),
    .X(_02895_));
 sky130_fd_sc_hd__buf_1 _17810_ (.A(_13714_),
    .X(_13719_));
 sky130_fd_sc_hd__buf_1 _17811_ (.A(_13717_),
    .X(_13720_));
 sky130_fd_sc_hd__a22o_1 _17812_ (.A1(\cpuregs[10][27] ),
    .A2(_13719_),
    .B1(_12583_),
    .B2(_13720_),
    .X(_02894_));
 sky130_fd_sc_hd__a22o_1 _17813_ (.A1(\cpuregs[10][26] ),
    .A2(_13719_),
    .B1(_12586_),
    .B2(_13720_),
    .X(_02893_));
 sky130_fd_sc_hd__a22o_1 _17814_ (.A1(\cpuregs[10][25] ),
    .A2(_13719_),
    .B1(_12588_),
    .B2(_13720_),
    .X(_02892_));
 sky130_fd_sc_hd__a22o_1 _17815_ (.A1(\cpuregs[10][24] ),
    .A2(_13719_),
    .B1(_12590_),
    .B2(_13720_),
    .X(_02891_));
 sky130_fd_sc_hd__buf_1 _17816_ (.A(_13714_),
    .X(_13721_));
 sky130_fd_sc_hd__buf_1 _17817_ (.A(_13717_),
    .X(_13722_));
 sky130_fd_sc_hd__a22o_1 _17818_ (.A1(\cpuregs[10][23] ),
    .A2(_13721_),
    .B1(_12593_),
    .B2(_13722_),
    .X(_02890_));
 sky130_fd_sc_hd__a22o_1 _17819_ (.A1(\cpuregs[10][22] ),
    .A2(_13721_),
    .B1(_12596_),
    .B2(_13722_),
    .X(_02889_));
 sky130_fd_sc_hd__a22o_1 _17820_ (.A1(\cpuregs[10][21] ),
    .A2(_13721_),
    .B1(_12598_),
    .B2(_13722_),
    .X(_02888_));
 sky130_fd_sc_hd__a22o_1 _17821_ (.A1(\cpuregs[10][20] ),
    .A2(_13721_),
    .B1(_12600_),
    .B2(_13722_),
    .X(_02887_));
 sky130_fd_sc_hd__buf_1 _17822_ (.A(_13714_),
    .X(_13723_));
 sky130_fd_sc_hd__buf_1 _17823_ (.A(_13717_),
    .X(_13724_));
 sky130_fd_sc_hd__a22o_1 _17824_ (.A1(\cpuregs[10][19] ),
    .A2(_13723_),
    .B1(_12603_),
    .B2(_13724_),
    .X(_02886_));
 sky130_fd_sc_hd__a22o_1 _17825_ (.A1(\cpuregs[10][18] ),
    .A2(_13723_),
    .B1(_12606_),
    .B2(_13724_),
    .X(_02885_));
 sky130_fd_sc_hd__a22o_1 _17826_ (.A1(\cpuregs[10][17] ),
    .A2(_13723_),
    .B1(_12608_),
    .B2(_13724_),
    .X(_02884_));
 sky130_fd_sc_hd__a22o_1 _17827_ (.A1(\cpuregs[10][16] ),
    .A2(_13723_),
    .B1(_12610_),
    .B2(_13724_),
    .X(_02883_));
 sky130_fd_sc_hd__clkbuf_2 _17828_ (.A(_13713_),
    .X(_13725_));
 sky130_fd_sc_hd__buf_1 _17829_ (.A(_13725_),
    .X(_13726_));
 sky130_fd_sc_hd__clkbuf_2 _17830_ (.A(_13716_),
    .X(_13727_));
 sky130_fd_sc_hd__buf_1 _17831_ (.A(_13727_),
    .X(_13728_));
 sky130_fd_sc_hd__a22o_1 _17832_ (.A1(\cpuregs[10][15] ),
    .A2(_13726_),
    .B1(_12614_),
    .B2(_13728_),
    .X(_02882_));
 sky130_fd_sc_hd__a22o_1 _17833_ (.A1(\cpuregs[10][14] ),
    .A2(_13726_),
    .B1(_12618_),
    .B2(_13728_),
    .X(_02881_));
 sky130_fd_sc_hd__a22o_1 _17834_ (.A1(\cpuregs[10][13] ),
    .A2(_13726_),
    .B1(_12620_),
    .B2(_13728_),
    .X(_02880_));
 sky130_fd_sc_hd__a22o_1 _17835_ (.A1(\cpuregs[10][12] ),
    .A2(_13726_),
    .B1(_12622_),
    .B2(_13728_),
    .X(_02879_));
 sky130_fd_sc_hd__clkbuf_2 _17836_ (.A(_13725_),
    .X(_13729_));
 sky130_fd_sc_hd__clkbuf_2 _17837_ (.A(_13727_),
    .X(_13730_));
 sky130_fd_sc_hd__a22o_1 _17838_ (.A1(\cpuregs[10][11] ),
    .A2(_13729_),
    .B1(_12625_),
    .B2(_13730_),
    .X(_02878_));
 sky130_fd_sc_hd__a22o_1 _17839_ (.A1(\cpuregs[10][10] ),
    .A2(_13729_),
    .B1(_12628_),
    .B2(_13730_),
    .X(_02877_));
 sky130_fd_sc_hd__a22o_1 _17840_ (.A1(\cpuregs[10][9] ),
    .A2(_13729_),
    .B1(_12630_),
    .B2(_13730_),
    .X(_02876_));
 sky130_fd_sc_hd__a22o_1 _17841_ (.A1(\cpuregs[10][8] ),
    .A2(_13729_),
    .B1(_12632_),
    .B2(_13730_),
    .X(_02875_));
 sky130_fd_sc_hd__buf_1 _17842_ (.A(_13725_),
    .X(_13731_));
 sky130_fd_sc_hd__buf_1 _17843_ (.A(_13727_),
    .X(_13732_));
 sky130_fd_sc_hd__a22o_1 _17844_ (.A1(\cpuregs[10][7] ),
    .A2(_13731_),
    .B1(_12635_),
    .B2(_13732_),
    .X(_02874_));
 sky130_fd_sc_hd__a22o_1 _17845_ (.A1(\cpuregs[10][6] ),
    .A2(_13731_),
    .B1(_12638_),
    .B2(_13732_),
    .X(_02873_));
 sky130_fd_sc_hd__a22o_1 _17846_ (.A1(\cpuregs[10][5] ),
    .A2(_13731_),
    .B1(_12640_),
    .B2(_13732_),
    .X(_02872_));
 sky130_fd_sc_hd__a22o_1 _17847_ (.A1(\cpuregs[10][4] ),
    .A2(_13731_),
    .B1(_12642_),
    .B2(_13732_),
    .X(_02871_));
 sky130_fd_sc_hd__buf_1 _17848_ (.A(_13725_),
    .X(_13733_));
 sky130_fd_sc_hd__buf_1 _17849_ (.A(_13727_),
    .X(_13734_));
 sky130_fd_sc_hd__a22o_1 _17850_ (.A1(\cpuregs[10][3] ),
    .A2(_13733_),
    .B1(_12645_),
    .B2(_13734_),
    .X(_02870_));
 sky130_fd_sc_hd__a22o_1 _17851_ (.A1(\cpuregs[10][2] ),
    .A2(_13733_),
    .B1(_12648_),
    .B2(_13734_),
    .X(_02869_));
 sky130_fd_sc_hd__a22o_1 _17852_ (.A1(\cpuregs[10][1] ),
    .A2(_13733_),
    .B1(_12650_),
    .B2(_13734_),
    .X(_02868_));
 sky130_fd_sc_hd__a22o_1 _17853_ (.A1(\cpuregs[10][0] ),
    .A2(_13733_),
    .B1(_12652_),
    .B2(_13734_),
    .X(_02867_));
 sky130_fd_sc_hd__clkbuf_1 _17854_ (.A(\cpuregs[0][31] ),
    .X(_02866_));
 sky130_fd_sc_hd__clkbuf_1 _17855_ (.A(\cpuregs[0][30] ),
    .X(_02865_));
 sky130_fd_sc_hd__clkbuf_1 _17856_ (.A(\cpuregs[0][29] ),
    .X(_02864_));
 sky130_fd_sc_hd__clkbuf_1 _17857_ (.A(\cpuregs[0][28] ),
    .X(_02863_));
 sky130_fd_sc_hd__clkbuf_1 _17858_ (.A(\cpuregs[0][27] ),
    .X(_02862_));
 sky130_fd_sc_hd__clkbuf_1 _17859_ (.A(\cpuregs[0][26] ),
    .X(_02861_));
 sky130_fd_sc_hd__clkbuf_1 _17860_ (.A(\cpuregs[0][25] ),
    .X(_02860_));
 sky130_fd_sc_hd__clkbuf_1 _17861_ (.A(\cpuregs[0][24] ),
    .X(_02859_));
 sky130_fd_sc_hd__clkbuf_1 _17862_ (.A(\cpuregs[0][23] ),
    .X(_02858_));
 sky130_fd_sc_hd__clkbuf_1 _17863_ (.A(\cpuregs[0][22] ),
    .X(_02857_));
 sky130_fd_sc_hd__clkbuf_1 _17864_ (.A(\cpuregs[0][21] ),
    .X(_02856_));
 sky130_fd_sc_hd__clkbuf_1 _17865_ (.A(\cpuregs[0][20] ),
    .X(_02855_));
 sky130_fd_sc_hd__clkbuf_1 _17866_ (.A(\cpuregs[0][19] ),
    .X(_02854_));
 sky130_fd_sc_hd__clkbuf_1 _17867_ (.A(\cpuregs[0][18] ),
    .X(_02853_));
 sky130_fd_sc_hd__clkbuf_1 _17868_ (.A(\cpuregs[0][17] ),
    .X(_02852_));
 sky130_fd_sc_hd__clkbuf_1 _17869_ (.A(\cpuregs[0][16] ),
    .X(_02851_));
 sky130_fd_sc_hd__clkbuf_1 _17870_ (.A(\cpuregs[0][15] ),
    .X(_02850_));
 sky130_fd_sc_hd__clkbuf_1 _17871_ (.A(\cpuregs[0][14] ),
    .X(_02849_));
 sky130_fd_sc_hd__clkbuf_1 _17872_ (.A(\cpuregs[0][13] ),
    .X(_02848_));
 sky130_fd_sc_hd__clkbuf_1 _17873_ (.A(\cpuregs[0][12] ),
    .X(_02847_));
 sky130_fd_sc_hd__clkbuf_1 _17874_ (.A(\cpuregs[0][11] ),
    .X(_02846_));
 sky130_fd_sc_hd__clkbuf_1 _17875_ (.A(\cpuregs[0][10] ),
    .X(_02845_));
 sky130_fd_sc_hd__clkbuf_1 _17876_ (.A(\cpuregs[0][9] ),
    .X(_02844_));
 sky130_fd_sc_hd__clkbuf_1 _17877_ (.A(\cpuregs[0][8] ),
    .X(_02843_));
 sky130_fd_sc_hd__clkbuf_1 _17878_ (.A(\cpuregs[0][7] ),
    .X(_02842_));
 sky130_fd_sc_hd__clkbuf_1 _17879_ (.A(\cpuregs[0][6] ),
    .X(_02841_));
 sky130_fd_sc_hd__clkbuf_1 _17880_ (.A(\cpuregs[0][5] ),
    .X(_02840_));
 sky130_fd_sc_hd__clkbuf_1 _17881_ (.A(\cpuregs[0][4] ),
    .X(_02839_));
 sky130_fd_sc_hd__clkbuf_1 _17882_ (.A(\cpuregs[0][3] ),
    .X(_02838_));
 sky130_fd_sc_hd__clkbuf_1 _17883_ (.A(\cpuregs[0][2] ),
    .X(_02837_));
 sky130_fd_sc_hd__clkbuf_1 _17884_ (.A(\cpuregs[0][1] ),
    .X(_02836_));
 sky130_fd_sc_hd__clkbuf_1 _17885_ (.A(\cpuregs[0][0] ),
    .X(_02835_));
 sky130_fd_sc_hd__or2_2 _17886_ (.A(_12567_),
    .B(_12876_),
    .X(_13735_));
 sky130_fd_sc_hd__clkbuf_4 _17887_ (.A(_13735_),
    .X(_13736_));
 sky130_fd_sc_hd__buf_1 _17888_ (.A(_13736_),
    .X(_13737_));
 sky130_vsdinv _17889_ (.A(_13735_),
    .Y(_13738_));
 sky130_fd_sc_hd__clkbuf_4 _17890_ (.A(_13738_),
    .X(_13739_));
 sky130_fd_sc_hd__buf_1 _17891_ (.A(_13739_),
    .X(_13740_));
 sky130_fd_sc_hd__a22o_1 _17892_ (.A1(\cpuregs[14][31] ),
    .A2(_13737_),
    .B1(_12571_),
    .B2(_13740_),
    .X(_02834_));
 sky130_fd_sc_hd__a22o_1 _17893_ (.A1(\cpuregs[14][30] ),
    .A2(_13737_),
    .B1(_12576_),
    .B2(_13740_),
    .X(_02833_));
 sky130_fd_sc_hd__a22o_1 _17894_ (.A1(\cpuregs[14][29] ),
    .A2(_13737_),
    .B1(_12578_),
    .B2(_13740_),
    .X(_02832_));
 sky130_fd_sc_hd__a22o_1 _17895_ (.A1(\cpuregs[14][28] ),
    .A2(_13737_),
    .B1(_12580_),
    .B2(_13740_),
    .X(_02831_));
 sky130_fd_sc_hd__buf_1 _17896_ (.A(_13736_),
    .X(_13741_));
 sky130_fd_sc_hd__buf_1 _17897_ (.A(_13739_),
    .X(_13742_));
 sky130_fd_sc_hd__a22o_1 _17898_ (.A1(\cpuregs[14][27] ),
    .A2(_13741_),
    .B1(_12583_),
    .B2(_13742_),
    .X(_02830_));
 sky130_fd_sc_hd__a22o_1 _17899_ (.A1(\cpuregs[14][26] ),
    .A2(_13741_),
    .B1(_12586_),
    .B2(_13742_),
    .X(_02829_));
 sky130_fd_sc_hd__a22o_1 _17900_ (.A1(\cpuregs[14][25] ),
    .A2(_13741_),
    .B1(_12588_),
    .B2(_13742_),
    .X(_02828_));
 sky130_fd_sc_hd__a22o_1 _17901_ (.A1(\cpuregs[14][24] ),
    .A2(_13741_),
    .B1(_12590_),
    .B2(_13742_),
    .X(_02827_));
 sky130_fd_sc_hd__buf_1 _17902_ (.A(_13736_),
    .X(_13743_));
 sky130_fd_sc_hd__buf_1 _17903_ (.A(_13739_),
    .X(_13744_));
 sky130_fd_sc_hd__a22o_1 _17904_ (.A1(\cpuregs[14][23] ),
    .A2(_13743_),
    .B1(_12593_),
    .B2(_13744_),
    .X(_02826_));
 sky130_fd_sc_hd__a22o_1 _17905_ (.A1(\cpuregs[14][22] ),
    .A2(_13743_),
    .B1(_12596_),
    .B2(_13744_),
    .X(_02825_));
 sky130_fd_sc_hd__a22o_1 _17906_ (.A1(\cpuregs[14][21] ),
    .A2(_13743_),
    .B1(_12598_),
    .B2(_13744_),
    .X(_02824_));
 sky130_fd_sc_hd__a22o_1 _17907_ (.A1(\cpuregs[14][20] ),
    .A2(_13743_),
    .B1(_12600_),
    .B2(_13744_),
    .X(_02823_));
 sky130_fd_sc_hd__buf_1 _17908_ (.A(_13736_),
    .X(_13745_));
 sky130_fd_sc_hd__buf_1 _17909_ (.A(_13739_),
    .X(_13746_));
 sky130_fd_sc_hd__a22o_1 _17910_ (.A1(\cpuregs[14][19] ),
    .A2(_13745_),
    .B1(_12603_),
    .B2(_13746_),
    .X(_02822_));
 sky130_fd_sc_hd__a22o_1 _17911_ (.A1(\cpuregs[14][18] ),
    .A2(_13745_),
    .B1(_12606_),
    .B2(_13746_),
    .X(_02821_));
 sky130_fd_sc_hd__a22o_1 _17912_ (.A1(\cpuregs[14][17] ),
    .A2(_13745_),
    .B1(_12608_),
    .B2(_13746_),
    .X(_02820_));
 sky130_fd_sc_hd__a22o_1 _17913_ (.A1(\cpuregs[14][16] ),
    .A2(_13745_),
    .B1(_12610_),
    .B2(_13746_),
    .X(_02819_));
 sky130_fd_sc_hd__buf_2 _17914_ (.A(_13735_),
    .X(_13747_));
 sky130_fd_sc_hd__buf_1 _17915_ (.A(_13747_),
    .X(_13748_));
 sky130_fd_sc_hd__buf_2 _17916_ (.A(_13738_),
    .X(_13749_));
 sky130_fd_sc_hd__buf_1 _17917_ (.A(_13749_),
    .X(_13750_));
 sky130_fd_sc_hd__a22o_1 _17918_ (.A1(\cpuregs[14][15] ),
    .A2(_13748_),
    .B1(_12614_),
    .B2(_13750_),
    .X(_02818_));
 sky130_fd_sc_hd__a22o_1 _17919_ (.A1(\cpuregs[14][14] ),
    .A2(_13748_),
    .B1(_12618_),
    .B2(_13750_),
    .X(_02817_));
 sky130_fd_sc_hd__a22o_1 _17920_ (.A1(\cpuregs[14][13] ),
    .A2(_13748_),
    .B1(_12620_),
    .B2(_13750_),
    .X(_02816_));
 sky130_fd_sc_hd__a22o_1 _17921_ (.A1(\cpuregs[14][12] ),
    .A2(_13748_),
    .B1(_12622_),
    .B2(_13750_),
    .X(_02815_));
 sky130_fd_sc_hd__buf_1 _17922_ (.A(_13747_),
    .X(_13751_));
 sky130_fd_sc_hd__buf_1 _17923_ (.A(_13749_),
    .X(_13752_));
 sky130_fd_sc_hd__a22o_1 _17924_ (.A1(\cpuregs[14][11] ),
    .A2(_13751_),
    .B1(_12625_),
    .B2(_13752_),
    .X(_02814_));
 sky130_fd_sc_hd__a22o_1 _17925_ (.A1(\cpuregs[14][10] ),
    .A2(_13751_),
    .B1(_12628_),
    .B2(_13752_),
    .X(_02813_));
 sky130_fd_sc_hd__a22o_1 _17926_ (.A1(\cpuregs[14][9] ),
    .A2(_13751_),
    .B1(_12630_),
    .B2(_13752_),
    .X(_02812_));
 sky130_fd_sc_hd__a22o_1 _17927_ (.A1(\cpuregs[14][8] ),
    .A2(_13751_),
    .B1(_12632_),
    .B2(_13752_),
    .X(_02811_));
 sky130_fd_sc_hd__buf_1 _17928_ (.A(_13747_),
    .X(_13753_));
 sky130_fd_sc_hd__buf_1 _17929_ (.A(_13749_),
    .X(_13754_));
 sky130_fd_sc_hd__a22o_1 _17930_ (.A1(\cpuregs[14][7] ),
    .A2(_13753_),
    .B1(_12635_),
    .B2(_13754_),
    .X(_02810_));
 sky130_fd_sc_hd__a22o_1 _17931_ (.A1(\cpuregs[14][6] ),
    .A2(_13753_),
    .B1(_12638_),
    .B2(_13754_),
    .X(_02809_));
 sky130_fd_sc_hd__a22o_1 _17932_ (.A1(\cpuregs[14][5] ),
    .A2(_13753_),
    .B1(_12640_),
    .B2(_13754_),
    .X(_02808_));
 sky130_fd_sc_hd__a22o_1 _17933_ (.A1(\cpuregs[14][4] ),
    .A2(_13753_),
    .B1(_12642_),
    .B2(_13754_),
    .X(_02807_));
 sky130_fd_sc_hd__buf_1 _17934_ (.A(_13747_),
    .X(_13755_));
 sky130_fd_sc_hd__buf_1 _17935_ (.A(_13749_),
    .X(_13756_));
 sky130_fd_sc_hd__a22o_1 _17936_ (.A1(\cpuregs[14][3] ),
    .A2(_13755_),
    .B1(_12645_),
    .B2(_13756_),
    .X(_02806_));
 sky130_fd_sc_hd__a22o_1 _17937_ (.A1(\cpuregs[14][2] ),
    .A2(_13755_),
    .B1(_12648_),
    .B2(_13756_),
    .X(_02805_));
 sky130_fd_sc_hd__a22o_1 _17938_ (.A1(\cpuregs[14][1] ),
    .A2(_13755_),
    .B1(_12650_),
    .B2(_13756_),
    .X(_02804_));
 sky130_fd_sc_hd__a22o_1 _17939_ (.A1(\cpuregs[14][0] ),
    .A2(_13755_),
    .B1(_12652_),
    .B2(_13756_),
    .X(_02803_));
 sky130_fd_sc_hd__or2_2 _17940_ (.A(_12655_),
    .B(_12746_),
    .X(_13757_));
 sky130_fd_sc_hd__clkbuf_4 _17941_ (.A(_13757_),
    .X(_13758_));
 sky130_fd_sc_hd__buf_1 _17942_ (.A(_13758_),
    .X(_13759_));
 sky130_vsdinv _17943_ (.A(_13757_),
    .Y(_13760_));
 sky130_fd_sc_hd__clkbuf_4 _17944_ (.A(_13760_),
    .X(_13761_));
 sky130_fd_sc_hd__buf_1 _17945_ (.A(_13761_),
    .X(_13762_));
 sky130_fd_sc_hd__a22o_1 _17946_ (.A1(\cpuregs[8][31] ),
    .A2(_13759_),
    .B1(_12571_),
    .B2(_13762_),
    .X(_02802_));
 sky130_fd_sc_hd__a22o_1 _17947_ (.A1(\cpuregs[8][30] ),
    .A2(_13759_),
    .B1(_12576_),
    .B2(_13762_),
    .X(_02801_));
 sky130_fd_sc_hd__a22o_1 _17948_ (.A1(\cpuregs[8][29] ),
    .A2(_13759_),
    .B1(_12578_),
    .B2(_13762_),
    .X(_02800_));
 sky130_fd_sc_hd__a22o_1 _17949_ (.A1(\cpuregs[8][28] ),
    .A2(_13759_),
    .B1(_12580_),
    .B2(_13762_),
    .X(_02799_));
 sky130_fd_sc_hd__buf_1 _17950_ (.A(_13758_),
    .X(_13763_));
 sky130_fd_sc_hd__buf_1 _17951_ (.A(_13761_),
    .X(_13764_));
 sky130_fd_sc_hd__a22o_1 _17952_ (.A1(\cpuregs[8][27] ),
    .A2(_13763_),
    .B1(_12583_),
    .B2(_13764_),
    .X(_02798_));
 sky130_fd_sc_hd__a22o_1 _17953_ (.A1(\cpuregs[8][26] ),
    .A2(_13763_),
    .B1(_12586_),
    .B2(_13764_),
    .X(_02797_));
 sky130_fd_sc_hd__a22o_1 _17954_ (.A1(\cpuregs[8][25] ),
    .A2(_13763_),
    .B1(_12588_),
    .B2(_13764_),
    .X(_02796_));
 sky130_fd_sc_hd__a22o_1 _17955_ (.A1(\cpuregs[8][24] ),
    .A2(_13763_),
    .B1(_12590_),
    .B2(_13764_),
    .X(_02795_));
 sky130_fd_sc_hd__buf_1 _17956_ (.A(_13758_),
    .X(_13765_));
 sky130_fd_sc_hd__buf_1 _17957_ (.A(_13761_),
    .X(_13766_));
 sky130_fd_sc_hd__a22o_1 _17958_ (.A1(\cpuregs[8][23] ),
    .A2(_13765_),
    .B1(_12593_),
    .B2(_13766_),
    .X(_02794_));
 sky130_fd_sc_hd__a22o_1 _17959_ (.A1(\cpuregs[8][22] ),
    .A2(_13765_),
    .B1(_12596_),
    .B2(_13766_),
    .X(_02793_));
 sky130_fd_sc_hd__a22o_1 _17960_ (.A1(\cpuregs[8][21] ),
    .A2(_13765_),
    .B1(_12598_),
    .B2(_13766_),
    .X(_02792_));
 sky130_fd_sc_hd__a22o_1 _17961_ (.A1(\cpuregs[8][20] ),
    .A2(_13765_),
    .B1(_12600_),
    .B2(_13766_),
    .X(_02791_));
 sky130_fd_sc_hd__buf_1 _17962_ (.A(_13758_),
    .X(_13767_));
 sky130_fd_sc_hd__buf_1 _17963_ (.A(_13761_),
    .X(_13768_));
 sky130_fd_sc_hd__a22o_1 _17964_ (.A1(\cpuregs[8][19] ),
    .A2(_13767_),
    .B1(_12603_),
    .B2(_13768_),
    .X(_02790_));
 sky130_fd_sc_hd__a22o_1 _17965_ (.A1(\cpuregs[8][18] ),
    .A2(_13767_),
    .B1(_12606_),
    .B2(_13768_),
    .X(_02789_));
 sky130_fd_sc_hd__a22o_1 _17966_ (.A1(\cpuregs[8][17] ),
    .A2(_13767_),
    .B1(_12608_),
    .B2(_13768_),
    .X(_02788_));
 sky130_fd_sc_hd__a22o_1 _17967_ (.A1(\cpuregs[8][16] ),
    .A2(_13767_),
    .B1(_12610_),
    .B2(_13768_),
    .X(_02787_));
 sky130_fd_sc_hd__clkbuf_2 _17968_ (.A(_13757_),
    .X(_13769_));
 sky130_fd_sc_hd__buf_1 _17969_ (.A(_13769_),
    .X(_13770_));
 sky130_fd_sc_hd__clkbuf_2 _17970_ (.A(_13760_),
    .X(_13771_));
 sky130_fd_sc_hd__buf_1 _17971_ (.A(_13771_),
    .X(_13772_));
 sky130_fd_sc_hd__a22o_1 _17972_ (.A1(\cpuregs[8][15] ),
    .A2(_13770_),
    .B1(_12614_),
    .B2(_13772_),
    .X(_02786_));
 sky130_fd_sc_hd__a22o_1 _17973_ (.A1(\cpuregs[8][14] ),
    .A2(_13770_),
    .B1(_12618_),
    .B2(_13772_),
    .X(_02785_));
 sky130_fd_sc_hd__a22o_1 _17974_ (.A1(\cpuregs[8][13] ),
    .A2(_13770_),
    .B1(_12620_),
    .B2(_13772_),
    .X(_02784_));
 sky130_fd_sc_hd__a22o_1 _17975_ (.A1(\cpuregs[8][12] ),
    .A2(_13770_),
    .B1(_12622_),
    .B2(_13772_),
    .X(_02783_));
 sky130_fd_sc_hd__buf_1 _17976_ (.A(_13769_),
    .X(_13773_));
 sky130_fd_sc_hd__buf_1 _17977_ (.A(_13771_),
    .X(_13774_));
 sky130_fd_sc_hd__a22o_1 _17978_ (.A1(\cpuregs[8][11] ),
    .A2(_13773_),
    .B1(_12625_),
    .B2(_13774_),
    .X(_02782_));
 sky130_fd_sc_hd__a22o_1 _17979_ (.A1(\cpuregs[8][10] ),
    .A2(_13773_),
    .B1(_12628_),
    .B2(_13774_),
    .X(_02781_));
 sky130_fd_sc_hd__a22o_1 _17980_ (.A1(\cpuregs[8][9] ),
    .A2(_13773_),
    .B1(_12630_),
    .B2(_13774_),
    .X(_02780_));
 sky130_fd_sc_hd__a22o_1 _17981_ (.A1(\cpuregs[8][8] ),
    .A2(_13773_),
    .B1(_12632_),
    .B2(_13774_),
    .X(_02779_));
 sky130_fd_sc_hd__buf_1 _17982_ (.A(_13769_),
    .X(_13775_));
 sky130_fd_sc_hd__buf_1 _17983_ (.A(_13771_),
    .X(_13776_));
 sky130_fd_sc_hd__a22o_1 _17984_ (.A1(\cpuregs[8][7] ),
    .A2(_13775_),
    .B1(_12635_),
    .B2(_13776_),
    .X(_02778_));
 sky130_fd_sc_hd__a22o_1 _17985_ (.A1(\cpuregs[8][6] ),
    .A2(_13775_),
    .B1(_12638_),
    .B2(_13776_),
    .X(_02777_));
 sky130_fd_sc_hd__a22o_1 _17986_ (.A1(\cpuregs[8][5] ),
    .A2(_13775_),
    .B1(_12640_),
    .B2(_13776_),
    .X(_02776_));
 sky130_fd_sc_hd__a22o_1 _17987_ (.A1(\cpuregs[8][4] ),
    .A2(_13775_),
    .B1(_12642_),
    .B2(_13776_),
    .X(_02775_));
 sky130_fd_sc_hd__buf_1 _17988_ (.A(_13769_),
    .X(_13777_));
 sky130_fd_sc_hd__buf_1 _17989_ (.A(_13771_),
    .X(_13778_));
 sky130_fd_sc_hd__a22o_1 _17990_ (.A1(\cpuregs[8][3] ),
    .A2(_13777_),
    .B1(_12645_),
    .B2(_13778_),
    .X(_02774_));
 sky130_fd_sc_hd__a22o_1 _17991_ (.A1(\cpuregs[8][2] ),
    .A2(_13777_),
    .B1(_12648_),
    .B2(_13778_),
    .X(_02773_));
 sky130_fd_sc_hd__a22o_1 _17992_ (.A1(\cpuregs[8][1] ),
    .A2(_13777_),
    .B1(_12650_),
    .B2(_13778_),
    .X(_02772_));
 sky130_fd_sc_hd__a22o_1 _17993_ (.A1(\cpuregs[8][0] ),
    .A2(_13777_),
    .B1(_12652_),
    .B2(_13778_),
    .X(_02771_));
 sky130_fd_sc_hd__buf_4 _17994_ (.A(_11575_),
    .X(_13779_));
 sky130_fd_sc_hd__nor2_8 _17995_ (.A(_13779_),
    .B(_11784_),
    .Y(_00292_));
 sky130_fd_sc_hd__o21ai_1 _17996_ (.A1(_12558_),
    .A2(latched_store),
    .B1(_12016_),
    .Y(_13780_));
 sky130_fd_sc_hd__clkbuf_2 _17997_ (.A(\reg_next_pc[0] ),
    .X(_13781_));
 sky130_fd_sc_hd__o211a_1 _17998_ (.A1(net425),
    .A2(_13780_),
    .B1(_12396_),
    .C1(_13781_),
    .X(_02770_));
 sky130_fd_sc_hd__and2_1 _17999_ (.A(_12406_),
    .B(_00008_),
    .X(_02769_));
 sky130_fd_sc_hd__and2_1 _18000_ (.A(_12406_),
    .B(_14321_),
    .X(_02768_));
 sky130_fd_sc_hd__buf_1 _18001_ (.A(_12405_),
    .X(_13782_));
 sky130_fd_sc_hd__and2_1 _18002_ (.A(_13782_),
    .B(_00031_),
    .X(_02767_));
 sky130_fd_sc_hd__and2_1 _18003_ (.A(_13782_),
    .B(_00032_),
    .X(_02766_));
 sky130_fd_sc_hd__and2_1 _18004_ (.A(_13782_),
    .B(_00033_),
    .X(_02765_));
 sky130_fd_sc_hd__and2_1 _18005_ (.A(_13782_),
    .B(_00034_),
    .X(_02764_));
 sky130_fd_sc_hd__buf_1 _18006_ (.A(_12405_),
    .X(_13783_));
 sky130_fd_sc_hd__and2_1 _18007_ (.A(_13783_),
    .B(_00035_),
    .X(_02763_));
 sky130_fd_sc_hd__and2_1 _18008_ (.A(_13783_),
    .B(_00036_),
    .X(_02762_));
 sky130_fd_sc_hd__and2_1 _18009_ (.A(_13783_),
    .B(_00037_),
    .X(_02761_));
 sky130_fd_sc_hd__and2_1 _18010_ (.A(_13783_),
    .B(_00009_),
    .X(_02760_));
 sky130_fd_sc_hd__buf_1 _18011_ (.A(_12405_),
    .X(_13784_));
 sky130_fd_sc_hd__and2_1 _18012_ (.A(_13784_),
    .B(_00010_),
    .X(_02759_));
 sky130_fd_sc_hd__and2_1 _18013_ (.A(_13784_),
    .B(_00011_),
    .X(_02758_));
 sky130_fd_sc_hd__and2_1 _18014_ (.A(_13784_),
    .B(_00012_),
    .X(_02757_));
 sky130_fd_sc_hd__and2_1 _18015_ (.A(_13784_),
    .B(_00013_),
    .X(_02756_));
 sky130_fd_sc_hd__clkbuf_2 _18016_ (.A(_12395_),
    .X(_13785_));
 sky130_fd_sc_hd__buf_1 _18017_ (.A(_13785_),
    .X(_13786_));
 sky130_fd_sc_hd__and2_1 _18018_ (.A(_13786_),
    .B(_00014_),
    .X(_02755_));
 sky130_fd_sc_hd__and2_1 _18019_ (.A(_13786_),
    .B(_00015_),
    .X(_02754_));
 sky130_fd_sc_hd__and2_1 _18020_ (.A(_13786_),
    .B(_00016_),
    .X(_02753_));
 sky130_fd_sc_hd__and2_1 _18021_ (.A(_13786_),
    .B(_00017_),
    .X(_02752_));
 sky130_fd_sc_hd__buf_1 _18022_ (.A(_13785_),
    .X(_13787_));
 sky130_fd_sc_hd__and2_1 _18023_ (.A(_13787_),
    .B(_00018_),
    .X(_02751_));
 sky130_fd_sc_hd__and2_1 _18024_ (.A(_13787_),
    .B(_00019_),
    .X(_02750_));
 sky130_fd_sc_hd__and2_1 _18025_ (.A(_13787_),
    .B(_00020_),
    .X(_02749_));
 sky130_fd_sc_hd__and2_1 _18026_ (.A(_13787_),
    .B(_00021_),
    .X(_02748_));
 sky130_fd_sc_hd__clkbuf_2 _18027_ (.A(_13785_),
    .X(_13788_));
 sky130_fd_sc_hd__and2_1 _18028_ (.A(_13788_),
    .B(_00022_),
    .X(_02747_));
 sky130_fd_sc_hd__and2_1 _18029_ (.A(_13788_),
    .B(_00023_),
    .X(_02746_));
 sky130_fd_sc_hd__and2_1 _18030_ (.A(_13788_),
    .B(_00024_),
    .X(_02745_));
 sky130_fd_sc_hd__and2_1 _18031_ (.A(_13788_),
    .B(_00025_),
    .X(_02744_));
 sky130_fd_sc_hd__buf_1 _18032_ (.A(_13785_),
    .X(_13789_));
 sky130_fd_sc_hd__and2_1 _18033_ (.A(_13789_),
    .B(_00026_),
    .X(_02743_));
 sky130_fd_sc_hd__and2_1 _18034_ (.A(_13789_),
    .B(_00027_),
    .X(_02742_));
 sky130_fd_sc_hd__and2_1 _18035_ (.A(_13789_),
    .B(_00028_),
    .X(_02741_));
 sky130_fd_sc_hd__and2_1 _18036_ (.A(_13789_),
    .B(_00029_),
    .X(_02740_));
 sky130_fd_sc_hd__and2_1 _18037_ (.A(_11566_),
    .B(_00030_),
    .X(_02739_));
 sky130_vsdinv _18038_ (.A(\decoded_imm[1] ),
    .Y(_13790_));
 sky130_vsdinv _18039_ (.A(\mem_rdata_q[8] ),
    .Y(_13791_));
 sky130_fd_sc_hd__nor2_4 _18040_ (.A(_11891_),
    .B(is_sb_sh_sw),
    .Y(_13792_));
 sky130_fd_sc_hd__buf_1 _18041_ (.A(_13792_),
    .X(_13793_));
 sky130_vsdinv _18042_ (.A(\decoded_imm_uj[1] ),
    .Y(_13794_));
 sky130_fd_sc_hd__or2_1 _18043_ (.A(_13794_),
    .B(_13370_),
    .X(_13795_));
 sky130_fd_sc_hd__o221a_1 _18044_ (.A1(_13791_),
    .A2(_13793_),
    .B1(_13325_),
    .B2(_13285_),
    .C1(_13795_),
    .X(_13796_));
 sky130_fd_sc_hd__o22ai_1 _18045_ (.A1(_13790_),
    .A2(_13346_),
    .B1(_13254_),
    .B2(_13796_),
    .Y(_02738_));
 sky130_vsdinv _18046_ (.A(\decoded_imm[2] ),
    .Y(_13797_));
 sky130_fd_sc_hd__buf_1 _18047_ (.A(_13247_),
    .X(_13798_));
 sky130_vsdinv _18048_ (.A(\mem_rdata_q[9] ),
    .Y(_13799_));
 sky130_vsdinv _18049_ (.A(\mem_rdata_q[22] ),
    .Y(_13800_));
 sky130_vsdinv _18050_ (.A(\decoded_imm_uj[2] ),
    .Y(_13801_));
 sky130_fd_sc_hd__buf_1 _18051_ (.A(_13369_),
    .X(_13802_));
 sky130_fd_sc_hd__or2_1 _18052_ (.A(_13801_),
    .B(_13802_),
    .X(_13803_));
 sky130_fd_sc_hd__o221a_1 _18053_ (.A1(_13799_),
    .A2(_13793_),
    .B1(_13800_),
    .B2(_13285_),
    .C1(_13803_),
    .X(_13804_));
 sky130_fd_sc_hd__o22ai_1 _18054_ (.A1(_13797_),
    .A2(_13346_),
    .B1(_13798_),
    .B2(_13804_),
    .Y(_02737_));
 sky130_vsdinv _18055_ (.A(\decoded_imm[3] ),
    .Y(_13805_));
 sky130_vsdinv _18056_ (.A(\mem_rdata_q[10] ),
    .Y(_13806_));
 sky130_vsdinv _18057_ (.A(\mem_rdata_q[23] ),
    .Y(_13807_));
 sky130_vsdinv _18058_ (.A(\decoded_imm_uj[3] ),
    .Y(_13808_));
 sky130_fd_sc_hd__or2_1 _18059_ (.A(_13808_),
    .B(_13802_),
    .X(_13809_));
 sky130_fd_sc_hd__o221a_1 _18060_ (.A1(_13806_),
    .A2(_13793_),
    .B1(_13807_),
    .B2(_13285_),
    .C1(_13809_),
    .X(_13810_));
 sky130_fd_sc_hd__o22ai_1 _18061_ (.A1(_13805_),
    .A2(_13346_),
    .B1(_13798_),
    .B2(_13810_),
    .Y(_02736_));
 sky130_vsdinv _18062_ (.A(\decoded_imm[4] ),
    .Y(_13811_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _18063_ (.A(_13811_),
    .X(_13812_));
 sky130_fd_sc_hd__buf_1 _18064_ (.A(_11999_),
    .X(_13813_));
 sky130_vsdinv _18065_ (.A(\mem_rdata_q[11] ),
    .Y(_13814_));
 sky130_vsdinv _18066_ (.A(_13338_),
    .Y(_13815_));
 sky130_fd_sc_hd__inv_2 _18067_ (.A(\decoded_imm_uj[4] ),
    .Y(_00367_));
 sky130_fd_sc_hd__or2_1 _18068_ (.A(_00367_),
    .B(_13802_),
    .X(_13816_));
 sky130_fd_sc_hd__o221a_1 _18069_ (.A1(_13814_),
    .A2(_13793_),
    .B1(_13815_),
    .B2(_13284_),
    .C1(_13816_),
    .X(_13817_));
 sky130_fd_sc_hd__o22ai_1 _18070_ (.A1(_13812_),
    .A2(_13813_),
    .B1(_13798_),
    .B2(_13817_),
    .Y(_02735_));
 sky130_vsdinv _18071_ (.A(\decoded_imm[5] ),
    .Y(_13818_));
 sky130_vsdinv _18072_ (.A(\decoded_imm_uj[5] ),
    .Y(_13819_));
 sky130_fd_sc_hd__or3_4 _18073_ (.A(is_sb_sh_sw),
    .B(_13283_),
    .C(_11891_),
    .X(_13820_));
 sky130_vsdinv _18074_ (.A(_13820_),
    .Y(_13821_));
 sky130_fd_sc_hd__buf_1 _18075_ (.A(_13821_),
    .X(_13822_));
 sky130_fd_sc_hd__o22a_1 _18076_ (.A1(_13819_),
    .A2(_00323_),
    .B1(_13296_),
    .B2(_13822_),
    .X(_13823_));
 sky130_fd_sc_hd__o22ai_1 _18077_ (.A1(_13818_),
    .A2(_13813_),
    .B1(_13798_),
    .B2(_13823_),
    .Y(_02734_));
 sky130_vsdinv _18078_ (.A(\decoded_imm[6] ),
    .Y(_13824_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _18079_ (.A(_13824_),
    .X(_13825_));
 sky130_fd_sc_hd__clkbuf_2 _18080_ (.A(_13253_),
    .X(_13826_));
 sky130_fd_sc_hd__o2bb2a_1 _18081_ (.A1_N(_13272_),
    .A2_N(instr_jal),
    .B1(_13304_),
    .B2(_13821_),
    .X(_13827_));
 sky130_fd_sc_hd__o22ai_1 _18082_ (.A1(_13825_),
    .A2(_13813_),
    .B1(_13826_),
    .B2(_13827_),
    .Y(_02733_));
 sky130_vsdinv _18083_ (.A(\decoded_imm[7] ),
    .Y(_13828_));
 sky130_vsdinv _18084_ (.A(\decoded_imm_uj[7] ),
    .Y(_13829_));
 sky130_fd_sc_hd__o22a_1 _18085_ (.A1(_13829_),
    .A2(_00323_),
    .B1(_13287_),
    .B2(_13822_),
    .X(_13830_));
 sky130_fd_sc_hd__o22ai_1 _18086_ (.A1(_13828_),
    .A2(_13813_),
    .B1(_13826_),
    .B2(_13830_),
    .Y(_02732_));
 sky130_vsdinv _18087_ (.A(\decoded_imm[8] ),
    .Y(_13831_));
 sky130_fd_sc_hd__clkbuf_2 _18088_ (.A(_13831_),
    .X(_13832_));
 sky130_fd_sc_hd__clkbuf_2 _18089_ (.A(_13832_),
    .X(_13833_));
 sky130_fd_sc_hd__clkbuf_2 _18090_ (.A(_11999_),
    .X(_13834_));
 sky130_vsdinv _18091_ (.A(\decoded_imm_uj[8] ),
    .Y(_13835_));
 sky130_fd_sc_hd__buf_1 _18092_ (.A(_13370_),
    .X(_13836_));
 sky130_vsdinv _18093_ (.A(_13294_),
    .Y(_13837_));
 sky130_fd_sc_hd__o22a_1 _18094_ (.A1(_13835_),
    .A2(_13836_),
    .B1(_13837_),
    .B2(_13822_),
    .X(_13838_));
 sky130_fd_sc_hd__o22ai_1 _18095_ (.A1(_13833_),
    .A2(_13834_),
    .B1(_13826_),
    .B2(_13838_),
    .Y(_02731_));
 sky130_vsdinv _18096_ (.A(\decoded_imm[9] ),
    .Y(_13839_));
 sky130_vsdinv _18097_ (.A(\decoded_imm_uj[9] ),
    .Y(_13840_));
 sky130_vsdinv _18098_ (.A(_13255_),
    .Y(_13841_));
 sky130_fd_sc_hd__o22a_1 _18099_ (.A1(_13840_),
    .A2(_13836_),
    .B1(_13841_),
    .B2(_13822_),
    .X(_13842_));
 sky130_fd_sc_hd__o22ai_2 _18100_ (.A1(_13839_),
    .A2(_13834_),
    .B1(_13826_),
    .B2(_13842_),
    .Y(_02730_));
 sky130_vsdinv _18101_ (.A(\decoded_imm[10] ),
    .Y(_13843_));
 sky130_fd_sc_hd__clkbuf_2 _18102_ (.A(_13843_),
    .X(_13844_));
 sky130_fd_sc_hd__buf_1 _18103_ (.A(_13253_),
    .X(_13845_));
 sky130_vsdinv _18104_ (.A(\decoded_imm_uj[10] ),
    .Y(_13846_));
 sky130_fd_sc_hd__o22a_1 _18105_ (.A1(_13846_),
    .A2(_13836_),
    .B1(_11926_),
    .B2(_13821_),
    .X(_13847_));
 sky130_fd_sc_hd__o22ai_1 _18106_ (.A1(_13844_),
    .A2(_13834_),
    .B1(_13845_),
    .B2(_13847_),
    .Y(_02729_));
 sky130_vsdinv _18107_ (.A(\decoded_imm[11] ),
    .Y(_13848_));
 sky130_fd_sc_hd__clkbuf_2 _18108_ (.A(_13848_),
    .X(_13849_));
 sky130_vsdinv _18109_ (.A(\decoded_imm_uj[11] ),
    .Y(_13850_));
 sky130_fd_sc_hd__clkbuf_2 _18110_ (.A(_13802_),
    .X(_13851_));
 sky130_fd_sc_hd__o21ai_1 _18111_ (.A1(_13353_),
    .A2(_13283_),
    .B1(_11923_),
    .Y(_13852_));
 sky130_fd_sc_hd__o221a_2 _18112_ (.A1(_13850_),
    .A2(_13851_),
    .B1(_11992_),
    .B2(_13281_),
    .C1(_13852_),
    .X(_13853_));
 sky130_fd_sc_hd__o22ai_1 _18113_ (.A1(_13849_),
    .A2(_13834_),
    .B1(_13845_),
    .B2(_13853_),
    .Y(_02728_));
 sky130_vsdinv _18114_ (.A(\decoded_imm[12] ),
    .Y(_13854_));
 sky130_fd_sc_hd__clkbuf_2 _18115_ (.A(_13854_),
    .X(_13855_));
 sky130_fd_sc_hd__buf_1 _18116_ (.A(_13301_),
    .X(_13856_));
 sky130_vsdinv _18117_ (.A(\decoded_imm_uj[12] ),
    .Y(_13857_));
 sky130_vsdinv _18118_ (.A(_11755_),
    .Y(_13858_));
 sky130_fd_sc_hd__clkbuf_2 _18119_ (.A(_13858_),
    .X(_13859_));
 sky130_fd_sc_hd__or2_2 _18120_ (.A(_13328_),
    .B(_13821_),
    .X(_13860_));
 sky130_fd_sc_hd__buf_1 _18121_ (.A(_13860_),
    .X(_13861_));
 sky130_fd_sc_hd__o221a_1 _18122_ (.A1(_13857_),
    .A2(_13851_),
    .B1(_11905_),
    .B2(_13859_),
    .C1(_13861_),
    .X(_13862_));
 sky130_fd_sc_hd__o22ai_1 _18123_ (.A1(_13855_),
    .A2(_13856_),
    .B1(_13845_),
    .B2(_13862_),
    .Y(_02727_));
 sky130_vsdinv _18124_ (.A(\decoded_imm[13] ),
    .Y(_13863_));
 sky130_fd_sc_hd__clkbuf_2 _18125_ (.A(_13863_),
    .X(_13864_));
 sky130_vsdinv _18126_ (.A(\decoded_imm_uj[13] ),
    .Y(_13865_));
 sky130_fd_sc_hd__clkbuf_2 _18127_ (.A(_13858_),
    .X(_13866_));
 sky130_fd_sc_hd__o221a_1 _18128_ (.A1(_13865_),
    .A2(_13851_),
    .B1(_11903_),
    .B2(_13866_),
    .C1(_13861_),
    .X(_13867_));
 sky130_fd_sc_hd__o22ai_1 _18129_ (.A1(_13864_),
    .A2(_13856_),
    .B1(_13845_),
    .B2(_13867_),
    .Y(_02726_));
 sky130_vsdinv _18130_ (.A(\decoded_imm[14] ),
    .Y(_13868_));
 sky130_fd_sc_hd__clkbuf_2 _18131_ (.A(_13868_),
    .X(_13869_));
 sky130_fd_sc_hd__buf_1 _18132_ (.A(_13253_),
    .X(_13870_));
 sky130_vsdinv _18133_ (.A(\decoded_imm_uj[14] ),
    .Y(_13871_));
 sky130_fd_sc_hd__o221a_1 _18134_ (.A1(_13871_),
    .A2(_13851_),
    .B1(_00334_),
    .B2(_13866_),
    .C1(_13861_),
    .X(_13872_));
 sky130_fd_sc_hd__o22ai_1 _18135_ (.A1(_13869_),
    .A2(_13856_),
    .B1(_13870_),
    .B2(_13872_),
    .Y(_02725_));
 sky130_vsdinv _18136_ (.A(\decoded_imm[15] ),
    .Y(_13873_));
 sky130_fd_sc_hd__clkbuf_2 _18137_ (.A(_13873_),
    .X(_13874_));
 sky130_vsdinv _18138_ (.A(\decoded_imm_uj[15] ),
    .Y(_13875_));
 sky130_fd_sc_hd__buf_1 _18139_ (.A(_13369_),
    .X(_13876_));
 sky130_vsdinv _18140_ (.A(\mem_rdata_q[15] ),
    .Y(_13877_));
 sky130_fd_sc_hd__o221a_1 _18141_ (.A1(_13875_),
    .A2(_13876_),
    .B1(_13877_),
    .B2(_13866_),
    .C1(_13861_),
    .X(_13878_));
 sky130_fd_sc_hd__o22ai_1 _18142_ (.A1(_13874_),
    .A2(_13856_),
    .B1(_13870_),
    .B2(_13878_),
    .Y(_02724_));
 sky130_vsdinv _18143_ (.A(\decoded_imm[16] ),
    .Y(_13879_));
 sky130_fd_sc_hd__clkbuf_2 _18144_ (.A(_13879_),
    .X(_13880_));
 sky130_fd_sc_hd__buf_2 _18145_ (.A(_13880_),
    .X(_13881_));
 sky130_fd_sc_hd__buf_1 _18146_ (.A(_13301_),
    .X(_13882_));
 sky130_vsdinv _18147_ (.A(\decoded_imm_uj[16] ),
    .Y(_13883_));
 sky130_vsdinv _18148_ (.A(\mem_rdata_q[16] ),
    .Y(_13884_));
 sky130_fd_sc_hd__buf_1 _18149_ (.A(_13860_),
    .X(_13885_));
 sky130_fd_sc_hd__o221a_1 _18150_ (.A1(_13883_),
    .A2(_13876_),
    .B1(_13884_),
    .B2(_13866_),
    .C1(_13885_),
    .X(_13886_));
 sky130_fd_sc_hd__o22ai_1 _18151_ (.A1(_13881_),
    .A2(_13882_),
    .B1(_13870_),
    .B2(_13886_),
    .Y(_02723_));
 sky130_vsdinv _18152_ (.A(\decoded_imm[17] ),
    .Y(_13887_));
 sky130_vsdinv _18153_ (.A(\decoded_imm_uj[17] ),
    .Y(_13888_));
 sky130_vsdinv _18154_ (.A(\mem_rdata_q[17] ),
    .Y(_13889_));
 sky130_fd_sc_hd__clkbuf_2 _18155_ (.A(_13858_),
    .X(_13890_));
 sky130_fd_sc_hd__o221a_1 _18156_ (.A1(_13888_),
    .A2(_13876_),
    .B1(_13889_),
    .B2(_13890_),
    .C1(_13885_),
    .X(_13891_));
 sky130_fd_sc_hd__o22ai_1 _18157_ (.A1(_13887_),
    .A2(_13882_),
    .B1(_13870_),
    .B2(_13891_),
    .Y(_02722_));
 sky130_vsdinv _18158_ (.A(\decoded_imm[18] ),
    .Y(_13892_));
 sky130_fd_sc_hd__clkbuf_2 _18159_ (.A(_13892_),
    .X(_13893_));
 sky130_vsdinv _18160_ (.A(\decoded_imm_uj[18] ),
    .Y(_13894_));
 sky130_vsdinv _18161_ (.A(\mem_rdata_q[18] ),
    .Y(_13895_));
 sky130_fd_sc_hd__o221a_1 _18162_ (.A1(_13894_),
    .A2(_13876_),
    .B1(_13895_),
    .B2(_13890_),
    .C1(_13885_),
    .X(_13896_));
 sky130_fd_sc_hd__o22ai_1 _18163_ (.A1(_13893_),
    .A2(_13882_),
    .B1(_12389_),
    .B2(_13896_),
    .Y(_02721_));
 sky130_vsdinv _18164_ (.A(\decoded_imm[19] ),
    .Y(_13897_));
 sky130_fd_sc_hd__clkbuf_2 _18165_ (.A(_13897_),
    .X(_13898_));
 sky130_vsdinv _18166_ (.A(\decoded_imm_uj[19] ),
    .Y(_13899_));
 sky130_vsdinv _18167_ (.A(\mem_rdata_q[19] ),
    .Y(_13900_));
 sky130_fd_sc_hd__o221a_1 _18168_ (.A1(_13899_),
    .A2(_13370_),
    .B1(_13900_),
    .B2(_13890_),
    .C1(_13885_),
    .X(_13901_));
 sky130_fd_sc_hd__o22ai_1 _18169_ (.A1(_13898_),
    .A2(_13882_),
    .B1(_12389_),
    .B2(_13901_),
    .Y(_02720_));
 sky130_fd_sc_hd__nor2_4 _18170_ (.A(_13339_),
    .B(_13284_),
    .Y(_13902_));
 sky130_fd_sc_hd__buf_1 _18171_ (.A(_13902_),
    .X(_13903_));
 sky130_fd_sc_hd__buf_1 _18172_ (.A(_13903_),
    .X(_13904_));
 sky130_fd_sc_hd__clkbuf_2 _18173_ (.A(_13890_),
    .X(_13905_));
 sky130_fd_sc_hd__o21ai_2 _18174_ (.A1(_13282_),
    .A2(_13905_),
    .B1(_13362_),
    .Y(_13906_));
 sky130_vsdinv _18175_ (.A(\decoded_imm_uj[20] ),
    .Y(_13907_));
 sky130_fd_sc_hd__buf_1 _18176_ (.A(_13907_),
    .X(_13908_));
 sky130_fd_sc_hd__buf_1 _18177_ (.A(_13908_),
    .X(_13909_));
 sky130_fd_sc_hd__buf_1 _18178_ (.A(_13909_),
    .X(_13910_));
 sky130_fd_sc_hd__buf_1 _18179_ (.A(_13910_),
    .X(_13911_));
 sky130_fd_sc_hd__buf_2 _18180_ (.A(_13911_),
    .X(_13912_));
 sky130_fd_sc_hd__o22ai_4 _18181_ (.A1(_13912_),
    .A2(_13369_),
    .B1(_13339_),
    .B2(_13792_),
    .Y(_13913_));
 sky130_fd_sc_hd__buf_1 _18182_ (.A(_13913_),
    .X(_13914_));
 sky130_fd_sc_hd__buf_1 _18183_ (.A(_13914_),
    .X(_13915_));
 sky130_fd_sc_hd__o32a_1 _18184_ (.A1(_13904_),
    .A2(_13906_),
    .A3(_13915_),
    .B1(\decoded_imm[20] ),
    .B2(_13250_),
    .X(_02719_));
 sky130_fd_sc_hd__o21ai_2 _18185_ (.A1(_13325_),
    .A2(_13905_),
    .B1(_13362_),
    .Y(_13916_));
 sky130_fd_sc_hd__buf_1 _18186_ (.A(_13249_),
    .X(_13917_));
 sky130_fd_sc_hd__o32a_1 _18187_ (.A1(_13904_),
    .A2(_13916_),
    .A3(_13915_),
    .B1(\decoded_imm[21] ),
    .B2(_13917_),
    .X(_02718_));
 sky130_fd_sc_hd__buf_1 _18188_ (.A(_13354_),
    .X(_13918_));
 sky130_fd_sc_hd__o21ai_1 _18189_ (.A1(_13800_),
    .A2(_13905_),
    .B1(_13918_),
    .Y(_13919_));
 sky130_fd_sc_hd__o32a_1 _18190_ (.A1(_13904_),
    .A2(_13919_),
    .A3(_13915_),
    .B1(\decoded_imm[22] ),
    .B2(_13917_),
    .X(_02717_));
 sky130_fd_sc_hd__o21ai_1 _18191_ (.A1(_13807_),
    .A2(_13905_),
    .B1(_13918_),
    .Y(_13920_));
 sky130_fd_sc_hd__o32a_1 _18192_ (.A1(_13904_),
    .A2(_13920_),
    .A3(_13915_),
    .B1(\decoded_imm[23] ),
    .B2(_13917_),
    .X(_02716_));
 sky130_fd_sc_hd__buf_1 _18193_ (.A(_13902_),
    .X(_13921_));
 sky130_fd_sc_hd__buf_1 _18194_ (.A(_13858_),
    .X(_13922_));
 sky130_fd_sc_hd__o21ai_1 _18195_ (.A1(_13815_),
    .A2(_13922_),
    .B1(_13918_),
    .Y(_13923_));
 sky130_fd_sc_hd__buf_1 _18196_ (.A(_13913_),
    .X(_13924_));
 sky130_fd_sc_hd__buf_2 _18197_ (.A(\decoded_imm[24] ),
    .X(_13925_));
 sky130_fd_sc_hd__o32a_1 _18198_ (.A1(_13921_),
    .A2(_13923_),
    .A3(_13924_),
    .B1(_13925_),
    .B2(_13917_),
    .X(_02715_));
 sky130_fd_sc_hd__o21ai_1 _18199_ (.A1(_13296_),
    .A2(_13922_),
    .B1(_13918_),
    .Y(_13926_));
 sky130_fd_sc_hd__buf_2 _18200_ (.A(\decoded_imm[25] ),
    .X(_13927_));
 sky130_fd_sc_hd__buf_1 _18201_ (.A(_13249_),
    .X(_13928_));
 sky130_fd_sc_hd__o32a_1 _18202_ (.A1(_13921_),
    .A2(_13926_),
    .A3(_13924_),
    .B1(_13927_),
    .B2(_13928_),
    .X(_02714_));
 sky130_fd_sc_hd__buf_1 _18203_ (.A(_13354_),
    .X(_13929_));
 sky130_fd_sc_hd__o21ai_1 _18204_ (.A1(_13304_),
    .A2(_13922_),
    .B1(_13929_),
    .Y(_13930_));
 sky130_fd_sc_hd__buf_2 _18205_ (.A(\decoded_imm[26] ),
    .X(_13931_));
 sky130_fd_sc_hd__o32a_1 _18206_ (.A1(_13921_),
    .A2(_13930_),
    .A3(_13924_),
    .B1(_13931_),
    .B2(_13928_),
    .X(_02713_));
 sky130_fd_sc_hd__o21ai_1 _18207_ (.A1(_13287_),
    .A2(_13922_),
    .B1(_13929_),
    .Y(_13932_));
 sky130_fd_sc_hd__buf_2 _18208_ (.A(\decoded_imm[27] ),
    .X(_13933_));
 sky130_fd_sc_hd__o32a_1 _18209_ (.A1(_13921_),
    .A2(_13932_),
    .A3(_13924_),
    .B1(_13933_),
    .B2(_13928_),
    .X(_02712_));
 sky130_fd_sc_hd__o21ai_1 _18210_ (.A1(_13837_),
    .A2(_13859_),
    .B1(_13929_),
    .Y(_13934_));
 sky130_fd_sc_hd__buf_2 _18211_ (.A(\decoded_imm[28] ),
    .X(_13935_));
 sky130_fd_sc_hd__o32a_1 _18212_ (.A1(_13903_),
    .A2(_13934_),
    .A3(_13914_),
    .B1(_13935_),
    .B2(_13928_),
    .X(_02711_));
 sky130_fd_sc_hd__o21ai_1 _18213_ (.A1(_13841_),
    .A2(_13859_),
    .B1(_13929_),
    .Y(_13936_));
 sky130_fd_sc_hd__buf_2 _18214_ (.A(\decoded_imm[29] ),
    .X(_13937_));
 sky130_fd_sc_hd__o32a_1 _18215_ (.A1(_13903_),
    .A2(_13936_),
    .A3(_13914_),
    .B1(_13937_),
    .B2(_13280_),
    .X(_02710_));
 sky130_fd_sc_hd__o21ai_1 _18216_ (.A1(_11926_),
    .A2(_13859_),
    .B1(_11932_),
    .Y(_13938_));
 sky130_fd_sc_hd__o32a_1 _18217_ (.A1(_13903_),
    .A2(_13938_),
    .A3(_13914_),
    .B1(\decoded_imm[30] ),
    .B2(_13280_),
    .X(_02709_));
 sky130_vsdinv _18218_ (.A(\decoded_imm[31] ),
    .Y(_13939_));
 sky130_fd_sc_hd__buf_2 _18219_ (.A(_13939_),
    .X(_13940_));
 sky130_fd_sc_hd__buf_2 _18220_ (.A(_13912_),
    .X(_13941_));
 sky130_fd_sc_hd__nor2_1 _18221_ (.A(_11755_),
    .B(_13820_),
    .Y(_13942_));
 sky130_fd_sc_hd__o22a_1 _18222_ (.A1(_13941_),
    .A2(_13836_),
    .B1(_13339_),
    .B2(_13942_),
    .X(_13943_));
 sky130_fd_sc_hd__o22ai_1 _18223_ (.A1(_13940_),
    .A2(_13376_),
    .B1(_12389_),
    .B2(_13943_),
    .Y(_02708_));
 sky130_fd_sc_hd__or2_1 _18224_ (.A(\cpu_state[4] ),
    .B(_11735_),
    .X(_13944_));
 sky130_fd_sc_hd__buf_4 _18225_ (.A(_13944_),
    .X(_02542_));
 sky130_vsdinv _18226_ (.A(_02542_),
    .Y(_13945_));
 sky130_fd_sc_hd__or4_4 _18227_ (.A(_11586_),
    .B(_00331_),
    .C(_12874_),
    .D(_11739_),
    .X(_13946_));
 sky130_vsdinv _18228_ (.A(_13946_),
    .Y(_13947_));
 sky130_fd_sc_hd__buf_1 _18229_ (.A(_13946_),
    .X(_13948_));
 sky130_fd_sc_hd__a32o_1 _18230_ (.A1(_14281_),
    .A2(_13945_),
    .A3(_13947_),
    .B1(_12557_),
    .B2(_13948_),
    .X(_02707_));
 sky130_fd_sc_hd__clkbuf_4 _18231_ (.A(_11672_),
    .X(_00308_));
 sky130_fd_sc_hd__nor2_2 _18232_ (.A(net410),
    .B(_02542_),
    .Y(_13949_));
 sky130_fd_sc_hd__a32o_1 _18233_ (.A1(\decoded_rd[1] ),
    .A2(_13947_),
    .A3(_13949_),
    .B1(_12564_),
    .B2(_13948_),
    .X(_02706_));
 sky130_fd_sc_hd__a32o_1 _18234_ (.A1(\decoded_rd[2] ),
    .A2(_13947_),
    .A3(_13949_),
    .B1(_12770_),
    .B2(_13948_),
    .X(_02705_));
 sky130_fd_sc_hd__a32o_2 _18235_ (.A1(\decoded_rd[3] ),
    .A2(_13947_),
    .A3(_13949_),
    .B1(_12771_),
    .B2(_13948_),
    .X(_02704_));
 sky130_fd_sc_hd__or3_4 _18236_ (.A(_13353_),
    .B(_12362_),
    .C(_00310_),
    .X(_13950_));
 sky130_fd_sc_hd__o31ai_4 _18237_ (.A1(is_jalr_addi_slti_sltiu_xori_ori_andi),
    .A2(is_slli_srli_srai),
    .A3(is_lui_auipc_jal),
    .B1(_12274_),
    .Y(_13951_));
 sky130_fd_sc_hd__a21oi_1 _18238_ (.A1(_13950_),
    .A2(_13951_),
    .B1(_12682_),
    .Y(_02703_));
 sky130_vsdinv _18239_ (.A(_12734_),
    .Y(_13952_));
 sky130_fd_sc_hd__buf_1 _18240_ (.A(_13952_),
    .X(_13953_));
 sky130_fd_sc_hd__buf_1 _18241_ (.A(_13953_),
    .X(_13954_));
 sky130_fd_sc_hd__clkbuf_2 _18242_ (.A(_13954_),
    .X(_02327_));
 sky130_fd_sc_hd__and2_1 _18243_ (.A(_02327_),
    .B(_02558_),
    .X(_02702_));
 sky130_fd_sc_hd__buf_1 _18244_ (.A(_13954_),
    .X(_13955_));
 sky130_fd_sc_hd__and2_1 _18245_ (.A(_13955_),
    .B(_02557_),
    .X(_02701_));
 sky130_fd_sc_hd__and2_1 _18246_ (.A(_13955_),
    .B(_02556_),
    .X(_02700_));
 sky130_fd_sc_hd__and2_1 _18247_ (.A(_13955_),
    .B(_02555_),
    .X(_02699_));
 sky130_fd_sc_hd__and2_1 _18248_ (.A(_13955_),
    .B(_02554_),
    .X(_02698_));
 sky130_fd_sc_hd__buf_1 _18249_ (.A(_13953_),
    .X(_13956_));
 sky130_fd_sc_hd__and2_1 _18250_ (.A(_13956_),
    .B(_02553_),
    .X(_02697_));
 sky130_fd_sc_hd__and2_1 _18251_ (.A(_13956_),
    .B(_02552_),
    .X(_02696_));
 sky130_fd_sc_hd__and2_1 _18252_ (.A(_13956_),
    .B(_02551_),
    .X(_02695_));
 sky130_vsdinv _18253_ (.A(_12737_),
    .Y(_13957_));
 sky130_fd_sc_hd__buf_1 _18254_ (.A(_13957_),
    .X(_13958_));
 sky130_fd_sc_hd__clkbuf_2 _18255_ (.A(_13958_),
    .X(_02324_));
 sky130_fd_sc_hd__and2_1 _18256_ (.A(_02324_),
    .B(_00122_),
    .X(_02550_));
 sky130_fd_sc_hd__buf_1 _18257_ (.A(_13958_),
    .X(_13959_));
 sky130_fd_sc_hd__and3_1 _18258_ (.A(_13959_),
    .B(_00122_),
    .C(_13956_),
    .X(_02694_));
 sky130_fd_sc_hd__and2_1 _18259_ (.A(_02324_),
    .B(_00116_),
    .X(_02549_));
 sky130_fd_sc_hd__buf_1 _18260_ (.A(_13953_),
    .X(_13960_));
 sky130_fd_sc_hd__and3_1 _18261_ (.A(_13959_),
    .B(_00116_),
    .C(_13960_),
    .X(_02693_));
 sky130_fd_sc_hd__and2_1 _18262_ (.A(_13959_),
    .B(_00110_),
    .X(_02548_));
 sky130_fd_sc_hd__buf_1 _18263_ (.A(_13958_),
    .X(_13961_));
 sky130_fd_sc_hd__and3_1 _18264_ (.A(_13961_),
    .B(_00110_),
    .C(_13960_),
    .X(_02692_));
 sky130_fd_sc_hd__and2_1 _18265_ (.A(_13959_),
    .B(_00104_),
    .X(_02547_));
 sky130_fd_sc_hd__and3_1 _18266_ (.A(_13961_),
    .B(_00104_),
    .C(_13960_),
    .X(_02691_));
 sky130_vsdinv _18267_ (.A(_12740_),
    .Y(_13962_));
 sky130_fd_sc_hd__buf_1 _18268_ (.A(_13962_),
    .X(_13963_));
 sky130_fd_sc_hd__clkbuf_2 _18269_ (.A(_13963_),
    .X(_02321_));
 sky130_fd_sc_hd__buf_1 _18270_ (.A(_13957_),
    .X(_13964_));
 sky130_fd_sc_hd__and3_1 _18271_ (.A(_02321_),
    .B(_00094_),
    .C(_13964_),
    .X(_02546_));
 sky130_fd_sc_hd__and2_1 _18272_ (.A(_13963_),
    .B(_00094_),
    .X(_00095_));
 sky130_fd_sc_hd__and3_1 _18273_ (.A(_13961_),
    .B(_00095_),
    .C(_13960_),
    .X(_02690_));
 sky130_fd_sc_hd__and3_1 _18274_ (.A(_02321_),
    .B(_00084_),
    .C(_13964_),
    .X(_02545_));
 sky130_fd_sc_hd__and2_1 _18275_ (.A(_13963_),
    .B(_00084_),
    .X(_00085_));
 sky130_fd_sc_hd__and3_1 _18276_ (.A(_13961_),
    .B(_00085_),
    .C(_13954_),
    .X(_02689_));
 sky130_vsdinv _18277_ (.A(_12742_),
    .Y(_13965_));
 sky130_fd_sc_hd__buf_1 _18278_ (.A(_13965_),
    .X(_13966_));
 sky130_fd_sc_hd__and3_1 _18279_ (.A(_13966_),
    .B(_00066_),
    .C(_13962_),
    .X(_13967_));
 sky130_fd_sc_hd__buf_1 _18280_ (.A(_13967_),
    .X(_00068_));
 sky130_fd_sc_hd__nand2_1 _18281_ (.A(_13958_),
    .B(_00068_),
    .Y(_13968_));
 sky130_vsdinv _18282_ (.A(_13968_),
    .Y(_02544_));
 sky130_fd_sc_hd__nor2_1 _18283_ (.A(_12735_),
    .B(_13968_),
    .Y(_02688_));
 sky130_vsdinv _18284_ (.A(net306),
    .Y(_13969_));
 sky130_fd_sc_hd__nor2_4 _18285_ (.A(_12744_),
    .B(_13969_),
    .Y(_00048_));
 sky130_fd_sc_hd__nand2_1 _18286_ (.A(_13965_),
    .B(_00048_),
    .Y(_13970_));
 sky130_fd_sc_hd__inv_2 _18287_ (.A(_13970_),
    .Y(_00049_));
 sky130_fd_sc_hd__and3_1 _18288_ (.A(_13963_),
    .B(_00049_),
    .C(_13964_),
    .X(_02543_));
 sky130_fd_sc_hd__nor2_2 _18289_ (.A(_12740_),
    .B(_13970_),
    .Y(_00050_));
 sky130_fd_sc_hd__and3_1 _18290_ (.A(_13964_),
    .B(_00050_),
    .C(_13954_),
    .X(_02687_));
 sky130_fd_sc_hd__clkbuf_4 _18291_ (.A(_12390_),
    .X(_00297_));
 sky130_fd_sc_hd__o211a_1 _18292_ (.A1(\reg_pc[1] ),
    .A2(_13781_),
    .B1(net101),
    .C1(mem_do_rinst),
    .X(_13971_));
 sky130_fd_sc_hd__buf_1 _18293_ (.A(_13971_),
    .X(_13972_));
 sky130_fd_sc_hd__clkbuf_2 _18294_ (.A(_13972_),
    .X(_00307_));
 sky130_fd_sc_hd__or2_1 _18295_ (.A(irq_active),
    .B(\irq_mask[2] ),
    .X(_13973_));
 sky130_fd_sc_hd__buf_1 _18296_ (.A(_13973_),
    .X(_13974_));
 sky130_fd_sc_hd__buf_1 _18297_ (.A(_13974_),
    .X(_13975_));
 sky130_fd_sc_hd__buf_1 _18298_ (.A(_13975_),
    .X(_13976_));
 sky130_fd_sc_hd__clkbuf_2 _18299_ (.A(_13976_),
    .X(_13977_));
 sky130_fd_sc_hd__nor2_1 _18300_ (.A(_12394_),
    .B(_13977_),
    .Y(_00312_));
 sky130_fd_sc_hd__o21ai_2 _18301_ (.A1(mem_do_wdata),
    .A2(_11557_),
    .B1(_11542_),
    .Y(_13978_));
 sky130_fd_sc_hd__buf_1 _18302_ (.A(_13978_),
    .X(_13979_));
 sky130_vsdinv _18303_ (.A(_13979_),
    .Y(_13980_));
 sky130_fd_sc_hd__clkbuf_2 _18304_ (.A(_13980_),
    .X(_00303_));
 sky130_vsdinv _18305_ (.A(_13971_),
    .Y(_13981_));
 sky130_fd_sc_hd__or2_1 _18306_ (.A(_13981_),
    .B(_13974_),
    .X(_13982_));
 sky130_fd_sc_hd__o21a_1 _18307_ (.A1(_11617_),
    .A2(_12385_),
    .B1(_11673_),
    .X(_13983_));
 sky130_fd_sc_hd__buf_1 _18308_ (.A(_13979_),
    .X(_13984_));
 sky130_vsdinv _18309_ (.A(\mem_wordsize[2] ),
    .Y(_13985_));
 sky130_fd_sc_hd__or2_4 _18310_ (.A(_13969_),
    .B(_13985_),
    .X(_13986_));
 sky130_vsdinv _18311_ (.A(_13986_),
    .Y(_13987_));
 sky130_fd_sc_hd__buf_1 _18312_ (.A(_13987_),
    .X(_00306_));
 sky130_vsdinv _18313_ (.A(\mem_wordsize[0] ),
    .Y(_13988_));
 sky130_fd_sc_hd__nor2_8 _18314_ (.A(_13485_),
    .B(_13487_),
    .Y(_00304_));
 sky130_fd_sc_hd__or2_2 _18315_ (.A(_13988_),
    .B(_00304_),
    .X(_13989_));
 sky130_fd_sc_hd__buf_1 _18316_ (.A(_13989_),
    .X(_13990_));
 sky130_fd_sc_hd__or3_4 _18317_ (.A(_13368_),
    .B(_11618_),
    .C(_11674_),
    .X(_13991_));
 sky130_fd_sc_hd__or2_1 _18318_ (.A(_11579_),
    .B(_13991_),
    .X(_13992_));
 sky130_fd_sc_hd__or3_4 _18319_ (.A(_11617_),
    .B(_00309_),
    .C(_12385_),
    .X(_13993_));
 sky130_vsdinv _18320_ (.A(_13989_),
    .Y(_13994_));
 sky130_fd_sc_hd__o32a_1 _18321_ (.A1(_13975_),
    .A2(_13990_),
    .A3(_13992_),
    .B1(_13993_),
    .B2(_13994_),
    .X(_13995_));
 sky130_fd_sc_hd__o41a_1 _18322_ (.A1(_13974_),
    .A2(_13990_),
    .A3(_13979_),
    .A4(_00306_),
    .B1(_13980_),
    .X(_13996_));
 sky130_fd_sc_hd__or2_1 _18323_ (.A(_13993_),
    .B(_13996_),
    .X(_13997_));
 sky130_fd_sc_hd__nor2_4 _18324_ (.A(_13987_),
    .B(_13994_),
    .Y(_13998_));
 sky130_fd_sc_hd__a21oi_4 _18325_ (.A1(_11878_),
    .A2(_11558_),
    .B1(_13998_),
    .Y(_13999_));
 sky130_fd_sc_hd__nand2_1 _18326_ (.A(_11542_),
    .B(_11672_),
    .Y(_14000_));
 sky130_fd_sc_hd__or3b_2 _18327_ (.A(_13975_),
    .B(_14000_),
    .C_N(_13999_),
    .X(_14001_));
 sky130_fd_sc_hd__o221a_1 _18328_ (.A1(_12386_),
    .A2(_00303_),
    .B1(_13999_),
    .B2(_13992_),
    .C1(_14001_),
    .X(_14002_));
 sky130_fd_sc_hd__o311a_1 _18329_ (.A1(_13984_),
    .A2(_00306_),
    .A3(_13995_),
    .B1(_13997_),
    .C1(_14002_),
    .X(_14003_));
 sky130_vsdinv _18330_ (.A(_13982_),
    .Y(_14004_));
 sky130_fd_sc_hd__o21a_1 _18331_ (.A1(_13978_),
    .A2(_13998_),
    .B1(_13981_),
    .X(_14005_));
 sky130_fd_sc_hd__nor2_1 _18332_ (.A(_14004_),
    .B(_14005_),
    .Y(_14006_));
 sky130_vsdinv _18333_ (.A(_13973_),
    .Y(_14007_));
 sky130_fd_sc_hd__a31o_1 _18334_ (.A1(_14007_),
    .A2(_00306_),
    .A3(_00303_),
    .B1(_14004_),
    .X(_14008_));
 sky130_vsdinv _18335_ (.A(_14008_),
    .Y(_14009_));
 sky130_fd_sc_hd__buf_1 _18336_ (.A(_13994_),
    .X(_00305_));
 sky130_fd_sc_hd__or2_1 _18337_ (.A(_13972_),
    .B(_13987_),
    .X(_14010_));
 sky130_fd_sc_hd__or2_1 _18338_ (.A(_13979_),
    .B(_14010_),
    .X(_14011_));
 sky130_fd_sc_hd__a211o_1 _18339_ (.A1(_13976_),
    .A2(_00305_),
    .B1(_14011_),
    .C1(_12386_),
    .X(_14012_));
 sky130_fd_sc_hd__o221a_1 _18340_ (.A1(_14000_),
    .A2(_14006_),
    .B1(_13992_),
    .B2(_14009_),
    .C1(_14012_),
    .X(_14013_));
 sky130_fd_sc_hd__o221a_1 _18341_ (.A1(_13982_),
    .A2(_13983_),
    .B1(_00307_),
    .B2(_14003_),
    .C1(_14013_),
    .X(_14014_));
 sky130_fd_sc_hd__or2_2 _18342_ (.A(_14007_),
    .B(_14005_),
    .X(_14015_));
 sky130_vsdinv _18343_ (.A(_14015_),
    .Y(_14016_));
 sky130_fd_sc_hd__clkbuf_2 _18344_ (.A(_14016_),
    .X(_14017_));
 sky130_fd_sc_hd__or4_4 _18345_ (.A(_11677_),
    .B(\irq_mask[1] ),
    .C(\pcpi_mul.active[1] ),
    .D(_00311_),
    .X(_14018_));
 sky130_fd_sc_hd__o31a_1 _18346_ (.A1(_13976_),
    .A2(_13990_),
    .A3(_14011_),
    .B1(_14006_),
    .X(_14019_));
 sky130_fd_sc_hd__o22a_1 _18347_ (.A1(_11748_),
    .A2(_14017_),
    .B1(_14018_),
    .B2(_14019_),
    .X(_14020_));
 sky130_fd_sc_hd__buf_1 _18348_ (.A(_14007_),
    .X(_14021_));
 sky130_fd_sc_hd__o21ai_1 _18349_ (.A1(_14021_),
    .A2(_13998_),
    .B1(_13981_),
    .Y(_14022_));
 sky130_fd_sc_hd__or3_1 _18350_ (.A(_13974_),
    .B(_13986_),
    .C(_13972_),
    .X(_14023_));
 sky130_fd_sc_hd__o32a_1 _18351_ (.A1(_11585_),
    .A2(_12363_),
    .A3(_14018_),
    .B1(_11773_),
    .B2(_13993_),
    .X(_14024_));
 sky130_fd_sc_hd__or3_2 _18352_ (.A(_11772_),
    .B(_12386_),
    .C(_14023_),
    .X(_14025_));
 sky130_fd_sc_hd__o221a_1 _18353_ (.A1(_12392_),
    .A2(_14022_),
    .B1(_14023_),
    .B2(_14024_),
    .C1(_14025_),
    .X(_14026_));
 sky130_fd_sc_hd__o21ai_1 _18354_ (.A1(_00307_),
    .A2(_13999_),
    .B1(_13975_),
    .Y(_14027_));
 sky130_fd_sc_hd__nand2_1 _18355_ (.A(_11678_),
    .B(_14027_),
    .Y(_14028_));
 sky130_fd_sc_hd__or4_4 _18356_ (.A(_11728_),
    .B(alu_wait),
    .C(_11732_),
    .D(_11555_),
    .X(_14029_));
 sky130_fd_sc_hd__o21a_1 _18357_ (.A1(_13972_),
    .A2(_13980_),
    .B1(_13982_),
    .X(_14030_));
 sky130_fd_sc_hd__a211oi_2 _18358_ (.A1(_12874_),
    .A2(_14015_),
    .B1(_11581_),
    .C1(_00314_),
    .Y(_14031_));
 sky130_fd_sc_hd__o221a_1 _18359_ (.A1(_14016_),
    .A2(_14029_),
    .B1(_12392_),
    .B2(_14030_),
    .C1(_14031_),
    .X(_14032_));
 sky130_fd_sc_hd__o31a_1 _18360_ (.A1(_11572_),
    .A2(_11746_),
    .A3(_14028_),
    .B1(_14032_),
    .X(_14033_));
 sky130_fd_sc_hd__o221a_1 _18361_ (.A1(_12364_),
    .A2(_14020_),
    .B1(_13984_),
    .B2(_14026_),
    .C1(_14033_),
    .X(_14034_));
 sky130_fd_sc_hd__o21ai_1 _18362_ (.A1(_00322_),
    .A2(_14014_),
    .B1(_14034_),
    .Y(_00039_));
 sky130_fd_sc_hd__nor2_1 _18363_ (.A(_11810_),
    .B(_14028_),
    .Y(_00040_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _18364_ (.A(_14005_),
    .X(_14035_));
 sky130_fd_sc_hd__and3_1 _18365_ (.A(_11563_),
    .B(_14035_),
    .C(_12009_),
    .X(_14036_));
 sky130_fd_sc_hd__a31oi_1 _18366_ (.A1(_12275_),
    .A2(_14015_),
    .A3(_11799_),
    .B1(_14036_),
    .Y(_14037_));
 sky130_fd_sc_hd__clkbuf_2 _18367_ (.A(_11560_),
    .X(_14038_));
 sky130_fd_sc_hd__buf_2 _18368_ (.A(_14038_),
    .X(_14039_));
 sky130_fd_sc_hd__clkbuf_2 _18369_ (.A(_14039_),
    .X(_14040_));
 sky130_vsdinv _18370_ (.A(_11545_),
    .Y(_14041_));
 sky130_fd_sc_hd__or2_2 _18371_ (.A(_14041_),
    .B(_11794_),
    .X(_14042_));
 sky130_fd_sc_hd__buf_1 _18372_ (.A(_14017_),
    .X(_14043_));
 sky130_fd_sc_hd__or2_1 _18373_ (.A(_11580_),
    .B(_12008_),
    .X(_14044_));
 sky130_vsdinv _18374_ (.A(_12391_),
    .Y(_14045_));
 sky130_fd_sc_hd__or2_1 _18375_ (.A(_14044_),
    .B(_14045_),
    .X(_14046_));
 sky130_fd_sc_hd__o32a_1 _18376_ (.A1(_13977_),
    .A2(_14035_),
    .A3(_14042_),
    .B1(_14043_),
    .B2(_14046_),
    .X(_14047_));
 sky130_fd_sc_hd__o22ai_1 _18377_ (.A1(_12545_),
    .A2(_14037_),
    .B1(_14040_),
    .B2(_14047_),
    .Y(_00044_));
 sky130_fd_sc_hd__nor2_8 _18378_ (.A(is_jalr_addi_slti_sltiu_xori_ori_andi),
    .B(is_slli_srli_srai),
    .Y(_01304_));
 sky130_fd_sc_hd__or4b_4 _18379_ (.A(is_lui_auipc_jal),
    .B(_14017_),
    .C(_11747_),
    .D_N(_01304_),
    .X(_14048_));
 sky130_fd_sc_hd__o32a_1 _18380_ (.A1(_12364_),
    .A2(_12368_),
    .A3(_14043_),
    .B1(_11799_),
    .B2(_14048_),
    .X(_14049_));
 sky130_fd_sc_hd__nor2_1 _18381_ (.A(_12393_),
    .B(_14049_),
    .Y(_00041_));
 sky130_fd_sc_hd__a211o_1 _18382_ (.A1(_11669_),
    .A2(_11619_),
    .B1(\pcpi_mul.active[1] ),
    .C1(_00311_),
    .X(_14050_));
 sky130_fd_sc_hd__or3_1 _18383_ (.A(_12364_),
    .B(_14050_),
    .C(_14043_),
    .X(_14051_));
 sky130_fd_sc_hd__a31oi_1 _18384_ (.A1(_12551_),
    .A2(_14027_),
    .A3(_14051_),
    .B1(_12213_),
    .Y(_00038_));
 sky130_vsdinv _18385_ (.A(_12267_),
    .Y(_00315_));
 sky130_fd_sc_hd__or3_4 _18386_ (.A(_11580_),
    .B(_11800_),
    .C(_12362_),
    .X(_14052_));
 sky130_fd_sc_hd__or3_2 _18387_ (.A(_13984_),
    .B(_13990_),
    .C(_13389_),
    .X(_14053_));
 sky130_fd_sc_hd__o32a_1 _18388_ (.A1(_13976_),
    .A2(_13984_),
    .A3(_14052_),
    .B1(_14042_),
    .B2(_14053_),
    .X(_14054_));
 sky130_fd_sc_hd__o21bai_1 _18389_ (.A1(_14008_),
    .A2(_14035_),
    .B1_N(_14052_),
    .Y(_14055_));
 sky130_fd_sc_hd__a41o_1 _18390_ (.A1(_00303_),
    .A2(_00305_),
    .A3(_13981_),
    .A4(_13986_),
    .B1(_14042_),
    .X(_14056_));
 sky130_fd_sc_hd__clkbuf_2 _18391_ (.A(_13389_),
    .X(_14057_));
 sky130_fd_sc_hd__a211o_1 _18392_ (.A1(_14046_),
    .A2(_14056_),
    .B1(_14057_),
    .C1(_14017_),
    .X(_14058_));
 sky130_fd_sc_hd__o311a_1 _18393_ (.A1(_13977_),
    .A2(_14010_),
    .A3(_14054_),
    .B1(_14055_),
    .C1(_14058_),
    .X(_14059_));
 sky130_vsdinv _18394_ (.A(_14059_),
    .Y(_00043_));
 sky130_fd_sc_hd__and3_4 _18395_ (.A(_11789_),
    .B(_00290_),
    .C(_11590_),
    .X(net199));
 sky130_fd_sc_hd__buf_1 _18396_ (.A(_12795_),
    .X(_14060_));
 sky130_vsdinv _18397_ (.A(_14060_),
    .Y(net232));
 sky130_fd_sc_hd__nor2_1 _18398_ (.A(_11878_),
    .B(_14057_),
    .Y(_00317_));
 sky130_fd_sc_hd__clkbuf_4 _18399_ (.A(_11734_),
    .X(_14061_));
 sky130_fd_sc_hd__clkbuf_2 _18400_ (.A(_14061_),
    .X(_14062_));
 sky130_fd_sc_hd__or3_1 _18401_ (.A(_11728_),
    .B(_11730_),
    .C(_11794_),
    .X(_14063_));
 sky130_fd_sc_hd__o21a_1 _18402_ (.A1(_00305_),
    .A2(_14011_),
    .B1(_14009_),
    .X(_14064_));
 sky130_fd_sc_hd__o32a_1 _18403_ (.A1(_11587_),
    .A2(_00302_),
    .A3(_14043_),
    .B1(_14063_),
    .B2(_14064_),
    .X(_14065_));
 sky130_fd_sc_hd__or2_1 _18404_ (.A(_11733_),
    .B(_13996_),
    .X(_14066_));
 sky130_fd_sc_hd__o32a_1 _18405_ (.A1(_11587_),
    .A2(_13999_),
    .A3(_13950_),
    .B1(_14063_),
    .B2(_14066_),
    .X(_14067_));
 sky130_fd_sc_hd__o32a_1 _18406_ (.A1(_13977_),
    .A2(_14035_),
    .A3(_13950_),
    .B1(_13951_),
    .B2(_14028_),
    .X(_14068_));
 sky130_fd_sc_hd__o221ai_1 _18407_ (.A1(_14062_),
    .A2(_14065_),
    .B1(_00307_),
    .B2(_14067_),
    .C1(_14068_),
    .Y(_00042_));
 sky130_vsdinv _18408_ (.A(_12744_),
    .Y(_14069_));
 sky130_fd_sc_hd__nor2_1 _18409_ (.A(_14069_),
    .B(_13487_),
    .Y(_14070_));
 sky130_fd_sc_hd__or2_2 _18410_ (.A(_00048_),
    .B(_14070_),
    .X(_02591_));
 sky130_fd_sc_hd__nor2_2 _18411_ (.A(net353),
    .B(_13419_),
    .Y(_14071_));
 sky130_fd_sc_hd__a21oi_4 _18412_ (.A1(net353),
    .A2(_13420_),
    .B1(_14071_),
    .Y(_14072_));
 sky130_fd_sc_hd__nor2_2 _18413_ (.A(net351),
    .B(_13424_),
    .Y(_14073_));
 sky130_fd_sc_hd__a21oi_2 _18414_ (.A1(net351),
    .A2(_13425_),
    .B1(_14073_),
    .Y(_14074_));
 sky130_fd_sc_hd__nor2_2 _18415_ (.A(net352),
    .B(_13422_),
    .Y(_14075_));
 sky130_fd_sc_hd__a21oi_2 _18416_ (.A1(_12699_),
    .A2(_13423_),
    .B1(_14075_),
    .Y(_14076_));
 sky130_fd_sc_hd__nor2_2 _18417_ (.A(net350),
    .B(_13426_),
    .Y(_14077_));
 sky130_fd_sc_hd__a21oi_4 _18418_ (.A1(_12701_),
    .A2(_13427_),
    .B1(_14077_),
    .Y(_14078_));
 sky130_fd_sc_hd__or4_4 _18419_ (.A(_14072_),
    .B(_14074_),
    .C(_14076_),
    .D(_14078_),
    .X(_14079_));
 sky130_fd_sc_hd__nor2_1 _18420_ (.A(_12707_),
    .B(_13437_),
    .Y(_14080_));
 sky130_fd_sc_hd__a21oi_2 _18421_ (.A1(_12707_),
    .A2(_13438_),
    .B1(_14080_),
    .Y(_14081_));
 sky130_fd_sc_hd__nor2_2 _18422_ (.A(net347),
    .B(_13432_),
    .Y(_14082_));
 sky130_fd_sc_hd__a21oi_4 _18423_ (.A1(_12705_),
    .A2(_13433_),
    .B1(_14082_),
    .Y(_14083_));
 sky130_fd_sc_hd__nor2_1 _18424_ (.A(net346),
    .B(_13434_),
    .Y(_14084_));
 sky130_fd_sc_hd__a21oi_2 _18425_ (.A1(net346),
    .A2(_13435_),
    .B1(_14084_),
    .Y(_14085_));
 sky130_fd_sc_hd__nor2_2 _18426_ (.A(net348),
    .B(_13429_),
    .Y(_14086_));
 sky130_fd_sc_hd__a21oi_4 _18427_ (.A1(_12703_),
    .A2(_13430_),
    .B1(_14086_),
    .Y(_14087_));
 sky130_fd_sc_hd__or4_4 _18428_ (.A(_14081_),
    .B(_14083_),
    .C(_14085_),
    .D(_14087_),
    .X(_14088_));
 sky130_fd_sc_hd__nor2_2 _18429_ (.A(net359),
    .B(net327),
    .Y(_14089_));
 sky130_fd_sc_hd__a21oi_4 _18430_ (.A1(net359),
    .A2(_13400_),
    .B1(_14089_),
    .Y(_14090_));
 sky130_fd_sc_hd__nor2_1 _18431_ (.A(net358),
    .B(net326),
    .Y(_14091_));
 sky130_fd_sc_hd__a21oi_2 _18432_ (.A1(_12688_),
    .A2(_13403_),
    .B1(_14091_),
    .Y(_14092_));
 sky130_fd_sc_hd__nor2_2 _18433_ (.A(net330),
    .B(net362),
    .Y(_14093_));
 sky130_fd_sc_hd__a21oi_4 _18434_ (.A1(net330),
    .A2(net362),
    .B1(_14093_),
    .Y(_14094_));
 sky130_fd_sc_hd__nor2_1 _18435_ (.A(net361),
    .B(net329),
    .Y(_14095_));
 sky130_fd_sc_hd__a21oi_1 _18436_ (.A1(net361),
    .A2(_13398_),
    .B1(_14095_),
    .Y(_14096_));
 sky130_fd_sc_hd__or2_1 _18437_ (.A(_14094_),
    .B(_14096_),
    .X(_14097_));
 sky130_fd_sc_hd__nor2_1 _18438_ (.A(net357),
    .B(net325),
    .Y(_14098_));
 sky130_fd_sc_hd__a21oi_2 _18439_ (.A1(net357),
    .A2(_13407_),
    .B1(_14098_),
    .Y(_14099_));
 sky130_fd_sc_hd__nor2_1 _18440_ (.A(net356),
    .B(net324),
    .Y(_14100_));
 sky130_fd_sc_hd__a21oi_2 _18441_ (.A1(_12693_),
    .A2(net324),
    .B1(_14100_),
    .Y(_14101_));
 sky130_fd_sc_hd__nor2_1 _18442_ (.A(net355),
    .B(net323),
    .Y(_14102_));
 sky130_fd_sc_hd__a21oi_2 _18443_ (.A1(net355),
    .A2(net323),
    .B1(_14102_),
    .Y(_14103_));
 sky130_fd_sc_hd__nor2_1 _18444_ (.A(_12695_),
    .B(_13416_),
    .Y(_14104_));
 sky130_fd_sc_hd__a21oi_2 _18445_ (.A1(_12695_),
    .A2(_13416_),
    .B1(_14104_),
    .Y(_14105_));
 sky130_fd_sc_hd__or4_4 _18446_ (.A(_14099_),
    .B(_14101_),
    .C(_14103_),
    .D(_14105_),
    .X(_14106_));
 sky130_fd_sc_hd__or4_4 _18447_ (.A(_14090_),
    .B(_14092_),
    .C(_14097_),
    .D(_14106_),
    .X(_14107_));
 sky130_fd_sc_hd__nor2_2 _18448_ (.A(net227),
    .B(_13471_),
    .Y(_14108_));
 sky130_fd_sc_hd__a21oi_4 _18449_ (.A1(_12732_),
    .A2(_13471_),
    .B1(_14108_),
    .Y(_14109_));
 sky130_fd_sc_hd__nor2_4 _18450_ (.A(net229),
    .B(_13464_),
    .Y(_14110_));
 sky130_fd_sc_hd__a21oi_4 _18451_ (.A1(_12727_),
    .A2(_13465_),
    .B1(_14110_),
    .Y(_14111_));
 sky130_fd_sc_hd__nor2_2 _18452_ (.A(_12742_),
    .B(_13485_),
    .Y(_14112_));
 sky130_fd_sc_hd__a21oi_2 _18453_ (.A1(_12742_),
    .A2(_13485_),
    .B1(_14112_),
    .Y(_14113_));
 sky130_fd_sc_hd__nor2_1 _18454_ (.A(net225),
    .B(_13478_),
    .Y(_14114_));
 sky130_fd_sc_hd__a21oi_2 _18455_ (.A1(_12737_),
    .A2(_13478_),
    .B1(_14114_),
    .Y(_14115_));
 sky130_fd_sc_hd__or4_4 _18456_ (.A(_14109_),
    .B(_14111_),
    .C(_14113_),
    .D(_14115_),
    .X(_14116_));
 sky130_fd_sc_hd__nor2_1 _18457_ (.A(net226),
    .B(_13474_),
    .Y(_14117_));
 sky130_fd_sc_hd__a21oi_2 _18458_ (.A1(_12734_),
    .A2(_13474_),
    .B1(_14117_),
    .Y(_14118_));
 sky130_fd_sc_hd__nor2_2 _18459_ (.A(_12730_),
    .B(_13468_),
    .Y(_14119_));
 sky130_fd_sc_hd__a21oi_4 _18460_ (.A1(_12730_),
    .A2(_13468_),
    .B1(_14119_),
    .Y(_14120_));
 sky130_fd_sc_hd__nor2_2 _18461_ (.A(net222),
    .B(_13482_),
    .Y(_14121_));
 sky130_fd_sc_hd__a21oi_4 _18462_ (.A1(net222),
    .A2(_13482_),
    .B1(_14121_),
    .Y(_14122_));
 sky130_fd_sc_hd__or4_4 _18463_ (.A(_02591_),
    .B(_14118_),
    .C(_14120_),
    .D(_14122_),
    .X(_14123_));
 sky130_fd_sc_hd__nor2_2 _18464_ (.A(_12710_),
    .B(_13441_),
    .Y(_14124_));
 sky130_fd_sc_hd__a21oi_4 _18465_ (.A1(_12710_),
    .A2(_13442_),
    .B1(_14124_),
    .Y(_14125_));
 sky130_fd_sc_hd__nor2_1 _18466_ (.A(net341),
    .B(_13449_),
    .Y(_14126_));
 sky130_fd_sc_hd__a21oi_2 _18467_ (.A1(_12717_),
    .A2(_13450_),
    .B1(_14126_),
    .Y(_14127_));
 sky130_fd_sc_hd__nor2_2 _18468_ (.A(_12715_),
    .B(_13447_),
    .Y(_14128_));
 sky130_fd_sc_hd__a21oi_2 _18469_ (.A1(_12715_),
    .A2(_13448_),
    .B1(_14128_),
    .Y(_14129_));
 sky130_fd_sc_hd__nor2_2 _18470_ (.A(net343),
    .B(_13445_),
    .Y(_14130_));
 sky130_fd_sc_hd__a21oi_4 _18471_ (.A1(net343),
    .A2(_13446_),
    .B1(_14130_),
    .Y(_14131_));
 sky130_fd_sc_hd__or4_4 _18472_ (.A(_14125_),
    .B(_14127_),
    .C(_14129_),
    .D(_14131_),
    .X(_14132_));
 sky130_fd_sc_hd__nor2_1 _18473_ (.A(_12719_),
    .B(_13452_),
    .Y(_14133_));
 sky130_fd_sc_hd__a21oi_2 _18474_ (.A1(_12719_),
    .A2(_13453_),
    .B1(_14133_),
    .Y(_14134_));
 sky130_fd_sc_hd__nor2_1 _18475_ (.A(net368),
    .B(_13460_),
    .Y(_14135_));
 sky130_fd_sc_hd__a21oi_2 _18476_ (.A1(_12725_),
    .A2(_13461_),
    .B1(_14135_),
    .Y(_14136_));
 sky130_fd_sc_hd__nor2_2 _18477_ (.A(_12723_),
    .B(_13457_),
    .Y(_14137_));
 sky130_fd_sc_hd__a21oi_4 _18478_ (.A1(_12723_),
    .A2(_13458_),
    .B1(_14137_),
    .Y(_14138_));
 sky130_fd_sc_hd__nor2_2 _18479_ (.A(net339),
    .B(_13455_),
    .Y(_14139_));
 sky130_fd_sc_hd__a21oi_4 _18480_ (.A1(_12722_),
    .A2(_13456_),
    .B1(_14139_),
    .Y(_14140_));
 sky130_fd_sc_hd__or4_4 _18481_ (.A(_14134_),
    .B(_14136_),
    .C(_14138_),
    .D(_14140_),
    .X(_14141_));
 sky130_fd_sc_hd__or4_4 _18482_ (.A(_14116_),
    .B(_14123_),
    .C(_14132_),
    .D(_14141_),
    .X(_14142_));
 sky130_fd_sc_hd__or4_4 _18483_ (.A(_14079_),
    .B(_14088_),
    .C(_14107_),
    .D(_14142_),
    .X(_14143_));
 sky130_fd_sc_hd__inv_2 _18484_ (.A(_14143_),
    .Y(_00000_));
 sky130_fd_sc_hd__or2_1 _18485_ (.A(_11697_),
    .B(_11698_),
    .X(\pcpi_mul.instr_any_mulh ));
 sky130_fd_sc_hd__or3_2 _18486_ (.A(instr_slt),
    .B(instr_slti),
    .C(instr_blt),
    .X(_00006_));
 sky130_fd_sc_hd__or3_2 _18487_ (.A(instr_sltu),
    .B(instr_sltiu),
    .C(instr_bltu),
    .X(_00007_));
 sky130_fd_sc_hd__or2_1 _18488_ (.A(net415),
    .B(_13183_),
    .X(_00299_));
 sky130_vsdinv _18489_ (.A(instr_sh),
    .Y(_14144_));
 sky130_fd_sc_hd__nor2_1 _18490_ (.A(instr_lhu),
    .B(instr_lh),
    .Y(_14145_));
 sky130_fd_sc_hd__o32a_1 _18491_ (.A1(_14144_),
    .A2(_14057_),
    .A3(_12010_),
    .B1(_12014_),
    .B2(_14145_),
    .X(_14146_));
 sky130_fd_sc_hd__clkbuf_2 _18492_ (.A(_13985_),
    .X(_14147_));
 sky130_fd_sc_hd__clkbuf_2 _18493_ (.A(_14147_),
    .X(_14148_));
 sky130_fd_sc_hd__nor2_1 _18494_ (.A(_00319_),
    .B(_00317_),
    .Y(_14149_));
 sky130_fd_sc_hd__o21a_1 _18495_ (.A1(_11781_),
    .A2(_11806_),
    .B1(_11678_),
    .X(_14150_));
 sky130_fd_sc_hd__o221a_1 _18496_ (.A1(_00297_),
    .A2(_14042_),
    .B1(_12009_),
    .B2(_14149_),
    .C1(_14150_),
    .X(_14151_));
 sky130_fd_sc_hd__o22ai_1 _18497_ (.A1(_00296_),
    .A2(_14146_),
    .B1(_14148_),
    .B2(_14151_),
    .Y(_00047_));
 sky130_fd_sc_hd__clkbuf_4 _18498_ (.A(_11879_),
    .X(_00301_));
 sky130_fd_sc_hd__clkbuf_4 _18499_ (.A(_11725_),
    .X(_14152_));
 sky130_fd_sc_hd__buf_2 _18500_ (.A(_14152_),
    .X(_14153_));
 sky130_fd_sc_hd__nor2_1 _18501_ (.A(_14153_),
    .B(_11806_),
    .Y(_00336_));
 sky130_fd_sc_hd__nor2_1 _18502_ (.A(_14286_),
    .B(_14045_),
    .Y(_00338_));
 sky130_vsdinv _18503_ (.A(alu_eq),
    .Y(_00340_));
 sky130_fd_sc_hd__or3_4 _18504_ (.A(instr_bne),
    .B(is_slti_blt_slt),
    .C(is_sltiu_bltu_sltu),
    .X(_14154_));
 sky130_fd_sc_hd__nor3_4 _18505_ (.A(instr_bgeu),
    .B(instr_bge),
    .C(_14154_),
    .Y(_00341_));
 sky130_fd_sc_hd__mux2_1 _18506_ (.A0(instr_bgeu),
    .A1(is_sltiu_bltu_sltu),
    .S(alu_ltu),
    .X(_14155_));
 sky130_fd_sc_hd__a21oi_1 _18507_ (.A1(is_slti_blt_slt),
    .A2(alu_lts),
    .B1(_14155_),
    .Y(_14156_));
 sky130_fd_sc_hd__o221a_1 _18508_ (.A1(_11995_),
    .A2(alu_eq),
    .B1(_11989_),
    .B2(alu_lts),
    .C1(_14156_),
    .X(_00342_));
 sky130_vsdinv _18509_ (.A(_00343_),
    .Y(_14157_));
 sky130_fd_sc_hd__or2_1 _18510_ (.A(_14157_),
    .B(_11896_),
    .X(_00344_));
 sky130_fd_sc_hd__o22ai_1 _18511_ (.A1(_00339_),
    .A2(_00297_),
    .B1(_14062_),
    .B2(_00346_),
    .Y(_00347_));
 sky130_fd_sc_hd__o21a_1 _18512_ (.A1(_11617_),
    .A2(do_waitirq),
    .B1(_11777_),
    .X(_00349_));
 sky130_fd_sc_hd__and2_1 _18513_ (.A(_02410_),
    .B(_00349_),
    .X(_00351_));
 sky130_fd_sc_hd__buf_2 _18514_ (.A(_12362_),
    .X(_14158_));
 sky130_fd_sc_hd__and3_1 _18515_ (.A(_12280_),
    .B(_14158_),
    .C(_11733_),
    .X(_00354_));
 sky130_fd_sc_hd__buf_2 _18516_ (.A(_11734_),
    .X(_14159_));
 sky130_fd_sc_hd__buf_1 _18517_ (.A(_12280_),
    .X(_14160_));
 sky130_fd_sc_hd__clkbuf_2 _18518_ (.A(_14160_),
    .X(_14161_));
 sky130_fd_sc_hd__o211a_1 _18519_ (.A1(_14159_),
    .A2(_14041_),
    .B1(_14161_),
    .C1(_14158_),
    .X(_00355_));
 sky130_vsdinv _18520_ (.A(\cpuregs[0][1] ),
    .Y(_00371_));
 sky130_vsdinv _18521_ (.A(\cpuregs[1][1] ),
    .Y(_00372_));
 sky130_vsdinv _18522_ (.A(\cpuregs[2][1] ),
    .Y(_00373_));
 sky130_vsdinv _18523_ (.A(\cpuregs[3][1] ),
    .Y(_00374_));
 sky130_vsdinv _18524_ (.A(\cpuregs[4][1] ),
    .Y(_00376_));
 sky130_vsdinv _18525_ (.A(\cpuregs[5][1] ),
    .Y(_00377_));
 sky130_vsdinv _18526_ (.A(\cpuregs[6][1] ),
    .Y(_00378_));
 sky130_vsdinv _18527_ (.A(\cpuregs[7][1] ),
    .Y(_00379_));
 sky130_vsdinv _18528_ (.A(\cpuregs[8][1] ),
    .Y(_00381_));
 sky130_vsdinv _18529_ (.A(\cpuregs[9][1] ),
    .Y(_00382_));
 sky130_vsdinv _18530_ (.A(\cpuregs[10][1] ),
    .Y(_00383_));
 sky130_vsdinv _18531_ (.A(\cpuregs[11][1] ),
    .Y(_00384_));
 sky130_vsdinv _18532_ (.A(\cpuregs[12][1] ),
    .Y(_00386_));
 sky130_vsdinv _18533_ (.A(\cpuregs[13][1] ),
    .Y(_00387_));
 sky130_vsdinv _18534_ (.A(\cpuregs[14][1] ),
    .Y(_00388_));
 sky130_vsdinv _18535_ (.A(\cpuregs[15][1] ),
    .Y(_00389_));
 sky130_vsdinv _18536_ (.A(\cpuregs[16][1] ),
    .Y(_00392_));
 sky130_vsdinv _18537_ (.A(\cpuregs[17][1] ),
    .Y(_00393_));
 sky130_vsdinv _18538_ (.A(\cpuregs[18][1] ),
    .Y(_00394_));
 sky130_vsdinv _18539_ (.A(\cpuregs[19][1] ),
    .Y(_00395_));
 sky130_vsdinv _18540_ (.A(\cpuregs[0][2] ),
    .Y(_00398_));
 sky130_vsdinv _18541_ (.A(\cpuregs[1][2] ),
    .Y(_00399_));
 sky130_vsdinv _18542_ (.A(\cpuregs[2][2] ),
    .Y(_00400_));
 sky130_vsdinv _18543_ (.A(\cpuregs[3][2] ),
    .Y(_00401_));
 sky130_vsdinv _18544_ (.A(\cpuregs[4][2] ),
    .Y(_00403_));
 sky130_vsdinv _18545_ (.A(\cpuregs[5][2] ),
    .Y(_00404_));
 sky130_vsdinv _18546_ (.A(\cpuregs[6][2] ),
    .Y(_00405_));
 sky130_vsdinv _18547_ (.A(\cpuregs[7][2] ),
    .Y(_00406_));
 sky130_vsdinv _18548_ (.A(\cpuregs[8][2] ),
    .Y(_00408_));
 sky130_vsdinv _18549_ (.A(\cpuregs[9][2] ),
    .Y(_00409_));
 sky130_vsdinv _18550_ (.A(\cpuregs[10][2] ),
    .Y(_00410_));
 sky130_vsdinv _18551_ (.A(\cpuregs[11][2] ),
    .Y(_00411_));
 sky130_vsdinv _18552_ (.A(\cpuregs[12][2] ),
    .Y(_00413_));
 sky130_vsdinv _18553_ (.A(\cpuregs[13][2] ),
    .Y(_00414_));
 sky130_vsdinv _18554_ (.A(\cpuregs[14][2] ),
    .Y(_00415_));
 sky130_vsdinv _18555_ (.A(\cpuregs[15][2] ),
    .Y(_00416_));
 sky130_vsdinv _18556_ (.A(\cpuregs[16][2] ),
    .Y(_00419_));
 sky130_vsdinv _18557_ (.A(\cpuregs[17][2] ),
    .Y(_00420_));
 sky130_vsdinv _18558_ (.A(\cpuregs[18][2] ),
    .Y(_00421_));
 sky130_vsdinv _18559_ (.A(\cpuregs[19][2] ),
    .Y(_00422_));
 sky130_vsdinv _18560_ (.A(\cpuregs[0][3] ),
    .Y(_00425_));
 sky130_vsdinv _18561_ (.A(\cpuregs[1][3] ),
    .Y(_00426_));
 sky130_vsdinv _18562_ (.A(\cpuregs[2][3] ),
    .Y(_00427_));
 sky130_vsdinv _18563_ (.A(\cpuregs[3][3] ),
    .Y(_00428_));
 sky130_vsdinv _18564_ (.A(\cpuregs[4][3] ),
    .Y(_00430_));
 sky130_vsdinv _18565_ (.A(\cpuregs[5][3] ),
    .Y(_00431_));
 sky130_vsdinv _18566_ (.A(\cpuregs[6][3] ),
    .Y(_00432_));
 sky130_vsdinv _18567_ (.A(\cpuregs[7][3] ),
    .Y(_00433_));
 sky130_vsdinv _18568_ (.A(\cpuregs[8][3] ),
    .Y(_00435_));
 sky130_vsdinv _18569_ (.A(\cpuregs[9][3] ),
    .Y(_00436_));
 sky130_vsdinv _18570_ (.A(\cpuregs[10][3] ),
    .Y(_00437_));
 sky130_vsdinv _18571_ (.A(\cpuregs[11][3] ),
    .Y(_00438_));
 sky130_vsdinv _18572_ (.A(\cpuregs[12][3] ),
    .Y(_00440_));
 sky130_vsdinv _18573_ (.A(\cpuregs[13][3] ),
    .Y(_00441_));
 sky130_vsdinv _18574_ (.A(\cpuregs[14][3] ),
    .Y(_00442_));
 sky130_vsdinv _18575_ (.A(\cpuregs[15][3] ),
    .Y(_00443_));
 sky130_vsdinv _18576_ (.A(\cpuregs[16][3] ),
    .Y(_00446_));
 sky130_vsdinv _18577_ (.A(\cpuregs[17][3] ),
    .Y(_00447_));
 sky130_vsdinv _18578_ (.A(\cpuregs[18][3] ),
    .Y(_00448_));
 sky130_vsdinv _18579_ (.A(\cpuregs[19][3] ),
    .Y(_00449_));
 sky130_vsdinv _18580_ (.A(\cpuregs[0][4] ),
    .Y(_00452_));
 sky130_vsdinv _18581_ (.A(\cpuregs[1][4] ),
    .Y(_00453_));
 sky130_vsdinv _18582_ (.A(\cpuregs[2][4] ),
    .Y(_00454_));
 sky130_vsdinv _18583_ (.A(\cpuregs[3][4] ),
    .Y(_00455_));
 sky130_vsdinv _18584_ (.A(\cpuregs[4][4] ),
    .Y(_00457_));
 sky130_vsdinv _18585_ (.A(\cpuregs[5][4] ),
    .Y(_00458_));
 sky130_vsdinv _18586_ (.A(\cpuregs[6][4] ),
    .Y(_00459_));
 sky130_vsdinv _18587_ (.A(\cpuregs[7][4] ),
    .Y(_00460_));
 sky130_vsdinv _18588_ (.A(\cpuregs[8][4] ),
    .Y(_00462_));
 sky130_vsdinv _18589_ (.A(\cpuregs[9][4] ),
    .Y(_00463_));
 sky130_vsdinv _18590_ (.A(\cpuregs[10][4] ),
    .Y(_00464_));
 sky130_vsdinv _18591_ (.A(\cpuregs[11][4] ),
    .Y(_00465_));
 sky130_vsdinv _18592_ (.A(\cpuregs[12][4] ),
    .Y(_00467_));
 sky130_vsdinv _18593_ (.A(\cpuregs[13][4] ),
    .Y(_00468_));
 sky130_vsdinv _18594_ (.A(\cpuregs[14][4] ),
    .Y(_00469_));
 sky130_vsdinv _18595_ (.A(\cpuregs[15][4] ),
    .Y(_00470_));
 sky130_vsdinv _18596_ (.A(\cpuregs[16][4] ),
    .Y(_00473_));
 sky130_vsdinv _18597_ (.A(\cpuregs[17][4] ),
    .Y(_00474_));
 sky130_vsdinv _18598_ (.A(\cpuregs[18][4] ),
    .Y(_00475_));
 sky130_vsdinv _18599_ (.A(\cpuregs[19][4] ),
    .Y(_00476_));
 sky130_vsdinv _18600_ (.A(\cpuregs[0][5] ),
    .Y(_00479_));
 sky130_vsdinv _18601_ (.A(\cpuregs[1][5] ),
    .Y(_00480_));
 sky130_vsdinv _18602_ (.A(\cpuregs[2][5] ),
    .Y(_00481_));
 sky130_vsdinv _18603_ (.A(\cpuregs[3][5] ),
    .Y(_00482_));
 sky130_vsdinv _18604_ (.A(\cpuregs[4][5] ),
    .Y(_00484_));
 sky130_vsdinv _18605_ (.A(\cpuregs[5][5] ),
    .Y(_00485_));
 sky130_vsdinv _18606_ (.A(\cpuregs[6][5] ),
    .Y(_00486_));
 sky130_vsdinv _18607_ (.A(\cpuregs[7][5] ),
    .Y(_00487_));
 sky130_vsdinv _18608_ (.A(\cpuregs[8][5] ),
    .Y(_00489_));
 sky130_vsdinv _18609_ (.A(\cpuregs[9][5] ),
    .Y(_00490_));
 sky130_vsdinv _18610_ (.A(\cpuregs[10][5] ),
    .Y(_00491_));
 sky130_vsdinv _18611_ (.A(\cpuregs[11][5] ),
    .Y(_00492_));
 sky130_vsdinv _18612_ (.A(\cpuregs[12][5] ),
    .Y(_00494_));
 sky130_vsdinv _18613_ (.A(\cpuregs[13][5] ),
    .Y(_00495_));
 sky130_vsdinv _18614_ (.A(\cpuregs[14][5] ),
    .Y(_00496_));
 sky130_vsdinv _18615_ (.A(\cpuregs[15][5] ),
    .Y(_00497_));
 sky130_vsdinv _18616_ (.A(\cpuregs[16][5] ),
    .Y(_00500_));
 sky130_vsdinv _18617_ (.A(\cpuregs[17][5] ),
    .Y(_00501_));
 sky130_vsdinv _18618_ (.A(\cpuregs[18][5] ),
    .Y(_00502_));
 sky130_vsdinv _18619_ (.A(\cpuregs[19][5] ),
    .Y(_00503_));
 sky130_vsdinv _18620_ (.A(\cpuregs[0][6] ),
    .Y(_00506_));
 sky130_vsdinv _18621_ (.A(\cpuregs[1][6] ),
    .Y(_00507_));
 sky130_vsdinv _18622_ (.A(\cpuregs[2][6] ),
    .Y(_00508_));
 sky130_vsdinv _18623_ (.A(\cpuregs[3][6] ),
    .Y(_00509_));
 sky130_vsdinv _18624_ (.A(\cpuregs[4][6] ),
    .Y(_00511_));
 sky130_vsdinv _18625_ (.A(\cpuregs[5][6] ),
    .Y(_00512_));
 sky130_vsdinv _18626_ (.A(\cpuregs[6][6] ),
    .Y(_00513_));
 sky130_vsdinv _18627_ (.A(\cpuregs[7][6] ),
    .Y(_00514_));
 sky130_vsdinv _18628_ (.A(\cpuregs[8][6] ),
    .Y(_00516_));
 sky130_vsdinv _18629_ (.A(\cpuregs[9][6] ),
    .Y(_00517_));
 sky130_vsdinv _18630_ (.A(\cpuregs[10][6] ),
    .Y(_00518_));
 sky130_vsdinv _18631_ (.A(\cpuregs[11][6] ),
    .Y(_00519_));
 sky130_vsdinv _18632_ (.A(\cpuregs[12][6] ),
    .Y(_00521_));
 sky130_vsdinv _18633_ (.A(\cpuregs[13][6] ),
    .Y(_00522_));
 sky130_vsdinv _18634_ (.A(\cpuregs[14][6] ),
    .Y(_00523_));
 sky130_vsdinv _18635_ (.A(\cpuregs[15][6] ),
    .Y(_00524_));
 sky130_vsdinv _18636_ (.A(\cpuregs[16][6] ),
    .Y(_00527_));
 sky130_vsdinv _18637_ (.A(\cpuregs[17][6] ),
    .Y(_00528_));
 sky130_vsdinv _18638_ (.A(\cpuregs[18][6] ),
    .Y(_00529_));
 sky130_vsdinv _18639_ (.A(\cpuregs[19][6] ),
    .Y(_00530_));
 sky130_vsdinv _18640_ (.A(\cpuregs[0][7] ),
    .Y(_00533_));
 sky130_vsdinv _18641_ (.A(\cpuregs[1][7] ),
    .Y(_00534_));
 sky130_vsdinv _18642_ (.A(\cpuregs[2][7] ),
    .Y(_00535_));
 sky130_vsdinv _18643_ (.A(\cpuregs[3][7] ),
    .Y(_00536_));
 sky130_vsdinv _18644_ (.A(\cpuregs[4][7] ),
    .Y(_00538_));
 sky130_vsdinv _18645_ (.A(\cpuregs[5][7] ),
    .Y(_00539_));
 sky130_vsdinv _18646_ (.A(\cpuregs[6][7] ),
    .Y(_00540_));
 sky130_vsdinv _18647_ (.A(\cpuregs[7][7] ),
    .Y(_00541_));
 sky130_vsdinv _18648_ (.A(\cpuregs[8][7] ),
    .Y(_00543_));
 sky130_vsdinv _18649_ (.A(\cpuregs[9][7] ),
    .Y(_00544_));
 sky130_vsdinv _18650_ (.A(\cpuregs[10][7] ),
    .Y(_00545_));
 sky130_vsdinv _18651_ (.A(\cpuregs[11][7] ),
    .Y(_00546_));
 sky130_vsdinv _18652_ (.A(\cpuregs[12][7] ),
    .Y(_00548_));
 sky130_vsdinv _18653_ (.A(\cpuregs[13][7] ),
    .Y(_00549_));
 sky130_vsdinv _18654_ (.A(\cpuregs[14][7] ),
    .Y(_00550_));
 sky130_vsdinv _18655_ (.A(\cpuregs[15][7] ),
    .Y(_00551_));
 sky130_vsdinv _18656_ (.A(\cpuregs[16][7] ),
    .Y(_00554_));
 sky130_vsdinv _18657_ (.A(\cpuregs[17][7] ),
    .Y(_00555_));
 sky130_vsdinv _18658_ (.A(\cpuregs[18][7] ),
    .Y(_00556_));
 sky130_vsdinv _18659_ (.A(\cpuregs[19][7] ),
    .Y(_00557_));
 sky130_vsdinv _18660_ (.A(\cpuregs[0][8] ),
    .Y(_00560_));
 sky130_vsdinv _18661_ (.A(\cpuregs[1][8] ),
    .Y(_00561_));
 sky130_vsdinv _18662_ (.A(\cpuregs[2][8] ),
    .Y(_00562_));
 sky130_vsdinv _18663_ (.A(\cpuregs[3][8] ),
    .Y(_00563_));
 sky130_vsdinv _18664_ (.A(\cpuregs[4][8] ),
    .Y(_00565_));
 sky130_vsdinv _18665_ (.A(\cpuregs[5][8] ),
    .Y(_00566_));
 sky130_vsdinv _18666_ (.A(\cpuregs[6][8] ),
    .Y(_00567_));
 sky130_vsdinv _18667_ (.A(\cpuregs[7][8] ),
    .Y(_00568_));
 sky130_vsdinv _18668_ (.A(\cpuregs[8][8] ),
    .Y(_00570_));
 sky130_vsdinv _18669_ (.A(\cpuregs[9][8] ),
    .Y(_00571_));
 sky130_vsdinv _18670_ (.A(\cpuregs[10][8] ),
    .Y(_00572_));
 sky130_vsdinv _18671_ (.A(\cpuregs[11][8] ),
    .Y(_00573_));
 sky130_vsdinv _18672_ (.A(\cpuregs[12][8] ),
    .Y(_00575_));
 sky130_vsdinv _18673_ (.A(\cpuregs[13][8] ),
    .Y(_00576_));
 sky130_vsdinv _18674_ (.A(\cpuregs[14][8] ),
    .Y(_00577_));
 sky130_vsdinv _18675_ (.A(\cpuregs[15][8] ),
    .Y(_00578_));
 sky130_vsdinv _18676_ (.A(\cpuregs[16][8] ),
    .Y(_00581_));
 sky130_vsdinv _18677_ (.A(\cpuregs[17][8] ),
    .Y(_00582_));
 sky130_vsdinv _18678_ (.A(\cpuregs[18][8] ),
    .Y(_00583_));
 sky130_vsdinv _18679_ (.A(\cpuregs[19][8] ),
    .Y(_00584_));
 sky130_vsdinv _18680_ (.A(\cpuregs[0][9] ),
    .Y(_00587_));
 sky130_vsdinv _18681_ (.A(\cpuregs[1][9] ),
    .Y(_00588_));
 sky130_vsdinv _18682_ (.A(\cpuregs[2][9] ),
    .Y(_00589_));
 sky130_vsdinv _18683_ (.A(\cpuregs[3][9] ),
    .Y(_00590_));
 sky130_vsdinv _18684_ (.A(\cpuregs[4][9] ),
    .Y(_00592_));
 sky130_vsdinv _18685_ (.A(\cpuregs[5][9] ),
    .Y(_00593_));
 sky130_vsdinv _18686_ (.A(\cpuregs[6][9] ),
    .Y(_00594_));
 sky130_vsdinv _18687_ (.A(\cpuregs[7][9] ),
    .Y(_00595_));
 sky130_vsdinv _18688_ (.A(\cpuregs[8][9] ),
    .Y(_00597_));
 sky130_vsdinv _18689_ (.A(\cpuregs[9][9] ),
    .Y(_00598_));
 sky130_vsdinv _18690_ (.A(\cpuregs[10][9] ),
    .Y(_00599_));
 sky130_vsdinv _18691_ (.A(\cpuregs[11][9] ),
    .Y(_00600_));
 sky130_vsdinv _18692_ (.A(\cpuregs[12][9] ),
    .Y(_00602_));
 sky130_vsdinv _18693_ (.A(\cpuregs[13][9] ),
    .Y(_00603_));
 sky130_vsdinv _18694_ (.A(\cpuregs[14][9] ),
    .Y(_00604_));
 sky130_vsdinv _18695_ (.A(\cpuregs[15][9] ),
    .Y(_00605_));
 sky130_vsdinv _18696_ (.A(\cpuregs[16][9] ),
    .Y(_00608_));
 sky130_vsdinv _18697_ (.A(\cpuregs[17][9] ),
    .Y(_00609_));
 sky130_vsdinv _18698_ (.A(\cpuregs[18][9] ),
    .Y(_00610_));
 sky130_vsdinv _18699_ (.A(\cpuregs[19][9] ),
    .Y(_00611_));
 sky130_vsdinv _18700_ (.A(\cpuregs[0][10] ),
    .Y(_00614_));
 sky130_vsdinv _18701_ (.A(\cpuregs[1][10] ),
    .Y(_00615_));
 sky130_vsdinv _18702_ (.A(\cpuregs[2][10] ),
    .Y(_00616_));
 sky130_vsdinv _18703_ (.A(\cpuregs[3][10] ),
    .Y(_00617_));
 sky130_vsdinv _18704_ (.A(\cpuregs[4][10] ),
    .Y(_00619_));
 sky130_vsdinv _18705_ (.A(\cpuregs[5][10] ),
    .Y(_00620_));
 sky130_vsdinv _18706_ (.A(\cpuregs[6][10] ),
    .Y(_00621_));
 sky130_vsdinv _18707_ (.A(\cpuregs[7][10] ),
    .Y(_00622_));
 sky130_vsdinv _18708_ (.A(\cpuregs[8][10] ),
    .Y(_00624_));
 sky130_vsdinv _18709_ (.A(\cpuregs[9][10] ),
    .Y(_00625_));
 sky130_vsdinv _18710_ (.A(\cpuregs[10][10] ),
    .Y(_00626_));
 sky130_vsdinv _18711_ (.A(\cpuregs[11][10] ),
    .Y(_00627_));
 sky130_vsdinv _18712_ (.A(\cpuregs[12][10] ),
    .Y(_00629_));
 sky130_vsdinv _18713_ (.A(\cpuregs[13][10] ),
    .Y(_00630_));
 sky130_vsdinv _18714_ (.A(\cpuregs[14][10] ),
    .Y(_00631_));
 sky130_vsdinv _18715_ (.A(\cpuregs[15][10] ),
    .Y(_00632_));
 sky130_vsdinv _18716_ (.A(\cpuregs[16][10] ),
    .Y(_00635_));
 sky130_vsdinv _18717_ (.A(\cpuregs[17][10] ),
    .Y(_00636_));
 sky130_vsdinv _18718_ (.A(\cpuregs[18][10] ),
    .Y(_00637_));
 sky130_vsdinv _18719_ (.A(\cpuregs[19][10] ),
    .Y(_00638_));
 sky130_vsdinv _18720_ (.A(\cpuregs[0][11] ),
    .Y(_00641_));
 sky130_vsdinv _18721_ (.A(\cpuregs[1][11] ),
    .Y(_00642_));
 sky130_vsdinv _18722_ (.A(\cpuregs[2][11] ),
    .Y(_00643_));
 sky130_vsdinv _18723_ (.A(\cpuregs[3][11] ),
    .Y(_00644_));
 sky130_vsdinv _18724_ (.A(\cpuregs[4][11] ),
    .Y(_00646_));
 sky130_vsdinv _18725_ (.A(\cpuregs[5][11] ),
    .Y(_00647_));
 sky130_vsdinv _18726_ (.A(\cpuregs[6][11] ),
    .Y(_00648_));
 sky130_vsdinv _18727_ (.A(\cpuregs[7][11] ),
    .Y(_00649_));
 sky130_vsdinv _18728_ (.A(\cpuregs[8][11] ),
    .Y(_00651_));
 sky130_vsdinv _18729_ (.A(\cpuregs[9][11] ),
    .Y(_00652_));
 sky130_vsdinv _18730_ (.A(\cpuregs[10][11] ),
    .Y(_00653_));
 sky130_vsdinv _18731_ (.A(\cpuregs[11][11] ),
    .Y(_00654_));
 sky130_vsdinv _18732_ (.A(\cpuregs[12][11] ),
    .Y(_00656_));
 sky130_vsdinv _18733_ (.A(\cpuregs[13][11] ),
    .Y(_00657_));
 sky130_vsdinv _18734_ (.A(\cpuregs[14][11] ),
    .Y(_00658_));
 sky130_vsdinv _18735_ (.A(\cpuregs[15][11] ),
    .Y(_00659_));
 sky130_vsdinv _18736_ (.A(\cpuregs[16][11] ),
    .Y(_00662_));
 sky130_vsdinv _18737_ (.A(\cpuregs[17][11] ),
    .Y(_00663_));
 sky130_vsdinv _18738_ (.A(\cpuregs[18][11] ),
    .Y(_00664_));
 sky130_vsdinv _18739_ (.A(\cpuregs[19][11] ),
    .Y(_00665_));
 sky130_vsdinv _18740_ (.A(\cpuregs[0][12] ),
    .Y(_00668_));
 sky130_vsdinv _18741_ (.A(\cpuregs[1][12] ),
    .Y(_00669_));
 sky130_vsdinv _18742_ (.A(\cpuregs[2][12] ),
    .Y(_00670_));
 sky130_vsdinv _18743_ (.A(\cpuregs[3][12] ),
    .Y(_00671_));
 sky130_vsdinv _18744_ (.A(\cpuregs[4][12] ),
    .Y(_00673_));
 sky130_vsdinv _18745_ (.A(\cpuregs[5][12] ),
    .Y(_00674_));
 sky130_vsdinv _18746_ (.A(\cpuregs[6][12] ),
    .Y(_00675_));
 sky130_vsdinv _18747_ (.A(\cpuregs[7][12] ),
    .Y(_00676_));
 sky130_vsdinv _18748_ (.A(\cpuregs[8][12] ),
    .Y(_00678_));
 sky130_vsdinv _18749_ (.A(\cpuregs[9][12] ),
    .Y(_00679_));
 sky130_vsdinv _18750_ (.A(\cpuregs[10][12] ),
    .Y(_00680_));
 sky130_vsdinv _18751_ (.A(\cpuregs[11][12] ),
    .Y(_00681_));
 sky130_vsdinv _18752_ (.A(\cpuregs[12][12] ),
    .Y(_00683_));
 sky130_vsdinv _18753_ (.A(\cpuregs[13][12] ),
    .Y(_00684_));
 sky130_vsdinv _18754_ (.A(\cpuregs[14][12] ),
    .Y(_00685_));
 sky130_vsdinv _18755_ (.A(\cpuregs[15][12] ),
    .Y(_00686_));
 sky130_vsdinv _18756_ (.A(\cpuregs[16][12] ),
    .Y(_00689_));
 sky130_vsdinv _18757_ (.A(\cpuregs[17][12] ),
    .Y(_00690_));
 sky130_vsdinv _18758_ (.A(\cpuregs[18][12] ),
    .Y(_00691_));
 sky130_vsdinv _18759_ (.A(\cpuregs[19][12] ),
    .Y(_00692_));
 sky130_vsdinv _18760_ (.A(\cpuregs[0][13] ),
    .Y(_00695_));
 sky130_vsdinv _18761_ (.A(\cpuregs[1][13] ),
    .Y(_00696_));
 sky130_vsdinv _18762_ (.A(\cpuregs[2][13] ),
    .Y(_00697_));
 sky130_vsdinv _18763_ (.A(\cpuregs[3][13] ),
    .Y(_00698_));
 sky130_vsdinv _18764_ (.A(\cpuregs[4][13] ),
    .Y(_00700_));
 sky130_vsdinv _18765_ (.A(\cpuregs[5][13] ),
    .Y(_00701_));
 sky130_vsdinv _18766_ (.A(\cpuregs[6][13] ),
    .Y(_00702_));
 sky130_vsdinv _18767_ (.A(\cpuregs[7][13] ),
    .Y(_00703_));
 sky130_vsdinv _18768_ (.A(\cpuregs[8][13] ),
    .Y(_00705_));
 sky130_vsdinv _18769_ (.A(\cpuregs[9][13] ),
    .Y(_00706_));
 sky130_vsdinv _18770_ (.A(\cpuregs[10][13] ),
    .Y(_00707_));
 sky130_vsdinv _18771_ (.A(\cpuregs[11][13] ),
    .Y(_00708_));
 sky130_vsdinv _18772_ (.A(\cpuregs[12][13] ),
    .Y(_00710_));
 sky130_vsdinv _18773_ (.A(\cpuregs[13][13] ),
    .Y(_00711_));
 sky130_vsdinv _18774_ (.A(\cpuregs[14][13] ),
    .Y(_00712_));
 sky130_vsdinv _18775_ (.A(\cpuregs[15][13] ),
    .Y(_00713_));
 sky130_vsdinv _18776_ (.A(\cpuregs[16][13] ),
    .Y(_00716_));
 sky130_vsdinv _18777_ (.A(\cpuregs[17][13] ),
    .Y(_00717_));
 sky130_vsdinv _18778_ (.A(\cpuregs[18][13] ),
    .Y(_00718_));
 sky130_vsdinv _18779_ (.A(\cpuregs[19][13] ),
    .Y(_00719_));
 sky130_vsdinv _18780_ (.A(\cpuregs[0][14] ),
    .Y(_00722_));
 sky130_vsdinv _18781_ (.A(\cpuregs[1][14] ),
    .Y(_00723_));
 sky130_vsdinv _18782_ (.A(\cpuregs[2][14] ),
    .Y(_00724_));
 sky130_vsdinv _18783_ (.A(\cpuregs[3][14] ),
    .Y(_00725_));
 sky130_vsdinv _18784_ (.A(\cpuregs[4][14] ),
    .Y(_00727_));
 sky130_vsdinv _18785_ (.A(\cpuregs[5][14] ),
    .Y(_00728_));
 sky130_vsdinv _18786_ (.A(\cpuregs[6][14] ),
    .Y(_00729_));
 sky130_vsdinv _18787_ (.A(\cpuregs[7][14] ),
    .Y(_00730_));
 sky130_vsdinv _18788_ (.A(\cpuregs[8][14] ),
    .Y(_00732_));
 sky130_vsdinv _18789_ (.A(\cpuregs[9][14] ),
    .Y(_00733_));
 sky130_vsdinv _18790_ (.A(\cpuregs[10][14] ),
    .Y(_00734_));
 sky130_vsdinv _18791_ (.A(\cpuregs[11][14] ),
    .Y(_00735_));
 sky130_vsdinv _18792_ (.A(\cpuregs[12][14] ),
    .Y(_00737_));
 sky130_vsdinv _18793_ (.A(\cpuregs[13][14] ),
    .Y(_00738_));
 sky130_vsdinv _18794_ (.A(\cpuregs[14][14] ),
    .Y(_00739_));
 sky130_vsdinv _18795_ (.A(\cpuregs[15][14] ),
    .Y(_00740_));
 sky130_vsdinv _18796_ (.A(\cpuregs[16][14] ),
    .Y(_00743_));
 sky130_vsdinv _18797_ (.A(\cpuregs[17][14] ),
    .Y(_00744_));
 sky130_vsdinv _18798_ (.A(\cpuregs[18][14] ),
    .Y(_00745_));
 sky130_vsdinv _18799_ (.A(\cpuregs[19][14] ),
    .Y(_00746_));
 sky130_vsdinv _18800_ (.A(\cpuregs[0][15] ),
    .Y(_00749_));
 sky130_vsdinv _18801_ (.A(\cpuregs[1][15] ),
    .Y(_00750_));
 sky130_vsdinv _18802_ (.A(\cpuregs[2][15] ),
    .Y(_00751_));
 sky130_vsdinv _18803_ (.A(\cpuregs[3][15] ),
    .Y(_00752_));
 sky130_vsdinv _18804_ (.A(\cpuregs[4][15] ),
    .Y(_00754_));
 sky130_vsdinv _18805_ (.A(\cpuregs[5][15] ),
    .Y(_00755_));
 sky130_vsdinv _18806_ (.A(\cpuregs[6][15] ),
    .Y(_00756_));
 sky130_vsdinv _18807_ (.A(\cpuregs[7][15] ),
    .Y(_00757_));
 sky130_vsdinv _18808_ (.A(\cpuregs[8][15] ),
    .Y(_00759_));
 sky130_vsdinv _18809_ (.A(\cpuregs[9][15] ),
    .Y(_00760_));
 sky130_vsdinv _18810_ (.A(\cpuregs[10][15] ),
    .Y(_00761_));
 sky130_vsdinv _18811_ (.A(\cpuregs[11][15] ),
    .Y(_00762_));
 sky130_vsdinv _18812_ (.A(\cpuregs[12][15] ),
    .Y(_00764_));
 sky130_vsdinv _18813_ (.A(\cpuregs[13][15] ),
    .Y(_00765_));
 sky130_vsdinv _18814_ (.A(\cpuregs[14][15] ),
    .Y(_00766_));
 sky130_vsdinv _18815_ (.A(\cpuregs[15][15] ),
    .Y(_00767_));
 sky130_vsdinv _18816_ (.A(\cpuregs[16][15] ),
    .Y(_00770_));
 sky130_vsdinv _18817_ (.A(\cpuregs[17][15] ),
    .Y(_00771_));
 sky130_vsdinv _18818_ (.A(\cpuregs[18][15] ),
    .Y(_00772_));
 sky130_vsdinv _18819_ (.A(\cpuregs[19][15] ),
    .Y(_00773_));
 sky130_vsdinv _18820_ (.A(\cpuregs[0][16] ),
    .Y(_00776_));
 sky130_vsdinv _18821_ (.A(\cpuregs[1][16] ),
    .Y(_00777_));
 sky130_vsdinv _18822_ (.A(\cpuregs[2][16] ),
    .Y(_00778_));
 sky130_vsdinv _18823_ (.A(\cpuregs[3][16] ),
    .Y(_00779_));
 sky130_vsdinv _18824_ (.A(\cpuregs[4][16] ),
    .Y(_00781_));
 sky130_vsdinv _18825_ (.A(\cpuregs[5][16] ),
    .Y(_00782_));
 sky130_vsdinv _18826_ (.A(\cpuregs[6][16] ),
    .Y(_00783_));
 sky130_vsdinv _18827_ (.A(\cpuregs[7][16] ),
    .Y(_00784_));
 sky130_vsdinv _18828_ (.A(\cpuregs[8][16] ),
    .Y(_00786_));
 sky130_vsdinv _18829_ (.A(\cpuregs[9][16] ),
    .Y(_00787_));
 sky130_vsdinv _18830_ (.A(\cpuregs[10][16] ),
    .Y(_00788_));
 sky130_vsdinv _18831_ (.A(\cpuregs[11][16] ),
    .Y(_00789_));
 sky130_vsdinv _18832_ (.A(\cpuregs[12][16] ),
    .Y(_00791_));
 sky130_vsdinv _18833_ (.A(\cpuregs[13][16] ),
    .Y(_00792_));
 sky130_vsdinv _18834_ (.A(\cpuregs[14][16] ),
    .Y(_00793_));
 sky130_vsdinv _18835_ (.A(\cpuregs[15][16] ),
    .Y(_00794_));
 sky130_vsdinv _18836_ (.A(\cpuregs[16][16] ),
    .Y(_00797_));
 sky130_vsdinv _18837_ (.A(\cpuregs[17][16] ),
    .Y(_00798_));
 sky130_vsdinv _18838_ (.A(\cpuregs[18][16] ),
    .Y(_00799_));
 sky130_vsdinv _18839_ (.A(\cpuregs[19][16] ),
    .Y(_00800_));
 sky130_vsdinv _18840_ (.A(\cpuregs[0][17] ),
    .Y(_00803_));
 sky130_vsdinv _18841_ (.A(\cpuregs[1][17] ),
    .Y(_00804_));
 sky130_vsdinv _18842_ (.A(\cpuregs[2][17] ),
    .Y(_00805_));
 sky130_vsdinv _18843_ (.A(\cpuregs[3][17] ),
    .Y(_00806_));
 sky130_vsdinv _18844_ (.A(\cpuregs[4][17] ),
    .Y(_00808_));
 sky130_vsdinv _18845_ (.A(\cpuregs[5][17] ),
    .Y(_00809_));
 sky130_vsdinv _18846_ (.A(\cpuregs[6][17] ),
    .Y(_00810_));
 sky130_vsdinv _18847_ (.A(\cpuregs[7][17] ),
    .Y(_00811_));
 sky130_vsdinv _18848_ (.A(\cpuregs[8][17] ),
    .Y(_00813_));
 sky130_vsdinv _18849_ (.A(\cpuregs[9][17] ),
    .Y(_00814_));
 sky130_vsdinv _18850_ (.A(\cpuregs[10][17] ),
    .Y(_00815_));
 sky130_vsdinv _18851_ (.A(\cpuregs[11][17] ),
    .Y(_00816_));
 sky130_vsdinv _18852_ (.A(\cpuregs[12][17] ),
    .Y(_00818_));
 sky130_vsdinv _18853_ (.A(\cpuregs[13][17] ),
    .Y(_00819_));
 sky130_vsdinv _18854_ (.A(\cpuregs[14][17] ),
    .Y(_00820_));
 sky130_vsdinv _18855_ (.A(\cpuregs[15][17] ),
    .Y(_00821_));
 sky130_vsdinv _18856_ (.A(\cpuregs[16][17] ),
    .Y(_00824_));
 sky130_vsdinv _18857_ (.A(\cpuregs[17][17] ),
    .Y(_00825_));
 sky130_vsdinv _18858_ (.A(\cpuregs[18][17] ),
    .Y(_00826_));
 sky130_vsdinv _18859_ (.A(\cpuregs[19][17] ),
    .Y(_00827_));
 sky130_vsdinv _18860_ (.A(\cpuregs[0][18] ),
    .Y(_00830_));
 sky130_vsdinv _18861_ (.A(\cpuregs[1][18] ),
    .Y(_00831_));
 sky130_vsdinv _18862_ (.A(\cpuregs[2][18] ),
    .Y(_00832_));
 sky130_vsdinv _18863_ (.A(\cpuregs[3][18] ),
    .Y(_00833_));
 sky130_vsdinv _18864_ (.A(\cpuregs[4][18] ),
    .Y(_00835_));
 sky130_vsdinv _18865_ (.A(\cpuregs[5][18] ),
    .Y(_00836_));
 sky130_vsdinv _18866_ (.A(\cpuregs[6][18] ),
    .Y(_00837_));
 sky130_vsdinv _18867_ (.A(\cpuregs[7][18] ),
    .Y(_00838_));
 sky130_vsdinv _18868_ (.A(\cpuregs[8][18] ),
    .Y(_00840_));
 sky130_vsdinv _18869_ (.A(\cpuregs[9][18] ),
    .Y(_00841_));
 sky130_vsdinv _18870_ (.A(\cpuregs[10][18] ),
    .Y(_00842_));
 sky130_vsdinv _18871_ (.A(\cpuregs[11][18] ),
    .Y(_00843_));
 sky130_vsdinv _18872_ (.A(\cpuregs[12][18] ),
    .Y(_00845_));
 sky130_vsdinv _18873_ (.A(\cpuregs[13][18] ),
    .Y(_00846_));
 sky130_vsdinv _18874_ (.A(\cpuregs[14][18] ),
    .Y(_00847_));
 sky130_vsdinv _18875_ (.A(\cpuregs[15][18] ),
    .Y(_00848_));
 sky130_vsdinv _18876_ (.A(\cpuregs[16][18] ),
    .Y(_00851_));
 sky130_vsdinv _18877_ (.A(\cpuregs[17][18] ),
    .Y(_00852_));
 sky130_vsdinv _18878_ (.A(\cpuregs[18][18] ),
    .Y(_00853_));
 sky130_vsdinv _18879_ (.A(\cpuregs[19][18] ),
    .Y(_00854_));
 sky130_vsdinv _18880_ (.A(\cpuregs[0][19] ),
    .Y(_00857_));
 sky130_vsdinv _18881_ (.A(\cpuregs[1][19] ),
    .Y(_00858_));
 sky130_vsdinv _18882_ (.A(\cpuregs[2][19] ),
    .Y(_00859_));
 sky130_vsdinv _18883_ (.A(\cpuregs[3][19] ),
    .Y(_00860_));
 sky130_vsdinv _18884_ (.A(\cpuregs[4][19] ),
    .Y(_00862_));
 sky130_vsdinv _18885_ (.A(\cpuregs[5][19] ),
    .Y(_00863_));
 sky130_vsdinv _18886_ (.A(\cpuregs[6][19] ),
    .Y(_00864_));
 sky130_vsdinv _18887_ (.A(\cpuregs[7][19] ),
    .Y(_00865_));
 sky130_vsdinv _18888_ (.A(\cpuregs[8][19] ),
    .Y(_00867_));
 sky130_vsdinv _18889_ (.A(\cpuregs[9][19] ),
    .Y(_00868_));
 sky130_vsdinv _18890_ (.A(\cpuregs[10][19] ),
    .Y(_00869_));
 sky130_vsdinv _18891_ (.A(\cpuregs[11][19] ),
    .Y(_00870_));
 sky130_vsdinv _18892_ (.A(\cpuregs[12][19] ),
    .Y(_00872_));
 sky130_vsdinv _18893_ (.A(\cpuregs[13][19] ),
    .Y(_00873_));
 sky130_vsdinv _18894_ (.A(\cpuregs[14][19] ),
    .Y(_00874_));
 sky130_vsdinv _18895_ (.A(\cpuregs[15][19] ),
    .Y(_00875_));
 sky130_vsdinv _18896_ (.A(\cpuregs[16][19] ),
    .Y(_00878_));
 sky130_vsdinv _18897_ (.A(\cpuregs[17][19] ),
    .Y(_00879_));
 sky130_vsdinv _18898_ (.A(\cpuregs[18][19] ),
    .Y(_00880_));
 sky130_vsdinv _18899_ (.A(\cpuregs[19][19] ),
    .Y(_00881_));
 sky130_vsdinv _18900_ (.A(\cpuregs[0][20] ),
    .Y(_00884_));
 sky130_vsdinv _18901_ (.A(\cpuregs[1][20] ),
    .Y(_00885_));
 sky130_vsdinv _18902_ (.A(\cpuregs[2][20] ),
    .Y(_00886_));
 sky130_vsdinv _18903_ (.A(\cpuregs[3][20] ),
    .Y(_00887_));
 sky130_vsdinv _18904_ (.A(\cpuregs[4][20] ),
    .Y(_00889_));
 sky130_vsdinv _18905_ (.A(\cpuregs[5][20] ),
    .Y(_00890_));
 sky130_vsdinv _18906_ (.A(\cpuregs[6][20] ),
    .Y(_00891_));
 sky130_vsdinv _18907_ (.A(\cpuregs[7][20] ),
    .Y(_00892_));
 sky130_vsdinv _18908_ (.A(\cpuregs[8][20] ),
    .Y(_00894_));
 sky130_vsdinv _18909_ (.A(\cpuregs[9][20] ),
    .Y(_00895_));
 sky130_vsdinv _18910_ (.A(\cpuregs[10][20] ),
    .Y(_00896_));
 sky130_vsdinv _18911_ (.A(\cpuregs[11][20] ),
    .Y(_00897_));
 sky130_vsdinv _18912_ (.A(\cpuregs[12][20] ),
    .Y(_00899_));
 sky130_vsdinv _18913_ (.A(\cpuregs[13][20] ),
    .Y(_00900_));
 sky130_vsdinv _18914_ (.A(\cpuregs[14][20] ),
    .Y(_00901_));
 sky130_vsdinv _18915_ (.A(\cpuregs[15][20] ),
    .Y(_00902_));
 sky130_vsdinv _18916_ (.A(\cpuregs[16][20] ),
    .Y(_00905_));
 sky130_vsdinv _18917_ (.A(\cpuregs[17][20] ),
    .Y(_00906_));
 sky130_vsdinv _18918_ (.A(\cpuregs[18][20] ),
    .Y(_00907_));
 sky130_vsdinv _18919_ (.A(\cpuregs[19][20] ),
    .Y(_00908_));
 sky130_vsdinv _18920_ (.A(\cpuregs[0][21] ),
    .Y(_00911_));
 sky130_vsdinv _18921_ (.A(\cpuregs[1][21] ),
    .Y(_00912_));
 sky130_vsdinv _18922_ (.A(\cpuregs[2][21] ),
    .Y(_00913_));
 sky130_vsdinv _18923_ (.A(\cpuregs[3][21] ),
    .Y(_00914_));
 sky130_vsdinv _18924_ (.A(\cpuregs[4][21] ),
    .Y(_00916_));
 sky130_vsdinv _18925_ (.A(\cpuregs[5][21] ),
    .Y(_00917_));
 sky130_vsdinv _18926_ (.A(\cpuregs[6][21] ),
    .Y(_00918_));
 sky130_vsdinv _18927_ (.A(\cpuregs[7][21] ),
    .Y(_00919_));
 sky130_vsdinv _18928_ (.A(\cpuregs[8][21] ),
    .Y(_00921_));
 sky130_vsdinv _18929_ (.A(\cpuregs[9][21] ),
    .Y(_00922_));
 sky130_vsdinv _18930_ (.A(\cpuregs[10][21] ),
    .Y(_00923_));
 sky130_vsdinv _18931_ (.A(\cpuregs[11][21] ),
    .Y(_00924_));
 sky130_vsdinv _18932_ (.A(\cpuregs[12][21] ),
    .Y(_00926_));
 sky130_vsdinv _18933_ (.A(\cpuregs[13][21] ),
    .Y(_00927_));
 sky130_vsdinv _18934_ (.A(\cpuregs[14][21] ),
    .Y(_00928_));
 sky130_vsdinv _18935_ (.A(\cpuregs[15][21] ),
    .Y(_00929_));
 sky130_vsdinv _18936_ (.A(\cpuregs[16][21] ),
    .Y(_00932_));
 sky130_vsdinv _18937_ (.A(\cpuregs[17][21] ),
    .Y(_00933_));
 sky130_vsdinv _18938_ (.A(\cpuregs[18][21] ),
    .Y(_00934_));
 sky130_vsdinv _18939_ (.A(\cpuregs[19][21] ),
    .Y(_00935_));
 sky130_vsdinv _18940_ (.A(\cpuregs[0][22] ),
    .Y(_00938_));
 sky130_vsdinv _18941_ (.A(\cpuregs[1][22] ),
    .Y(_00939_));
 sky130_vsdinv _18942_ (.A(\cpuregs[2][22] ),
    .Y(_00940_));
 sky130_vsdinv _18943_ (.A(\cpuregs[3][22] ),
    .Y(_00941_));
 sky130_vsdinv _18944_ (.A(\cpuregs[4][22] ),
    .Y(_00943_));
 sky130_vsdinv _18945_ (.A(\cpuregs[5][22] ),
    .Y(_00944_));
 sky130_vsdinv _18946_ (.A(\cpuregs[6][22] ),
    .Y(_00945_));
 sky130_vsdinv _18947_ (.A(\cpuregs[7][22] ),
    .Y(_00946_));
 sky130_fd_sc_hd__o32a_1 _18948_ (.A1(_13351_),
    .A2(_14057_),
    .A3(_12010_),
    .B1(_13360_),
    .B2(_12014_),
    .X(_14162_));
 sky130_fd_sc_hd__or2_1 _18949_ (.A(_12009_),
    .B(_14162_),
    .X(_14163_));
 sky130_fd_sc_hd__o221ai_1 _18950_ (.A1(_12545_),
    .A2(_00322_),
    .B1(_13988_),
    .B2(_14151_),
    .C1(_14163_),
    .Y(_00045_));
 sky130_vsdinv _18951_ (.A(\cpuregs[8][22] ),
    .Y(_00948_));
 sky130_vsdinv _18952_ (.A(\cpuregs[9][22] ),
    .Y(_00949_));
 sky130_vsdinv _18953_ (.A(\cpuregs[10][22] ),
    .Y(_00950_));
 sky130_vsdinv _18954_ (.A(\cpuregs[11][22] ),
    .Y(_00951_));
 sky130_vsdinv _18955_ (.A(\cpuregs[12][22] ),
    .Y(_00953_));
 sky130_vsdinv _18956_ (.A(\cpuregs[13][22] ),
    .Y(_00954_));
 sky130_vsdinv _18957_ (.A(\cpuregs[14][22] ),
    .Y(_00955_));
 sky130_vsdinv _18958_ (.A(\cpuregs[15][22] ),
    .Y(_00956_));
 sky130_vsdinv _18959_ (.A(\cpuregs[16][22] ),
    .Y(_00959_));
 sky130_vsdinv _18960_ (.A(\cpuregs[17][22] ),
    .Y(_00960_));
 sky130_vsdinv _18961_ (.A(\cpuregs[18][22] ),
    .Y(_00961_));
 sky130_vsdinv _18962_ (.A(\cpuregs[19][22] ),
    .Y(_00962_));
 sky130_vsdinv _18963_ (.A(\cpuregs[0][23] ),
    .Y(_00965_));
 sky130_vsdinv _18964_ (.A(\cpuregs[1][23] ),
    .Y(_00966_));
 sky130_vsdinv _18965_ (.A(\cpuregs[2][23] ),
    .Y(_00967_));
 sky130_vsdinv _18966_ (.A(\cpuregs[3][23] ),
    .Y(_00968_));
 sky130_vsdinv _18967_ (.A(\cpuregs[4][23] ),
    .Y(_00970_));
 sky130_vsdinv _18968_ (.A(\cpuregs[5][23] ),
    .Y(_00971_));
 sky130_vsdinv _18969_ (.A(\cpuregs[6][23] ),
    .Y(_00972_));
 sky130_vsdinv _18970_ (.A(\cpuregs[7][23] ),
    .Y(_00973_));
 sky130_vsdinv _18971_ (.A(\cpuregs[8][23] ),
    .Y(_00975_));
 sky130_vsdinv _18972_ (.A(\cpuregs[9][23] ),
    .Y(_00976_));
 sky130_vsdinv _18973_ (.A(\cpuregs[10][23] ),
    .Y(_00977_));
 sky130_vsdinv _18974_ (.A(\cpuregs[11][23] ),
    .Y(_00978_));
 sky130_vsdinv _18975_ (.A(\cpuregs[12][23] ),
    .Y(_00980_));
 sky130_vsdinv _18976_ (.A(\cpuregs[13][23] ),
    .Y(_00981_));
 sky130_vsdinv _18977_ (.A(\cpuregs[14][23] ),
    .Y(_00982_));
 sky130_vsdinv _18978_ (.A(\cpuregs[15][23] ),
    .Y(_00983_));
 sky130_vsdinv _18979_ (.A(\cpuregs[16][23] ),
    .Y(_00986_));
 sky130_vsdinv _18980_ (.A(\cpuregs[17][23] ),
    .Y(_00987_));
 sky130_vsdinv _18981_ (.A(\cpuregs[18][23] ),
    .Y(_00988_));
 sky130_vsdinv _18982_ (.A(\cpuregs[19][23] ),
    .Y(_00989_));
 sky130_vsdinv _18983_ (.A(\cpuregs[0][24] ),
    .Y(_00992_));
 sky130_vsdinv _18984_ (.A(\cpuregs[1][24] ),
    .Y(_00993_));
 sky130_vsdinv _18985_ (.A(\cpuregs[2][24] ),
    .Y(_00994_));
 sky130_vsdinv _18986_ (.A(\cpuregs[3][24] ),
    .Y(_00995_));
 sky130_vsdinv _18987_ (.A(\cpuregs[4][24] ),
    .Y(_00997_));
 sky130_vsdinv _18988_ (.A(\cpuregs[5][24] ),
    .Y(_00998_));
 sky130_vsdinv _18989_ (.A(\cpuregs[6][24] ),
    .Y(_00999_));
 sky130_vsdinv _18990_ (.A(\cpuregs[7][24] ),
    .Y(_01000_));
 sky130_vsdinv _18991_ (.A(\cpuregs[8][24] ),
    .Y(_01002_));
 sky130_vsdinv _18992_ (.A(\cpuregs[9][24] ),
    .Y(_01003_));
 sky130_vsdinv _18993_ (.A(\cpuregs[10][24] ),
    .Y(_01004_));
 sky130_vsdinv _18994_ (.A(\cpuregs[11][24] ),
    .Y(_01005_));
 sky130_vsdinv _18995_ (.A(\cpuregs[12][24] ),
    .Y(_01007_));
 sky130_vsdinv _18996_ (.A(\cpuregs[13][24] ),
    .Y(_01008_));
 sky130_vsdinv _18997_ (.A(\cpuregs[14][24] ),
    .Y(_01009_));
 sky130_vsdinv _18998_ (.A(\cpuregs[15][24] ),
    .Y(_01010_));
 sky130_vsdinv _18999_ (.A(\cpuregs[16][24] ),
    .Y(_01013_));
 sky130_vsdinv _19000_ (.A(\cpuregs[17][24] ),
    .Y(_01014_));
 sky130_vsdinv _19001_ (.A(\cpuregs[18][24] ),
    .Y(_01015_));
 sky130_vsdinv _19002_ (.A(\cpuregs[19][24] ),
    .Y(_01016_));
 sky130_vsdinv _19003_ (.A(\cpuregs[0][25] ),
    .Y(_01019_));
 sky130_vsdinv _19004_ (.A(\cpuregs[1][25] ),
    .Y(_01020_));
 sky130_vsdinv _19005_ (.A(\cpuregs[2][25] ),
    .Y(_01021_));
 sky130_vsdinv _19006_ (.A(\cpuregs[3][25] ),
    .Y(_01022_));
 sky130_vsdinv _19007_ (.A(\cpuregs[4][25] ),
    .Y(_01024_));
 sky130_vsdinv _19008_ (.A(\cpuregs[5][25] ),
    .Y(_01025_));
 sky130_vsdinv _19009_ (.A(\cpuregs[6][25] ),
    .Y(_01026_));
 sky130_vsdinv _19010_ (.A(\cpuregs[7][25] ),
    .Y(_01027_));
 sky130_fd_sc_hd__nor2_2 _19011_ (.A(\mem_state[1] ),
    .B(_11549_),
    .Y(_00289_));
 sky130_fd_sc_hd__nand2_1 _19012_ (.A(_13184_),
    .B(_00289_),
    .Y(_00298_));
 sky130_vsdinv _19013_ (.A(\cpuregs[8][25] ),
    .Y(_01029_));
 sky130_vsdinv _19014_ (.A(\cpuregs[9][25] ),
    .Y(_01030_));
 sky130_vsdinv _19015_ (.A(\cpuregs[10][25] ),
    .Y(_01031_));
 sky130_vsdinv _19016_ (.A(\cpuregs[11][25] ),
    .Y(_01032_));
 sky130_vsdinv _19017_ (.A(\cpuregs[12][25] ),
    .Y(_01034_));
 sky130_vsdinv _19018_ (.A(\cpuregs[13][25] ),
    .Y(_01035_));
 sky130_vsdinv _19019_ (.A(\cpuregs[14][25] ),
    .Y(_01036_));
 sky130_vsdinv _19020_ (.A(\cpuregs[15][25] ),
    .Y(_01037_));
 sky130_vsdinv _19021_ (.A(\cpuregs[16][25] ),
    .Y(_01040_));
 sky130_vsdinv _19022_ (.A(\cpuregs[17][25] ),
    .Y(_01041_));
 sky130_vsdinv _19023_ (.A(\cpuregs[18][25] ),
    .Y(_01042_));
 sky130_vsdinv _19024_ (.A(\cpuregs[19][25] ),
    .Y(_01043_));
 sky130_vsdinv _19025_ (.A(\cpuregs[0][26] ),
    .Y(_01046_));
 sky130_vsdinv _19026_ (.A(\cpuregs[1][26] ),
    .Y(_01047_));
 sky130_vsdinv _19027_ (.A(\cpuregs[2][26] ),
    .Y(_01048_));
 sky130_vsdinv _19028_ (.A(\cpuregs[3][26] ),
    .Y(_01049_));
 sky130_vsdinv _19029_ (.A(\cpuregs[4][26] ),
    .Y(_01051_));
 sky130_vsdinv _19030_ (.A(\cpuregs[5][26] ),
    .Y(_01052_));
 sky130_vsdinv _19031_ (.A(\cpuregs[6][26] ),
    .Y(_01053_));
 sky130_vsdinv _19032_ (.A(\cpuregs[7][26] ),
    .Y(_01054_));
 sky130_vsdinv _19033_ (.A(\cpuregs[8][26] ),
    .Y(_01056_));
 sky130_vsdinv _19034_ (.A(\cpuregs[9][26] ),
    .Y(_01057_));
 sky130_vsdinv _19035_ (.A(\cpuregs[10][26] ),
    .Y(_01058_));
 sky130_vsdinv _19036_ (.A(\cpuregs[11][26] ),
    .Y(_01059_));
 sky130_vsdinv _19037_ (.A(\cpuregs[12][26] ),
    .Y(_01061_));
 sky130_vsdinv _19038_ (.A(\cpuregs[13][26] ),
    .Y(_01062_));
 sky130_vsdinv _19039_ (.A(\cpuregs[14][26] ),
    .Y(_01063_));
 sky130_vsdinv _19040_ (.A(\cpuregs[15][26] ),
    .Y(_01064_));
 sky130_vsdinv _19041_ (.A(\cpuregs[16][26] ),
    .Y(_01067_));
 sky130_vsdinv _19042_ (.A(\cpuregs[17][26] ),
    .Y(_01068_));
 sky130_vsdinv _19043_ (.A(\cpuregs[18][26] ),
    .Y(_01069_));
 sky130_vsdinv _19044_ (.A(\cpuregs[19][26] ),
    .Y(_01070_));
 sky130_vsdinv _19045_ (.A(\mem_wordsize[1] ),
    .Y(_14164_));
 sky130_fd_sc_hd__clkbuf_2 _19046_ (.A(_14164_),
    .X(_14165_));
 sky130_fd_sc_hd__o211a_1 _19047_ (.A1(instr_lbu),
    .A2(instr_lb),
    .B1(_12012_),
    .C1(_11563_),
    .X(_14166_));
 sky130_fd_sc_hd__a31oi_2 _19048_ (.A1(_00291_),
    .A2(instr_sb),
    .A3(\cpu_state[5] ),
    .B1(_14166_),
    .Y(_14167_));
 sky130_fd_sc_hd__o22ai_1 _19049_ (.A1(_14165_),
    .A2(_14151_),
    .B1(_14044_),
    .B2(_14167_),
    .Y(_00046_));
 sky130_vsdinv _19050_ (.A(\cpuregs[0][27] ),
    .Y(_01073_));
 sky130_vsdinv _19051_ (.A(\cpuregs[1][27] ),
    .Y(_01074_));
 sky130_vsdinv _19052_ (.A(\cpuregs[2][27] ),
    .Y(_01075_));
 sky130_vsdinv _19053_ (.A(\cpuregs[3][27] ),
    .Y(_01076_));
 sky130_vsdinv _19054_ (.A(\cpuregs[4][27] ),
    .Y(_01078_));
 sky130_vsdinv _19055_ (.A(\cpuregs[5][27] ),
    .Y(_01079_));
 sky130_vsdinv _19056_ (.A(\cpuregs[6][27] ),
    .Y(_01080_));
 sky130_vsdinv _19057_ (.A(\cpuregs[7][27] ),
    .Y(_01081_));
 sky130_vsdinv _19058_ (.A(\cpuregs[8][27] ),
    .Y(_01083_));
 sky130_vsdinv _19059_ (.A(\cpuregs[9][27] ),
    .Y(_01084_));
 sky130_vsdinv _19060_ (.A(\cpuregs[10][27] ),
    .Y(_01085_));
 sky130_vsdinv _19061_ (.A(\cpuregs[11][27] ),
    .Y(_01086_));
 sky130_vsdinv _19062_ (.A(\cpuregs[12][27] ),
    .Y(_01088_));
 sky130_vsdinv _19063_ (.A(\cpuregs[13][27] ),
    .Y(_01089_));
 sky130_vsdinv _19064_ (.A(\cpuregs[14][27] ),
    .Y(_01090_));
 sky130_vsdinv _19065_ (.A(\cpuregs[15][27] ),
    .Y(_01091_));
 sky130_vsdinv _19066_ (.A(\cpuregs[16][27] ),
    .Y(_01094_));
 sky130_vsdinv _19067_ (.A(\cpuregs[17][27] ),
    .Y(_01095_));
 sky130_vsdinv _19068_ (.A(\cpuregs[18][27] ),
    .Y(_01096_));
 sky130_vsdinv _19069_ (.A(\cpuregs[19][27] ),
    .Y(_01097_));
 sky130_vsdinv _19070_ (.A(\cpuregs[0][28] ),
    .Y(_01100_));
 sky130_vsdinv _19071_ (.A(\cpuregs[1][28] ),
    .Y(_01101_));
 sky130_vsdinv _19072_ (.A(\cpuregs[2][28] ),
    .Y(_01102_));
 sky130_vsdinv _19073_ (.A(\cpuregs[3][28] ),
    .Y(_01103_));
 sky130_vsdinv _19074_ (.A(\cpuregs[4][28] ),
    .Y(_01105_));
 sky130_vsdinv _19075_ (.A(\cpuregs[5][28] ),
    .Y(_01106_));
 sky130_vsdinv _19076_ (.A(\cpuregs[6][28] ),
    .Y(_01107_));
 sky130_vsdinv _19077_ (.A(\cpuregs[7][28] ),
    .Y(_01108_));
 sky130_vsdinv _19078_ (.A(\cpuregs[8][28] ),
    .Y(_01110_));
 sky130_vsdinv _19079_ (.A(\cpuregs[9][28] ),
    .Y(_01111_));
 sky130_vsdinv _19080_ (.A(\cpuregs[10][28] ),
    .Y(_01112_));
 sky130_vsdinv _19081_ (.A(\cpuregs[11][28] ),
    .Y(_01113_));
 sky130_vsdinv _19082_ (.A(\cpuregs[12][28] ),
    .Y(_01115_));
 sky130_vsdinv _19083_ (.A(\cpuregs[13][28] ),
    .Y(_01116_));
 sky130_vsdinv _19084_ (.A(\cpuregs[14][28] ),
    .Y(_01117_));
 sky130_vsdinv _19085_ (.A(\cpuregs[15][28] ),
    .Y(_01118_));
 sky130_vsdinv _19086_ (.A(\cpuregs[16][28] ),
    .Y(_01121_));
 sky130_vsdinv _19087_ (.A(\cpuregs[17][28] ),
    .Y(_01122_));
 sky130_vsdinv _19088_ (.A(\cpuregs[18][28] ),
    .Y(_01123_));
 sky130_vsdinv _19089_ (.A(\cpuregs[19][28] ),
    .Y(_01124_));
 sky130_vsdinv _19090_ (.A(\cpuregs[0][29] ),
    .Y(_01127_));
 sky130_vsdinv _19091_ (.A(\cpuregs[1][29] ),
    .Y(_01128_));
 sky130_vsdinv _19092_ (.A(\cpuregs[2][29] ),
    .Y(_01129_));
 sky130_vsdinv _19093_ (.A(\cpuregs[3][29] ),
    .Y(_01130_));
 sky130_vsdinv _19094_ (.A(\cpuregs[4][29] ),
    .Y(_01132_));
 sky130_vsdinv _19095_ (.A(\cpuregs[5][29] ),
    .Y(_01133_));
 sky130_vsdinv _19096_ (.A(\cpuregs[6][29] ),
    .Y(_01134_));
 sky130_vsdinv _19097_ (.A(\cpuregs[7][29] ),
    .Y(_01135_));
 sky130_vsdinv _19098_ (.A(\cpuregs[8][29] ),
    .Y(_01137_));
 sky130_vsdinv _19099_ (.A(\cpuregs[9][29] ),
    .Y(_01138_));
 sky130_vsdinv _19100_ (.A(\cpuregs[10][29] ),
    .Y(_01139_));
 sky130_vsdinv _19101_ (.A(\cpuregs[11][29] ),
    .Y(_01140_));
 sky130_vsdinv _19102_ (.A(\cpuregs[12][29] ),
    .Y(_01142_));
 sky130_vsdinv _19103_ (.A(\cpuregs[13][29] ),
    .Y(_01143_));
 sky130_fd_sc_hd__buf_1 _19104_ (.A(_13779_),
    .X(_14168_));
 sky130_fd_sc_hd__and2_1 _19105_ (.A(_14168_),
    .B(_00294_),
    .X(_00295_));
 sky130_vsdinv _19106_ (.A(\cpuregs[14][29] ),
    .Y(_01144_));
 sky130_vsdinv _19107_ (.A(\cpuregs[15][29] ),
    .Y(_01145_));
 sky130_vsdinv _19108_ (.A(\cpuregs[16][29] ),
    .Y(_01148_));
 sky130_vsdinv _19109_ (.A(\cpuregs[17][29] ),
    .Y(_01149_));
 sky130_vsdinv _19110_ (.A(\cpuregs[18][29] ),
    .Y(_01150_));
 sky130_vsdinv _19111_ (.A(\cpuregs[19][29] ),
    .Y(_01151_));
 sky130_vsdinv _19112_ (.A(\cpuregs[0][30] ),
    .Y(_01154_));
 sky130_vsdinv _19113_ (.A(\cpuregs[1][30] ),
    .Y(_01155_));
 sky130_vsdinv _19114_ (.A(\cpuregs[2][30] ),
    .Y(_01156_));
 sky130_vsdinv _19115_ (.A(\cpuregs[3][30] ),
    .Y(_01157_));
 sky130_vsdinv _19116_ (.A(\cpuregs[4][30] ),
    .Y(_01159_));
 sky130_vsdinv _19117_ (.A(\cpuregs[5][30] ),
    .Y(_01160_));
 sky130_vsdinv _19118_ (.A(\cpuregs[6][30] ),
    .Y(_01161_));
 sky130_vsdinv _19119_ (.A(\cpuregs[7][30] ),
    .Y(_01162_));
 sky130_vsdinv _19120_ (.A(\cpuregs[8][30] ),
    .Y(_01164_));
 sky130_vsdinv _19121_ (.A(\cpuregs[9][30] ),
    .Y(_01165_));
 sky130_vsdinv _19122_ (.A(\cpuregs[10][30] ),
    .Y(_01166_));
 sky130_vsdinv _19123_ (.A(\cpuregs[11][30] ),
    .Y(_01167_));
 sky130_vsdinv _19124_ (.A(\cpuregs[12][30] ),
    .Y(_01169_));
 sky130_vsdinv _19125_ (.A(\cpuregs[13][30] ),
    .Y(_01170_));
 sky130_vsdinv _19126_ (.A(\cpuregs[14][30] ),
    .Y(_01171_));
 sky130_vsdinv _19127_ (.A(\cpuregs[15][30] ),
    .Y(_01172_));
 sky130_vsdinv _19128_ (.A(\cpuregs[16][30] ),
    .Y(_01175_));
 sky130_vsdinv _19129_ (.A(\cpuregs[17][30] ),
    .Y(_01176_));
 sky130_vsdinv _19130_ (.A(\cpuregs[18][30] ),
    .Y(_01177_));
 sky130_vsdinv _19131_ (.A(\cpuregs[19][30] ),
    .Y(_01178_));
 sky130_vsdinv _19132_ (.A(\cpuregs[0][31] ),
    .Y(_01181_));
 sky130_vsdinv _19133_ (.A(\cpuregs[1][31] ),
    .Y(_01182_));
 sky130_vsdinv _19134_ (.A(\cpuregs[2][31] ),
    .Y(_01183_));
 sky130_vsdinv _19135_ (.A(\cpuregs[3][31] ),
    .Y(_01184_));
 sky130_vsdinv _19136_ (.A(\cpuregs[4][31] ),
    .Y(_01186_));
 sky130_vsdinv _19137_ (.A(\cpuregs[5][31] ),
    .Y(_01187_));
 sky130_vsdinv _19138_ (.A(\cpuregs[6][31] ),
    .Y(_01188_));
 sky130_vsdinv _19139_ (.A(\cpuregs[7][31] ),
    .Y(_01189_));
 sky130_vsdinv _19140_ (.A(\cpuregs[8][31] ),
    .Y(_01191_));
 sky130_vsdinv _19141_ (.A(\cpuregs[9][31] ),
    .Y(_01192_));
 sky130_vsdinv _19142_ (.A(\cpuregs[10][31] ),
    .Y(_01193_));
 sky130_vsdinv _19143_ (.A(\cpuregs[11][31] ),
    .Y(_01194_));
 sky130_vsdinv _19144_ (.A(\cpuregs[12][31] ),
    .Y(_01196_));
 sky130_vsdinv _19145_ (.A(\cpuregs[13][31] ),
    .Y(_01197_));
 sky130_vsdinv _19146_ (.A(\cpuregs[14][31] ),
    .Y(_01198_));
 sky130_vsdinv _19147_ (.A(\cpuregs[15][31] ),
    .Y(_01199_));
 sky130_vsdinv _19148_ (.A(\cpuregs[16][31] ),
    .Y(_01202_));
 sky130_vsdinv _19149_ (.A(\cpuregs[17][31] ),
    .Y(_01203_));
 sky130_vsdinv _19150_ (.A(\cpuregs[18][31] ),
    .Y(_01204_));
 sky130_vsdinv _19151_ (.A(\cpuregs[19][31] ),
    .Y(_01205_));
 sky130_vsdinv _19152_ (.A(\timer[26] ),
    .Y(_14169_));
 sky130_vsdinv _19153_ (.A(\timer[18] ),
    .Y(_14170_));
 sky130_fd_sc_hd__or2_1 _19154_ (.A(\timer[1] ),
    .B(\timer[0] ),
    .X(_14171_));
 sky130_fd_sc_hd__or2_1 _19155_ (.A(\timer[2] ),
    .B(_14171_),
    .X(_14172_));
 sky130_fd_sc_hd__or2_1 _19156_ (.A(\timer[3] ),
    .B(_14172_),
    .X(_14173_));
 sky130_fd_sc_hd__or3_1 _19157_ (.A(\timer[5] ),
    .B(\timer[4] ),
    .C(_14173_),
    .X(_14174_));
 sky130_fd_sc_hd__or2_1 _19158_ (.A(\timer[6] ),
    .B(_14174_),
    .X(_14175_));
 sky130_fd_sc_hd__or2_1 _19159_ (.A(\timer[7] ),
    .B(_14175_),
    .X(_14176_));
 sky130_fd_sc_hd__or2_1 _19160_ (.A(\timer[8] ),
    .B(_14176_),
    .X(_14177_));
 sky130_fd_sc_hd__or2_1 _19161_ (.A(\timer[9] ),
    .B(_14177_),
    .X(_14178_));
 sky130_fd_sc_hd__or2_1 _19162_ (.A(\timer[10] ),
    .B(_14178_),
    .X(_14179_));
 sky130_fd_sc_hd__or2_1 _19163_ (.A(\timer[11] ),
    .B(_14179_),
    .X(_14180_));
 sky130_fd_sc_hd__or2_1 _19164_ (.A(\timer[12] ),
    .B(_14180_),
    .X(_14181_));
 sky130_fd_sc_hd__or2_1 _19165_ (.A(\timer[13] ),
    .B(_14181_),
    .X(_14182_));
 sky130_fd_sc_hd__or2_1 _19166_ (.A(\timer[14] ),
    .B(_14182_),
    .X(_14183_));
 sky130_fd_sc_hd__or2_1 _19167_ (.A(\timer[15] ),
    .B(_14183_),
    .X(_14184_));
 sky130_fd_sc_hd__or2_2 _19168_ (.A(\timer[16] ),
    .B(_14184_),
    .X(_14185_));
 sky130_fd_sc_hd__nor2_2 _19169_ (.A(\timer[17] ),
    .B(_14185_),
    .Y(_14186_));
 sky130_fd_sc_hd__nand2_1 _19170_ (.A(_14170_),
    .B(_14186_),
    .Y(_14187_));
 sky130_fd_sc_hd__or2_1 _19171_ (.A(\timer[19] ),
    .B(_14187_),
    .X(_14188_));
 sky130_fd_sc_hd__or2_1 _19172_ (.A(\timer[20] ),
    .B(_14188_),
    .X(_14189_));
 sky130_fd_sc_hd__or2_1 _19173_ (.A(\timer[21] ),
    .B(_14189_),
    .X(_14190_));
 sky130_fd_sc_hd__or2_1 _19174_ (.A(\timer[22] ),
    .B(_14190_),
    .X(_14191_));
 sky130_fd_sc_hd__or2_1 _19175_ (.A(\timer[23] ),
    .B(_14191_),
    .X(_14192_));
 sky130_fd_sc_hd__or2_2 _19176_ (.A(\timer[24] ),
    .B(_14192_),
    .X(_14193_));
 sky130_fd_sc_hd__nor2_2 _19177_ (.A(\timer[25] ),
    .B(_14193_),
    .Y(_14194_));
 sky130_fd_sc_hd__nand2_1 _19178_ (.A(_14169_),
    .B(_14194_),
    .Y(_14195_));
 sky130_fd_sc_hd__or2_1 _19179_ (.A(\timer[27] ),
    .B(_14195_),
    .X(_14196_));
 sky130_fd_sc_hd__or2_1 _19180_ (.A(\timer[28] ),
    .B(_14196_),
    .X(_14197_));
 sky130_fd_sc_hd__or2_1 _19181_ (.A(\timer[29] ),
    .B(_14197_),
    .X(_14198_));
 sky130_fd_sc_hd__or2_4 _19182_ (.A(\timer[30] ),
    .B(_14198_),
    .X(_14199_));
 sky130_fd_sc_hd__nor2_8 _19183_ (.A(\timer[31] ),
    .B(_14199_),
    .Y(_01208_));
 sky130_fd_sc_hd__nor2_1 _19184_ (.A(\timer[0] ),
    .B(_01208_),
    .Y(_01209_));
 sky130_vsdinv _19185_ (.A(\timer[1] ),
    .Y(_14200_));
 sky130_vsdinv _19186_ (.A(\timer[0] ),
    .Y(_14201_));
 sky130_fd_sc_hd__o21ai_1 _19187_ (.A1(_14200_),
    .A2(_14201_),
    .B1(_14171_),
    .Y(_01211_));
 sky130_fd_sc_hd__a21bo_1 _19188_ (.A1(\timer[2] ),
    .A2(_14171_),
    .B1_N(_14172_),
    .X(_01214_));
 sky130_fd_sc_hd__a21bo_1 _19189_ (.A1(\timer[3] ),
    .A2(_14172_),
    .B1_N(_14173_),
    .X(_01217_));
 sky130_fd_sc_hd__clkbuf_2 _19190_ (.A(\timer[4] ),
    .X(_14202_));
 sky130_fd_sc_hd__nor2_1 _19191_ (.A(_14202_),
    .B(_14173_),
    .Y(_14203_));
 sky130_fd_sc_hd__a21o_1 _19192_ (.A1(_14202_),
    .A2(_14173_),
    .B1(_14203_),
    .X(_01220_));
 sky130_vsdinv _19193_ (.A(\timer[5] ),
    .Y(_14204_));
 sky130_fd_sc_hd__o21ai_1 _19194_ (.A1(_14204_),
    .A2(_14203_),
    .B1(_14174_),
    .Y(_01223_));
 sky130_vsdinv _19195_ (.A(_14175_),
    .Y(_14205_));
 sky130_fd_sc_hd__a21o_1 _19196_ (.A1(\timer[6] ),
    .A2(_14174_),
    .B1(_14205_),
    .X(_01226_));
 sky130_vsdinv _19197_ (.A(\timer[7] ),
    .Y(_14206_));
 sky130_fd_sc_hd__o21ai_1 _19198_ (.A1(_14206_),
    .A2(_14205_),
    .B1(_14176_),
    .Y(_01229_));
 sky130_vsdinv _19199_ (.A(_14177_),
    .Y(_14207_));
 sky130_fd_sc_hd__a21o_1 _19200_ (.A1(\timer[8] ),
    .A2(_14176_),
    .B1(_14207_),
    .X(_01232_));
 sky130_vsdinv _19201_ (.A(\timer[9] ),
    .Y(_14208_));
 sky130_fd_sc_hd__o21ai_1 _19202_ (.A1(_14208_),
    .A2(_14207_),
    .B1(_14178_),
    .Y(_01235_));
 sky130_vsdinv _19203_ (.A(_14179_),
    .Y(_14209_));
 sky130_fd_sc_hd__a21o_1 _19204_ (.A1(\timer[10] ),
    .A2(_14178_),
    .B1(_14209_),
    .X(_01238_));
 sky130_vsdinv _19205_ (.A(\timer[11] ),
    .Y(_14210_));
 sky130_fd_sc_hd__o21ai_1 _19206_ (.A1(_14210_),
    .A2(_14209_),
    .B1(_14180_),
    .Y(_01241_));
 sky130_vsdinv _19207_ (.A(_14181_),
    .Y(_14211_));
 sky130_fd_sc_hd__a21o_1 _19208_ (.A1(\timer[12] ),
    .A2(_14180_),
    .B1(_14211_),
    .X(_01244_));
 sky130_vsdinv _19209_ (.A(\timer[13] ),
    .Y(_14212_));
 sky130_fd_sc_hd__o21ai_1 _19210_ (.A1(_14212_),
    .A2(_14211_),
    .B1(_14182_),
    .Y(_01247_));
 sky130_vsdinv _19211_ (.A(_14183_),
    .Y(_14213_));
 sky130_fd_sc_hd__a21o_1 _19212_ (.A1(\timer[14] ),
    .A2(_14182_),
    .B1(_14213_),
    .X(_01250_));
 sky130_vsdinv _19213_ (.A(\timer[15] ),
    .Y(_14214_));
 sky130_fd_sc_hd__o21ai_1 _19214_ (.A1(_14214_),
    .A2(_14213_),
    .B1(_14184_),
    .Y(_01253_));
 sky130_fd_sc_hd__a21bo_1 _19215_ (.A1(\timer[16] ),
    .A2(_14184_),
    .B1_N(_14185_),
    .X(_01256_));
 sky130_fd_sc_hd__a21o_1 _19216_ (.A1(\timer[17] ),
    .A2(_14185_),
    .B1(_14186_),
    .X(_01259_));
 sky130_fd_sc_hd__o21ai_1 _19217_ (.A1(_14170_),
    .A2(_14186_),
    .B1(_14187_),
    .Y(_01262_));
 sky130_vsdinv _19218_ (.A(_14188_),
    .Y(_14215_));
 sky130_fd_sc_hd__a21o_1 _19219_ (.A1(\timer[19] ),
    .A2(_14187_),
    .B1(_14215_),
    .X(_01265_));
 sky130_vsdinv _19220_ (.A(\timer[20] ),
    .Y(_14216_));
 sky130_fd_sc_hd__o21ai_1 _19221_ (.A1(_14216_),
    .A2(_14215_),
    .B1(_14189_),
    .Y(_01268_));
 sky130_vsdinv _19222_ (.A(_14190_),
    .Y(_14217_));
 sky130_fd_sc_hd__a21o_1 _19223_ (.A1(\timer[21] ),
    .A2(_14189_),
    .B1(_14217_),
    .X(_01271_));
 sky130_vsdinv _19224_ (.A(\timer[22] ),
    .Y(_14218_));
 sky130_fd_sc_hd__o21ai_1 _19225_ (.A1(_14218_),
    .A2(_14217_),
    .B1(_14191_),
    .Y(_01274_));
 sky130_vsdinv _19226_ (.A(_14192_),
    .Y(_14219_));
 sky130_fd_sc_hd__a21o_1 _19227_ (.A1(\timer[23] ),
    .A2(_14191_),
    .B1(_14219_),
    .X(_01277_));
 sky130_vsdinv _19228_ (.A(\timer[24] ),
    .Y(_14220_));
 sky130_fd_sc_hd__o21ai_1 _19229_ (.A1(_14220_),
    .A2(_14219_),
    .B1(_14193_),
    .Y(_01280_));
 sky130_fd_sc_hd__a21o_1 _19230_ (.A1(\timer[25] ),
    .A2(_14193_),
    .B1(_14194_),
    .X(_01283_));
 sky130_fd_sc_hd__o21ai_1 _19231_ (.A1(_14169_),
    .A2(_14194_),
    .B1(_14195_),
    .Y(_01286_));
 sky130_vsdinv _19232_ (.A(_14196_),
    .Y(_14221_));
 sky130_fd_sc_hd__a21o_1 _19233_ (.A1(\timer[27] ),
    .A2(_14195_),
    .B1(_14221_),
    .X(_01289_));
 sky130_vsdinv _19234_ (.A(\timer[28] ),
    .Y(_14222_));
 sky130_fd_sc_hd__o21ai_1 _19235_ (.A1(_14222_),
    .A2(_14221_),
    .B1(_14197_),
    .Y(_01292_));
 sky130_vsdinv _19236_ (.A(_14198_),
    .Y(_14223_));
 sky130_fd_sc_hd__a21o_1 _19237_ (.A1(\timer[29] ),
    .A2(_14197_),
    .B1(_14223_),
    .X(_01295_));
 sky130_vsdinv _19238_ (.A(\timer[30] ),
    .Y(_14224_));
 sky130_fd_sc_hd__o21ai_1 _19239_ (.A1(_14224_),
    .A2(_14223_),
    .B1(_14199_),
    .Y(_01298_));
 sky130_fd_sc_hd__a21o_1 _19240_ (.A1(\timer[31] ),
    .A2(_14199_),
    .B1(_01208_),
    .X(_01301_));
 sky130_fd_sc_hd__nor2_1 _19241_ (.A(_13252_),
    .B(_13818_),
    .Y(_01315_));
 sky130_fd_sc_hd__nor2_1 _19242_ (.A(_13252_),
    .B(_13825_),
    .Y(_01317_));
 sky130_fd_sc_hd__nor2_1 _19243_ (.A(_13252_),
    .B(_13828_),
    .Y(_01319_));
 sky130_fd_sc_hd__buf_2 _19244_ (.A(_13251_),
    .X(_14225_));
 sky130_fd_sc_hd__buf_1 _19245_ (.A(_14225_),
    .X(_14226_));
 sky130_fd_sc_hd__nor2_1 _19246_ (.A(_14226_),
    .B(_13833_),
    .Y(_01321_));
 sky130_fd_sc_hd__nor2_1 _19247_ (.A(_14226_),
    .B(_13839_),
    .Y(_01323_));
 sky130_fd_sc_hd__nor2_1 _19248_ (.A(_14226_),
    .B(_13844_),
    .Y(_01325_));
 sky130_fd_sc_hd__nor2_1 _19249_ (.A(_14226_),
    .B(_13849_),
    .Y(_01327_));
 sky130_fd_sc_hd__buf_1 _19250_ (.A(_14225_),
    .X(_14227_));
 sky130_fd_sc_hd__nor2_1 _19251_ (.A(_14227_),
    .B(_13855_),
    .Y(_01329_));
 sky130_fd_sc_hd__nor2_1 _19252_ (.A(_14227_),
    .B(_13864_),
    .Y(_01331_));
 sky130_fd_sc_hd__nor2_1 _19253_ (.A(_14227_),
    .B(_13869_),
    .Y(_01333_));
 sky130_fd_sc_hd__nor2_1 _19254_ (.A(_14227_),
    .B(_13874_),
    .Y(_01335_));
 sky130_fd_sc_hd__clkbuf_2 _19255_ (.A(_14225_),
    .X(_14228_));
 sky130_fd_sc_hd__nor2_1 _19256_ (.A(_14228_),
    .B(_13881_),
    .Y(_01337_));
 sky130_fd_sc_hd__nor2_1 _19257_ (.A(_14228_),
    .B(_13887_),
    .Y(_01339_));
 sky130_fd_sc_hd__nor2_1 _19258_ (.A(_14228_),
    .B(_13893_),
    .Y(_01341_));
 sky130_fd_sc_hd__nor2_1 _19259_ (.A(_14228_),
    .B(_13898_),
    .Y(_01343_));
 sky130_fd_sc_hd__buf_1 _19260_ (.A(_14225_),
    .X(_14229_));
 sky130_vsdinv _19261_ (.A(\decoded_imm[20] ),
    .Y(_14230_));
 sky130_fd_sc_hd__clkbuf_2 _19262_ (.A(_14230_),
    .X(_14231_));
 sky130_fd_sc_hd__nor2_1 _19263_ (.A(_14229_),
    .B(_14231_),
    .Y(_01345_));
 sky130_vsdinv _19264_ (.A(\decoded_imm[21] ),
    .Y(_14232_));
 sky130_fd_sc_hd__clkbuf_2 _19265_ (.A(_14232_),
    .X(_14233_));
 sky130_fd_sc_hd__nor2_1 _19266_ (.A(_14229_),
    .B(_14233_),
    .Y(_01347_));
 sky130_vsdinv _19267_ (.A(\decoded_imm[22] ),
    .Y(_14234_));
 sky130_fd_sc_hd__clkbuf_2 _19268_ (.A(_14234_),
    .X(_14235_));
 sky130_fd_sc_hd__nor2_1 _19269_ (.A(_14229_),
    .B(_14235_),
    .Y(_01349_));
 sky130_vsdinv _19270_ (.A(\decoded_imm[23] ),
    .Y(_14236_));
 sky130_fd_sc_hd__buf_2 _19271_ (.A(_14236_),
    .X(_14237_));
 sky130_fd_sc_hd__nor2_1 _19272_ (.A(_14229_),
    .B(_14237_),
    .Y(_01351_));
 sky130_fd_sc_hd__clkbuf_2 _19273_ (.A(_13251_),
    .X(_14238_));
 sky130_vsdinv _19274_ (.A(\decoded_imm[24] ),
    .Y(_14239_));
 sky130_fd_sc_hd__clkbuf_2 _19275_ (.A(_14239_),
    .X(_14240_));
 sky130_fd_sc_hd__nor2_1 _19276_ (.A(_14238_),
    .B(_14240_),
    .Y(_01353_));
 sky130_vsdinv _19277_ (.A(\decoded_imm[25] ),
    .Y(_14241_));
 sky130_fd_sc_hd__nor2_1 _19278_ (.A(_14238_),
    .B(_14241_),
    .Y(_01355_));
 sky130_vsdinv _19279_ (.A(\decoded_imm[26] ),
    .Y(_14242_));
 sky130_fd_sc_hd__clkbuf_2 _19280_ (.A(_14242_),
    .X(_14243_));
 sky130_fd_sc_hd__nor2_1 _19281_ (.A(_14238_),
    .B(_14243_),
    .Y(_01357_));
 sky130_vsdinv _19282_ (.A(\decoded_imm[27] ),
    .Y(_14244_));
 sky130_fd_sc_hd__nor2_1 _19283_ (.A(_14238_),
    .B(_14244_),
    .Y(_01359_));
 sky130_fd_sc_hd__clkbuf_2 _19284_ (.A(_13251_),
    .X(_14245_));
 sky130_vsdinv _19285_ (.A(\decoded_imm[28] ),
    .Y(_14246_));
 sky130_fd_sc_hd__nor2_1 _19286_ (.A(_14245_),
    .B(_14246_),
    .Y(_01361_));
 sky130_vsdinv _19287_ (.A(\decoded_imm[29] ),
    .Y(_14247_));
 sky130_fd_sc_hd__nor2_1 _19288_ (.A(_14245_),
    .B(_14247_),
    .Y(_01363_));
 sky130_vsdinv _19289_ (.A(\decoded_imm[30] ),
    .Y(_14248_));
 sky130_fd_sc_hd__buf_2 _19290_ (.A(_14248_),
    .X(_14249_));
 sky130_fd_sc_hd__nor2_1 _19291_ (.A(_14245_),
    .B(_14249_),
    .Y(_01365_));
 sky130_fd_sc_hd__nor2_1 _19292_ (.A(_14245_),
    .B(_13940_),
    .Y(_01367_));
 sky130_fd_sc_hd__clkbuf_2 _19293_ (.A(instr_lui),
    .X(_14250_));
 sky130_vsdinv _19294_ (.A(\reg_next_pc[0] ),
    .Y(_14251_));
 sky130_fd_sc_hd__nor2_1 _19295_ (.A(_14250_),
    .B(_14251_),
    .Y(_01369_));
 sky130_fd_sc_hd__clkbuf_2 _19296_ (.A(_13969_),
    .X(_14252_));
 sky130_fd_sc_hd__nor2_2 _19297_ (.A(_13277_),
    .B(_13969_),
    .Y(_14253_));
 sky130_fd_sc_hd__a21oi_1 _19298_ (.A1(_13278_),
    .A2(_14252_),
    .B1(_14253_),
    .Y(_01371_));
 sky130_vsdinv _19299_ (.A(\reg_pc[1] ),
    .Y(_14254_));
 sky130_fd_sc_hd__buf_1 _19300_ (.A(_13373_),
    .X(_14255_));
 sky130_fd_sc_hd__nor2_1 _19301_ (.A(_14254_),
    .B(_14255_),
    .Y(_01372_));
 sky130_vsdinv _19302_ (.A(net317),
    .Y(_14256_));
 sky130_fd_sc_hd__o22a_1 _19303_ (.A1(_14256_),
    .A2(_13790_),
    .B1(net317),
    .B2(\decoded_imm[1] ),
    .X(_14257_));
 sky130_fd_sc_hd__o2bb2a_1 _19304_ (.A1_N(_14253_),
    .A2_N(_14257_),
    .B1(_14253_),
    .B2(_14257_),
    .X(_01374_));
 sky130_vsdinv _19305_ (.A(\reg_pc[2] ),
    .Y(_14258_));
 sky130_fd_sc_hd__clkbuf_2 _19306_ (.A(_14258_),
    .X(_02073_));
 sky130_fd_sc_hd__nor2_1 _19307_ (.A(_02073_),
    .B(_14255_),
    .Y(_01375_));
 sky130_fd_sc_hd__a22o_1 _19308_ (.A1(_13484_),
    .A2(\decoded_imm[1] ),
    .B1(_14253_),
    .B2(_14257_),
    .X(_14259_));
 sky130_fd_sc_hd__clkbuf_2 _19309_ (.A(\decoded_imm[2] ),
    .X(_14260_));
 sky130_fd_sc_hd__nor2_1 _19310_ (.A(net328),
    .B(_14260_),
    .Y(_14261_));
 sky130_fd_sc_hd__a21oi_1 _19311_ (.A1(_13483_),
    .A2(_14260_),
    .B1(_14261_),
    .Y(_14262_));
 sky130_vsdinv _19312_ (.A(_14259_),
    .Y(_14263_));
 sky130_vsdinv _19313_ (.A(_14262_),
    .Y(_14264_));
 sky130_fd_sc_hd__o22a_1 _19314_ (.A1(_14259_),
    .A2(_14262_),
    .B1(_14263_),
    .B2(_14264_),
    .X(_01377_));
 sky130_vsdinv _19315_ (.A(\reg_pc[3] ),
    .Y(_14265_));
 sky130_fd_sc_hd__nor2_1 _19316_ (.A(_14265_),
    .B(_14255_),
    .Y(_01378_));
 sky130_vsdinv _19317_ (.A(_13481_),
    .Y(_14266_));
 sky130_fd_sc_hd__o22a_1 _19318_ (.A1(_14266_),
    .A2(_13797_),
    .B1(_14263_),
    .B2(_14261_),
    .X(_14267_));
 sky130_fd_sc_hd__clkbuf_2 _19319_ (.A(\decoded_imm[3] ),
    .X(_14268_));
 sky130_fd_sc_hd__nor2_1 _19320_ (.A(_13477_),
    .B(_14268_),
    .Y(_14269_));
 sky130_fd_sc_hd__a21o_1 _19321_ (.A1(_13479_),
    .A2(_14268_),
    .B1(_14269_),
    .X(_14270_));
 sky130_fd_sc_hd__o2bb2a_1 _19322_ (.A1_N(_14267_),
    .A2_N(_14270_),
    .B1(_14267_),
    .B2(_14270_),
    .X(_01380_));
 sky130_vsdinv _19323_ (.A(_12081_),
    .Y(_14271_));
 sky130_fd_sc_hd__nor2_1 _19324_ (.A(_14271_),
    .B(_14255_),
    .Y(_01381_));
 sky130_vsdinv _19325_ (.A(net331),
    .Y(_14272_));
 sky130_fd_sc_hd__o22a_1 _19326_ (.A1(_14272_),
    .A2(_13805_),
    .B1(_14267_),
    .B2(_14269_),
    .X(_14273_));
 sky130_fd_sc_hd__nor2_1 _19327_ (.A(_13473_),
    .B(\decoded_imm[4] ),
    .Y(_14274_));
 sky130_fd_sc_hd__a21o_1 _19328_ (.A1(_13475_),
    .A2(\decoded_imm[4] ),
    .B1(_14274_),
    .X(_14275_));
 sky130_fd_sc_hd__o2bb2a_1 _19329_ (.A1_N(_14273_),
    .A2_N(_14275_),
    .B1(_14273_),
    .B2(_14275_),
    .X(_01383_));
 sky130_vsdinv _19330_ (.A(\reg_pc[5] ),
    .Y(_14276_));
 sky130_fd_sc_hd__buf_1 _19331_ (.A(_13373_),
    .X(_14277_));
 sky130_fd_sc_hd__nor2_1 _19332_ (.A(_14276_),
    .B(_14277_),
    .Y(_01384_));
 sky130_vsdinv _19333_ (.A(net332),
    .Y(_14278_));
 sky130_fd_sc_hd__o22a_2 _19334_ (.A1(_14278_),
    .A2(_13812_),
    .B1(_14273_),
    .B2(_14274_),
    .X(_14279_));
 sky130_fd_sc_hd__clkbuf_2 _19335_ (.A(\decoded_imm[5] ),
    .X(_14280_));
 sky130_fd_sc_hd__nor2_2 _19336_ (.A(_13470_),
    .B(_14280_),
    .Y(_04073_));
 sky130_fd_sc_hd__a21o_1 _19337_ (.A1(_13472_),
    .A2(_14280_),
    .B1(_04073_),
    .X(_04074_));
 sky130_fd_sc_hd__o2bb2a_1 _19338_ (.A1_N(_14279_),
    .A2_N(_04074_),
    .B1(_14279_),
    .B2(_04074_),
    .X(_01386_));
 sky130_vsdinv _19339_ (.A(_12076_),
    .Y(_04075_));
 sky130_fd_sc_hd__nor2_1 _19340_ (.A(_04075_),
    .B(_14277_),
    .Y(_01387_));
 sky130_vsdinv _19341_ (.A(net333),
    .Y(_04076_));
 sky130_fd_sc_hd__o22ai_4 _19342_ (.A1(_04076_),
    .A2(_13818_),
    .B1(_14279_),
    .B2(_04073_),
    .Y(_04077_));
 sky130_vsdinv _19343_ (.A(net334),
    .Y(_04078_));
 sky130_fd_sc_hd__o22a_1 _19344_ (.A1(_04078_),
    .A2(_13825_),
    .B1(net334),
    .B2(\decoded_imm[6] ),
    .X(_04079_));
 sky130_fd_sc_hd__o2bb2a_1 _19345_ (.A1_N(_04077_),
    .A2_N(_04079_),
    .B1(_04077_),
    .B2(_04079_),
    .X(_01389_));
 sky130_vsdinv _19346_ (.A(\reg_pc[7] ),
    .Y(_04080_));
 sky130_fd_sc_hd__nor2_1 _19347_ (.A(_04080_),
    .B(_14277_),
    .Y(_01390_));
 sky130_fd_sc_hd__clkbuf_2 _19348_ (.A(\decoded_imm[7] ),
    .X(_04081_));
 sky130_fd_sc_hd__nor2_1 _19349_ (.A(net335),
    .B(_04081_),
    .Y(_04082_));
 sky130_fd_sc_hd__a21oi_2 _19350_ (.A1(_13463_),
    .A2(_04081_),
    .B1(_04082_),
    .Y(_04083_));
 sky130_fd_sc_hd__a22o_1 _19351_ (.A1(_13469_),
    .A2(\decoded_imm[6] ),
    .B1(_04077_),
    .B2(_04079_),
    .X(_04084_));
 sky130_fd_sc_hd__a2bb2oi_1 _19352_ (.A1_N(_04083_),
    .A2_N(_04084_),
    .B1(_04083_),
    .B2(_04084_),
    .Y(_01392_));
 sky130_vsdinv _19353_ (.A(\reg_pc[8] ),
    .Y(_04085_));
 sky130_fd_sc_hd__buf_1 _19354_ (.A(_04085_),
    .X(_04086_));
 sky130_fd_sc_hd__nor2_1 _19355_ (.A(_04086_),
    .B(_14277_),
    .Y(_01393_));
 sky130_vsdinv _19356_ (.A(net335),
    .Y(_04087_));
 sky130_fd_sc_hd__o32a_1 _19357_ (.A1(_04078_),
    .A2(_13824_),
    .A3(_04082_),
    .B1(_04087_),
    .B2(_13828_),
    .X(_04088_));
 sky130_vsdinv _19358_ (.A(_04088_),
    .Y(_04089_));
 sky130_fd_sc_hd__a31o_1 _19359_ (.A1(_04079_),
    .A2(_04083_),
    .A3(_04077_),
    .B1(_04089_),
    .X(_04090_));
 sky130_vsdinv _19360_ (.A(_04090_),
    .Y(_04091_));
 sky130_vsdinv _19361_ (.A(net336),
    .Y(_04092_));
 sky130_fd_sc_hd__o22a_1 _19362_ (.A1(_04092_),
    .A2(_13832_),
    .B1(_13459_),
    .B2(\decoded_imm[8] ),
    .X(_04093_));
 sky130_vsdinv _19363_ (.A(_04093_),
    .Y(_04094_));
 sky130_fd_sc_hd__o22a_1 _19364_ (.A1(_04091_),
    .A2(_04094_),
    .B1(_04090_),
    .B2(_04093_),
    .X(_01395_));
 sky130_vsdinv _19365_ (.A(\reg_pc[9] ),
    .Y(_04095_));
 sky130_fd_sc_hd__clkbuf_2 _19366_ (.A(_13373_),
    .X(_04096_));
 sky130_fd_sc_hd__nor2_1 _19367_ (.A(_04095_),
    .B(_04096_),
    .Y(_01396_));
 sky130_fd_sc_hd__buf_1 _19368_ (.A(net337),
    .X(_04097_));
 sky130_fd_sc_hd__clkbuf_2 _19369_ (.A(\decoded_imm[9] ),
    .X(_04098_));
 sky130_fd_sc_hd__nor2_1 _19370_ (.A(_04097_),
    .B(_04098_),
    .Y(_04099_));
 sky130_fd_sc_hd__a21o_1 _19371_ (.A1(_04097_),
    .A2(_04098_),
    .B1(_04099_),
    .X(_04100_));
 sky130_fd_sc_hd__o22a_1 _19372_ (.A1(_04092_),
    .A2(_13833_),
    .B1(_04091_),
    .B2(_04094_),
    .X(_04101_));
 sky130_fd_sc_hd__o2bb2a_1 _19373_ (.A1_N(_04100_),
    .A2_N(_04101_),
    .B1(_04100_),
    .B2(_04101_),
    .X(_01398_));
 sky130_vsdinv _19374_ (.A(\reg_pc[10] ),
    .Y(_04102_));
 sky130_fd_sc_hd__nor2_1 _19375_ (.A(_04102_),
    .B(_04096_),
    .Y(_01399_));
 sky130_vsdinv _19376_ (.A(net307),
    .Y(_04103_));
 sky130_fd_sc_hd__a22o_1 _19377_ (.A1(_13455_),
    .A2(\decoded_imm[10] ),
    .B1(_04103_),
    .B2(_13844_),
    .X(_04104_));
 sky130_vsdinv _19378_ (.A(_04097_),
    .Y(_04105_));
 sky130_fd_sc_hd__o32a_1 _19379_ (.A1(_04092_),
    .A2(_13832_),
    .A3(_04099_),
    .B1(_04105_),
    .B2(_13839_),
    .X(_04106_));
 sky130_fd_sc_hd__o31a_1 _19380_ (.A1(_04094_),
    .A2(_04100_),
    .A3(_04091_),
    .B1(_04106_),
    .X(_04107_));
 sky130_fd_sc_hd__a2bb2oi_1 _19381_ (.A1_N(_04104_),
    .A2_N(_04107_),
    .B1(_04104_),
    .B2(_04107_),
    .Y(_01401_));
 sky130_vsdinv _19382_ (.A(\reg_pc[11] ),
    .Y(_04108_));
 sky130_fd_sc_hd__buf_1 _19383_ (.A(_04108_),
    .X(_04109_));
 sky130_fd_sc_hd__nor2_1 _19384_ (.A(_04109_),
    .B(_04096_),
    .Y(_01402_));
 sky130_vsdinv _19385_ (.A(net308),
    .Y(_04110_));
 sky130_fd_sc_hd__a22o_1 _19386_ (.A1(_13452_),
    .A2(\decoded_imm[11] ),
    .B1(_04110_),
    .B2(_13849_),
    .X(_04111_));
 sky130_fd_sc_hd__buf_1 _19387_ (.A(_04103_),
    .X(_04112_));
 sky130_fd_sc_hd__o22a_1 _19388_ (.A1(_04112_),
    .A2(_13844_),
    .B1(_04104_),
    .B2(_04107_),
    .X(_04113_));
 sky130_fd_sc_hd__a2bb2oi_1 _19389_ (.A1_N(_04111_),
    .A2_N(_04113_),
    .B1(_04111_),
    .B2(_04113_),
    .Y(_01404_));
 sky130_vsdinv _19390_ (.A(\reg_pc[12] ),
    .Y(_04114_));
 sky130_fd_sc_hd__nor2_1 _19391_ (.A(_04114_),
    .B(_04096_),
    .Y(_01405_));
 sky130_vsdinv _19392_ (.A(net309),
    .Y(_04115_));
 sky130_fd_sc_hd__a22o_1 _19393_ (.A1(_13449_),
    .A2(\decoded_imm[12] ),
    .B1(_04115_),
    .B2(_13855_),
    .X(_04116_));
 sky130_fd_sc_hd__buf_1 _19394_ (.A(_04110_),
    .X(_04117_));
 sky130_fd_sc_hd__o22a_1 _19395_ (.A1(_04117_),
    .A2(_13849_),
    .B1(_04111_),
    .B2(_04113_),
    .X(_04118_));
 sky130_fd_sc_hd__a2bb2oi_1 _19396_ (.A1_N(_04116_),
    .A2_N(_04118_),
    .B1(_04116_),
    .B2(_04118_),
    .Y(_01407_));
 sky130_vsdinv _19397_ (.A(\reg_pc[13] ),
    .Y(_04119_));
 sky130_fd_sc_hd__buf_1 _19398_ (.A(_04119_),
    .X(_04120_));
 sky130_fd_sc_hd__clkbuf_4 _19399_ (.A(instr_lui),
    .X(_04121_));
 sky130_fd_sc_hd__buf_1 _19400_ (.A(_04121_),
    .X(_04122_));
 sky130_fd_sc_hd__nor2_1 _19401_ (.A(_04120_),
    .B(_04122_),
    .Y(_01408_));
 sky130_vsdinv _19402_ (.A(net310),
    .Y(_04123_));
 sky130_fd_sc_hd__a22o_1 _19403_ (.A1(_13447_),
    .A2(\decoded_imm[13] ),
    .B1(_04123_),
    .B2(_13864_),
    .X(_04124_));
 sky130_fd_sc_hd__buf_1 _19404_ (.A(_04115_),
    .X(_04125_));
 sky130_fd_sc_hd__o22a_1 _19405_ (.A1(_04125_),
    .A2(_13855_),
    .B1(_04116_),
    .B2(_04118_),
    .X(_04126_));
 sky130_fd_sc_hd__a2bb2oi_1 _19406_ (.A1_N(_04124_),
    .A2_N(_04126_),
    .B1(_04124_),
    .B2(_04126_),
    .Y(_01410_));
 sky130_vsdinv _19407_ (.A(\reg_pc[14] ),
    .Y(_04127_));
 sky130_fd_sc_hd__nor2_1 _19408_ (.A(_04127_),
    .B(_04122_),
    .Y(_01411_));
 sky130_vsdinv _19409_ (.A(net311),
    .Y(_04128_));
 sky130_fd_sc_hd__a22o_1 _19410_ (.A1(_13445_),
    .A2(\decoded_imm[14] ),
    .B1(_04128_),
    .B2(_13869_),
    .X(_04129_));
 sky130_fd_sc_hd__buf_1 _19411_ (.A(_04123_),
    .X(_04130_));
 sky130_fd_sc_hd__o22a_1 _19412_ (.A1(_04130_),
    .A2(_13864_),
    .B1(_04124_),
    .B2(_04126_),
    .X(_04131_));
 sky130_fd_sc_hd__a2bb2oi_1 _19413_ (.A1_N(_04129_),
    .A2_N(_04131_),
    .B1(_04129_),
    .B2(_04131_),
    .Y(_01413_));
 sky130_vsdinv _19414_ (.A(\reg_pc[15] ),
    .Y(_04132_));
 sky130_fd_sc_hd__buf_1 _19415_ (.A(_04132_),
    .X(_04133_));
 sky130_fd_sc_hd__nor2_1 _19416_ (.A(_04133_),
    .B(_04122_),
    .Y(_01414_));
 sky130_vsdinv _19417_ (.A(net312),
    .Y(_04134_));
 sky130_fd_sc_hd__a22o_1 _19418_ (.A1(_13441_),
    .A2(\decoded_imm[15] ),
    .B1(_04134_),
    .B2(_13874_),
    .X(_04135_));
 sky130_fd_sc_hd__buf_1 _19419_ (.A(_04128_),
    .X(_04136_));
 sky130_fd_sc_hd__o22a_1 _19420_ (.A1(_04136_),
    .A2(_13869_),
    .B1(_04129_),
    .B2(_04131_),
    .X(_04137_));
 sky130_fd_sc_hd__a2bb2oi_1 _19421_ (.A1_N(_04135_),
    .A2_N(_04137_),
    .B1(_04135_),
    .B2(_04137_),
    .Y(_01416_));
 sky130_vsdinv _19422_ (.A(\reg_pc[16] ),
    .Y(_04138_));
 sky130_fd_sc_hd__clkbuf_2 _19423_ (.A(_04138_),
    .X(_04139_));
 sky130_fd_sc_hd__nor2_1 _19424_ (.A(_04139_),
    .B(_04122_),
    .Y(_01417_));
 sky130_fd_sc_hd__clkbuf_2 _19425_ (.A(_04134_),
    .X(_04140_));
 sky130_fd_sc_hd__o22a_1 _19426_ (.A1(_04140_),
    .A2(_13874_),
    .B1(_04135_),
    .B2(_04137_),
    .X(_04141_));
 sky130_vsdinv _19427_ (.A(net313),
    .Y(_04142_));
 sky130_fd_sc_hd__o22a_1 _19428_ (.A1(_04142_),
    .A2(_13880_),
    .B1(_13436_),
    .B2(\decoded_imm[16] ),
    .X(_04143_));
 sky130_vsdinv _19429_ (.A(_04143_),
    .Y(_04144_));
 sky130_vsdinv _19430_ (.A(_04141_),
    .Y(_04145_));
 sky130_fd_sc_hd__o22a_1 _19431_ (.A1(_04141_),
    .A2(_04144_),
    .B1(_04145_),
    .B2(_04143_),
    .X(_01419_));
 sky130_vsdinv _19432_ (.A(\reg_pc[17] ),
    .Y(_04146_));
 sky130_fd_sc_hd__buf_1 _19433_ (.A(_04121_),
    .X(_04147_));
 sky130_fd_sc_hd__nor2_1 _19434_ (.A(_04146_),
    .B(_04147_),
    .Y(_01420_));
 sky130_fd_sc_hd__buf_2 _19435_ (.A(\decoded_imm[17] ),
    .X(_04148_));
 sky130_fd_sc_hd__buf_1 _19436_ (.A(net314),
    .X(_04149_));
 sky130_fd_sc_hd__nor2_1 _19437_ (.A(_04149_),
    .B(_04148_),
    .Y(_04150_));
 sky130_fd_sc_hd__a21o_1 _19438_ (.A1(_13434_),
    .A2(_04148_),
    .B1(_04150_),
    .X(_04151_));
 sky130_fd_sc_hd__o22a_1 _19439_ (.A1(_04142_),
    .A2(_13881_),
    .B1(_04141_),
    .B2(_04144_),
    .X(_04152_));
 sky130_fd_sc_hd__o2bb2a_1 _19440_ (.A1_N(_04151_),
    .A2_N(_04152_),
    .B1(_04151_),
    .B2(_04152_),
    .X(_01422_));
 sky130_vsdinv _19441_ (.A(\reg_pc[18] ),
    .Y(_04153_));
 sky130_fd_sc_hd__nor2_1 _19442_ (.A(_04153_),
    .B(_04147_),
    .Y(_01423_));
 sky130_vsdinv _19443_ (.A(net315),
    .Y(_04154_));
 sky130_fd_sc_hd__buf_1 _19444_ (.A(_04154_),
    .X(_04155_));
 sky130_fd_sc_hd__a22o_1 _19445_ (.A1(_13432_),
    .A2(\decoded_imm[18] ),
    .B1(_04155_),
    .B2(_13893_),
    .X(_04156_));
 sky130_vsdinv _19446_ (.A(_04149_),
    .Y(_04157_));
 sky130_fd_sc_hd__o32a_1 _19447_ (.A1(_04142_),
    .A2(_13880_),
    .A3(_04150_),
    .B1(_04157_),
    .B2(_13887_),
    .X(_04158_));
 sky130_fd_sc_hd__o31a_1 _19448_ (.A1(_04144_),
    .A2(_04151_),
    .A3(_04141_),
    .B1(_04158_),
    .X(_04159_));
 sky130_fd_sc_hd__a2bb2oi_1 _19449_ (.A1_N(_04156_),
    .A2_N(_04159_),
    .B1(_04156_),
    .B2(_04159_),
    .Y(_01425_));
 sky130_vsdinv _19450_ (.A(\reg_pc[19] ),
    .Y(_04160_));
 sky130_fd_sc_hd__buf_1 _19451_ (.A(_04160_),
    .X(_04161_));
 sky130_fd_sc_hd__nor2_1 _19452_ (.A(_04161_),
    .B(_04147_),
    .Y(_01426_));
 sky130_vsdinv _19453_ (.A(net316),
    .Y(_04162_));
 sky130_fd_sc_hd__buf_1 _19454_ (.A(_04162_),
    .X(_04163_));
 sky130_fd_sc_hd__a22o_1 _19455_ (.A1(_13429_),
    .A2(\decoded_imm[19] ),
    .B1(_04163_),
    .B2(_13898_),
    .X(_04164_));
 sky130_fd_sc_hd__o22a_1 _19456_ (.A1(_04155_),
    .A2(_13893_),
    .B1(_04156_),
    .B2(_04159_),
    .X(_04165_));
 sky130_fd_sc_hd__a2bb2oi_1 _19457_ (.A1_N(_04164_),
    .A2_N(_04165_),
    .B1(_04164_),
    .B2(_04165_),
    .Y(_01428_));
 sky130_vsdinv _19458_ (.A(\reg_pc[20] ),
    .Y(_04166_));
 sky130_fd_sc_hd__nor2_1 _19459_ (.A(_04166_),
    .B(_04147_),
    .Y(_01429_));
 sky130_vsdinv _19460_ (.A(net318),
    .Y(_04167_));
 sky130_fd_sc_hd__buf_1 _19461_ (.A(_04167_),
    .X(_04168_));
 sky130_fd_sc_hd__a22o_1 _19462_ (.A1(_13426_),
    .A2(\decoded_imm[20] ),
    .B1(_04168_),
    .B2(_14231_),
    .X(_04169_));
 sky130_fd_sc_hd__o22a_1 _19463_ (.A1(_04163_),
    .A2(_13898_),
    .B1(_04164_),
    .B2(_04165_),
    .X(_04170_));
 sky130_fd_sc_hd__a2bb2oi_1 _19464_ (.A1_N(_04169_),
    .A2_N(_04170_),
    .B1(_04169_),
    .B2(_04170_),
    .Y(_01431_));
 sky130_vsdinv _19465_ (.A(\reg_pc[21] ),
    .Y(_04171_));
 sky130_fd_sc_hd__buf_1 _19466_ (.A(_04171_),
    .X(_04172_));
 sky130_fd_sc_hd__buf_1 _19467_ (.A(_04121_),
    .X(_04173_));
 sky130_fd_sc_hd__nor2_1 _19468_ (.A(_04172_),
    .B(_04173_),
    .Y(_01432_));
 sky130_vsdinv _19469_ (.A(net319),
    .Y(_04174_));
 sky130_fd_sc_hd__clkbuf_2 _19470_ (.A(_04174_),
    .X(_04175_));
 sky130_fd_sc_hd__a22o_1 _19471_ (.A1(_13424_),
    .A2(\decoded_imm[21] ),
    .B1(_04175_),
    .B2(_14233_),
    .X(_04176_));
 sky130_fd_sc_hd__o22a_1 _19472_ (.A1(_04168_),
    .A2(_14231_),
    .B1(_04169_),
    .B2(_04170_),
    .X(_04177_));
 sky130_fd_sc_hd__a2bb2oi_1 _19473_ (.A1_N(_04176_),
    .A2_N(_04177_),
    .B1(_04176_),
    .B2(_04177_),
    .Y(_01434_));
 sky130_vsdinv _19474_ (.A(\reg_pc[22] ),
    .Y(_04178_));
 sky130_fd_sc_hd__nor2_1 _19475_ (.A(_04178_),
    .B(_04173_),
    .Y(_01435_));
 sky130_vsdinv _19476_ (.A(net320),
    .Y(_04179_));
 sky130_fd_sc_hd__clkbuf_2 _19477_ (.A(_04179_),
    .X(_04180_));
 sky130_fd_sc_hd__a22o_1 _19478_ (.A1(_13422_),
    .A2(\decoded_imm[22] ),
    .B1(_04180_),
    .B2(_14235_),
    .X(_04181_));
 sky130_fd_sc_hd__o22a_1 _19479_ (.A1(_04175_),
    .A2(_14233_),
    .B1(_04176_),
    .B2(_04177_),
    .X(_04182_));
 sky130_fd_sc_hd__a2bb2oi_1 _19480_ (.A1_N(_04181_),
    .A2_N(_04182_),
    .B1(_04181_),
    .B2(_04182_),
    .Y(_01437_));
 sky130_vsdinv _19481_ (.A(\reg_pc[23] ),
    .Y(_04183_));
 sky130_fd_sc_hd__clkbuf_2 _19482_ (.A(_04183_),
    .X(_04184_));
 sky130_fd_sc_hd__nor2_1 _19483_ (.A(_04184_),
    .B(_04173_),
    .Y(_01438_));
 sky130_vsdinv _19484_ (.A(net321),
    .Y(_04185_));
 sky130_fd_sc_hd__buf_2 _19485_ (.A(_04185_),
    .X(_04186_));
 sky130_fd_sc_hd__a22o_1 _19486_ (.A1(_13419_),
    .A2(\decoded_imm[23] ),
    .B1(_04186_),
    .B2(_14237_),
    .X(_04187_));
 sky130_fd_sc_hd__o22a_2 _19487_ (.A1(_04180_),
    .A2(_14235_),
    .B1(_04181_),
    .B2(_04182_),
    .X(_04188_));
 sky130_fd_sc_hd__a2bb2oi_1 _19488_ (.A1_N(_04187_),
    .A2_N(_04188_),
    .B1(_04187_),
    .B2(_04188_),
    .Y(_01440_));
 sky130_vsdinv _19489_ (.A(\reg_pc[24] ),
    .Y(_04189_));
 sky130_fd_sc_hd__clkbuf_2 _19490_ (.A(_04189_),
    .X(_04190_));
 sky130_fd_sc_hd__nor2_1 _19491_ (.A(_04190_),
    .B(_04173_),
    .Y(_01441_));
 sky130_fd_sc_hd__o22ai_4 _19492_ (.A1(_04186_),
    .A2(_14237_),
    .B1(_04187_),
    .B2(_04188_),
    .Y(_04191_));
 sky130_vsdinv _19493_ (.A(net322),
    .Y(_04192_));
 sky130_fd_sc_hd__o22a_1 _19494_ (.A1(_04192_),
    .A2(_14240_),
    .B1(_13415_),
    .B2(_13925_),
    .X(_04193_));
 sky130_fd_sc_hd__o2bb2a_1 _19495_ (.A1_N(_04191_),
    .A2_N(_04193_),
    .B1(_04191_),
    .B2(_04193_),
    .X(_01443_));
 sky130_vsdinv _19496_ (.A(\reg_pc[25] ),
    .Y(_04194_));
 sky130_fd_sc_hd__clkbuf_2 _19497_ (.A(_04121_),
    .X(_04195_));
 sky130_fd_sc_hd__nor2_1 _19498_ (.A(_04194_),
    .B(_04195_),
    .Y(_01444_));
 sky130_fd_sc_hd__nor2_1 _19499_ (.A(_13413_),
    .B(_13927_),
    .Y(_04196_));
 sky130_fd_sc_hd__a21oi_2 _19500_ (.A1(_13414_),
    .A2(_13927_),
    .B1(_04196_),
    .Y(_04197_));
 sky130_fd_sc_hd__a22o_1 _19501_ (.A1(_13417_),
    .A2(_13925_),
    .B1(_04191_),
    .B2(_04193_),
    .X(_04198_));
 sky130_fd_sc_hd__a2bb2oi_1 _19502_ (.A1_N(_04197_),
    .A2_N(_04198_),
    .B1(_04197_),
    .B2(_04198_),
    .Y(_01446_));
 sky130_vsdinv _19503_ (.A(\reg_pc[26] ),
    .Y(_04199_));
 sky130_fd_sc_hd__buf_1 _19504_ (.A(_04199_),
    .X(_04200_));
 sky130_fd_sc_hd__nor2_1 _19505_ (.A(_04200_),
    .B(_04195_),
    .Y(_01447_));
 sky130_fd_sc_hd__buf_1 _19506_ (.A(_13413_),
    .X(_04201_));
 sky130_vsdinv _19507_ (.A(_04201_),
    .Y(_04202_));
 sky130_fd_sc_hd__o32a_1 _19508_ (.A1(_04192_),
    .A2(_14240_),
    .A3(_04196_),
    .B1(_04202_),
    .B2(_14241_),
    .X(_04203_));
 sky130_vsdinv _19509_ (.A(_04203_),
    .Y(_04204_));
 sky130_fd_sc_hd__a31o_1 _19510_ (.A1(_04193_),
    .A2(_04197_),
    .A3(_04191_),
    .B1(_04204_),
    .X(_04205_));
 sky130_vsdinv _19511_ (.A(_13410_),
    .Y(_04206_));
 sky130_fd_sc_hd__o22a_1 _19512_ (.A1(_04206_),
    .A2(_14243_),
    .B1(_13411_),
    .B2(_13931_),
    .X(_04207_));
 sky130_fd_sc_hd__o2bb2a_1 _19513_ (.A1_N(_04205_),
    .A2_N(_04207_),
    .B1(_04205_),
    .B2(_04207_),
    .X(_01449_));
 sky130_vsdinv _19514_ (.A(\reg_pc[27] ),
    .Y(_04208_));
 sky130_fd_sc_hd__nor2_1 _19515_ (.A(_04208_),
    .B(_04195_),
    .Y(_01450_));
 sky130_fd_sc_hd__nor2_2 _19516_ (.A(_13407_),
    .B(_13933_),
    .Y(_04209_));
 sky130_fd_sc_hd__a21oi_2 _19517_ (.A1(_13408_),
    .A2(_13933_),
    .B1(_04209_),
    .Y(_04210_));
 sky130_fd_sc_hd__a22o_1 _19518_ (.A1(_13412_),
    .A2(_13931_),
    .B1(_04205_),
    .B2(_04207_),
    .X(_04211_));
 sky130_fd_sc_hd__a2bb2oi_1 _19519_ (.A1_N(_04210_),
    .A2_N(_04211_),
    .B1(_04210_),
    .B2(_04211_),
    .Y(_01452_));
 sky130_vsdinv _19520_ (.A(\reg_pc[28] ),
    .Y(_04212_));
 sky130_fd_sc_hd__nor2_1 _19521_ (.A(_04212_),
    .B(_04195_),
    .Y(_01453_));
 sky130_fd_sc_hd__buf_1 _19522_ (.A(net325),
    .X(_04213_));
 sky130_vsdinv _19523_ (.A(_04213_),
    .Y(_04214_));
 sky130_fd_sc_hd__o32a_1 _19524_ (.A1(_04206_),
    .A2(_14243_),
    .A3(_04209_),
    .B1(_04214_),
    .B2(_14244_),
    .X(_04215_));
 sky130_vsdinv _19525_ (.A(_04215_),
    .Y(_04216_));
 sky130_fd_sc_hd__a31o_1 _19526_ (.A1(_04207_),
    .A2(_04210_),
    .A3(_04205_),
    .B1(_04216_),
    .X(_04217_));
 sky130_fd_sc_hd__nor2_1 _19527_ (.A(_13404_),
    .B(_13935_),
    .Y(_04218_));
 sky130_fd_sc_hd__a21oi_1 _19528_ (.A1(_13405_),
    .A2(_13935_),
    .B1(_04218_),
    .Y(_04219_));
 sky130_vsdinv _19529_ (.A(_04217_),
    .Y(_04220_));
 sky130_vsdinv _19530_ (.A(_04219_),
    .Y(_04221_));
 sky130_fd_sc_hd__o22a_1 _19531_ (.A1(_04217_),
    .A2(_04219_),
    .B1(_04220_),
    .B2(_04221_),
    .X(_01455_));
 sky130_vsdinv _19532_ (.A(\reg_pc[29] ),
    .Y(_04222_));
 sky130_fd_sc_hd__nor2_1 _19533_ (.A(_04222_),
    .B(_14250_),
    .Y(_01456_));
 sky130_vsdinv _19534_ (.A(_13404_),
    .Y(_04223_));
 sky130_fd_sc_hd__o22a_1 _19535_ (.A1(_04223_),
    .A2(_14246_),
    .B1(_04220_),
    .B2(_04218_),
    .X(_04224_));
 sky130_fd_sc_hd__nor2_1 _19536_ (.A(_13401_),
    .B(_13937_),
    .Y(_04225_));
 sky130_fd_sc_hd__a21o_1 _19537_ (.A1(_13402_),
    .A2(_13937_),
    .B1(_04225_),
    .X(_04226_));
 sky130_fd_sc_hd__o2bb2a_1 _19538_ (.A1_N(_04224_),
    .A2_N(_04226_),
    .B1(_04224_),
    .B2(_04226_),
    .X(_01458_));
 sky130_vsdinv _19539_ (.A(\reg_pc[30] ),
    .Y(_04227_));
 sky130_fd_sc_hd__nor2_1 _19540_ (.A(_04227_),
    .B(_14250_),
    .Y(_01459_));
 sky130_vsdinv _19541_ (.A(_13398_),
    .Y(_04228_));
 sky130_fd_sc_hd__a22o_1 _19542_ (.A1(_13399_),
    .A2(\decoded_imm[30] ),
    .B1(_04228_),
    .B2(_14249_),
    .X(_04229_));
 sky130_vsdinv _19543_ (.A(_13400_),
    .Y(_04230_));
 sky130_fd_sc_hd__o22a_1 _19544_ (.A1(_04230_),
    .A2(_14247_),
    .B1(_04224_),
    .B2(_04225_),
    .X(_04231_));
 sky130_fd_sc_hd__a2bb2oi_1 _19545_ (.A1_N(_04229_),
    .A2_N(_04231_),
    .B1(_04229_),
    .B2(_04231_),
    .Y(_01461_));
 sky130_vsdinv _19546_ (.A(\reg_pc[31] ),
    .Y(_04232_));
 sky130_fd_sc_hd__nor2_1 _19547_ (.A(_04232_),
    .B(_14250_),
    .Y(_01462_));
 sky130_fd_sc_hd__buf_1 _19548_ (.A(_04228_),
    .X(_04233_));
 sky130_fd_sc_hd__o22a_1 _19549_ (.A1(_04233_),
    .A2(_14249_),
    .B1(_04229_),
    .B2(_04231_),
    .X(_04234_));
 sky130_fd_sc_hd__o22a_1 _19550_ (.A1(_11682_),
    .A2(\decoded_imm[31] ),
    .B1(_11684_),
    .B2(_13940_),
    .X(_04235_));
 sky130_fd_sc_hd__o2bb2ai_1 _19551_ (.A1_N(_04234_),
    .A2_N(_04235_),
    .B1(_04234_),
    .B2(_04235_),
    .Y(_01464_));
 sky130_fd_sc_hd__and2_1 _19552_ (.A(_14168_),
    .B(_01466_),
    .X(_01467_));
 sky130_fd_sc_hd__and2_1 _19553_ (.A(_14168_),
    .B(_01469_),
    .X(_01470_));
 sky130_vsdinv _19554_ (.A(\reg_next_pc[4] ),
    .Y(_01471_));
 sky130_fd_sc_hd__a21oi_1 _19555_ (.A1(_14168_),
    .A2(_01473_),
    .B1(_11785_),
    .Y(_01474_));
 sky130_fd_sc_hd__buf_2 _19556_ (.A(_11575_),
    .X(_04236_));
 sky130_fd_sc_hd__buf_1 _19557_ (.A(_04236_),
    .X(_04237_));
 sky130_fd_sc_hd__and2_1 _19558_ (.A(_04237_),
    .B(_01477_),
    .X(_01478_));
 sky130_fd_sc_hd__and2_1 _19559_ (.A(_04237_),
    .B(_01480_),
    .X(_01481_));
 sky130_fd_sc_hd__and2_1 _19560_ (.A(_04237_),
    .B(_01483_),
    .X(_01484_));
 sky130_fd_sc_hd__and2_1 _19561_ (.A(_04237_),
    .B(_01486_),
    .X(_01487_));
 sky130_fd_sc_hd__buf_1 _19562_ (.A(_04236_),
    .X(_04238_));
 sky130_fd_sc_hd__and2_1 _19563_ (.A(_04238_),
    .B(_01489_),
    .X(_01490_));
 sky130_fd_sc_hd__and2_1 _19564_ (.A(_04238_),
    .B(_01492_),
    .X(_01493_));
 sky130_fd_sc_hd__and2_1 _19565_ (.A(_04238_),
    .B(_01495_),
    .X(_01496_));
 sky130_fd_sc_hd__and2_1 _19566_ (.A(_04238_),
    .B(_01498_),
    .X(_01499_));
 sky130_fd_sc_hd__buf_1 _19567_ (.A(_04236_),
    .X(_04239_));
 sky130_fd_sc_hd__and2_1 _19568_ (.A(_04239_),
    .B(_01501_),
    .X(_01502_));
 sky130_fd_sc_hd__and2_1 _19569_ (.A(_04239_),
    .B(_01504_),
    .X(_01505_));
 sky130_fd_sc_hd__and2_1 _19570_ (.A(_04239_),
    .B(_01507_),
    .X(_01508_));
 sky130_fd_sc_hd__and2_1 _19571_ (.A(_04239_),
    .B(_01510_),
    .X(_01511_));
 sky130_fd_sc_hd__buf_1 _19572_ (.A(_04236_),
    .X(_04240_));
 sky130_fd_sc_hd__and2_1 _19573_ (.A(_04240_),
    .B(_01513_),
    .X(_01514_));
 sky130_fd_sc_hd__and2_1 _19574_ (.A(_04240_),
    .B(_01516_),
    .X(_01517_));
 sky130_fd_sc_hd__and2_1 _19575_ (.A(_04240_),
    .B(_01519_),
    .X(_01520_));
 sky130_fd_sc_hd__and2_1 _19576_ (.A(_04240_),
    .B(_01522_),
    .X(_01523_));
 sky130_fd_sc_hd__buf_1 _19577_ (.A(_13779_),
    .X(_04241_));
 sky130_fd_sc_hd__and2_1 _19578_ (.A(_04241_),
    .B(_01525_),
    .X(_01526_));
 sky130_fd_sc_hd__and2_1 _19579_ (.A(_04241_),
    .B(_01528_),
    .X(_01529_));
 sky130_fd_sc_hd__and2_1 _19580_ (.A(_04241_),
    .B(_01531_),
    .X(_01532_));
 sky130_fd_sc_hd__and2_1 _19581_ (.A(_04241_),
    .B(_01534_),
    .X(_01535_));
 sky130_fd_sc_hd__buf_1 _19582_ (.A(_13779_),
    .X(_04242_));
 sky130_fd_sc_hd__and2_1 _19583_ (.A(_04242_),
    .B(_01537_),
    .X(_01538_));
 sky130_fd_sc_hd__and2_1 _19584_ (.A(_04242_),
    .B(_01540_),
    .X(_01541_));
 sky130_fd_sc_hd__and2_1 _19585_ (.A(_04242_),
    .B(_01543_),
    .X(_01544_));
 sky130_fd_sc_hd__and2_1 _19586_ (.A(_04242_),
    .B(_01546_),
    .X(_01547_));
 sky130_fd_sc_hd__and2_1 _19587_ (.A(_11576_),
    .B(_01549_),
    .X(_01550_));
 sky130_fd_sc_hd__and2_1 _19588_ (.A(_11576_),
    .B(_01552_),
    .X(_01553_));
 sky130_fd_sc_hd__and2_1 _19589_ (.A(_11576_),
    .B(_01555_),
    .X(_01556_));
 sky130_vsdinv _19590_ (.A(_02590_),
    .Y(_04243_));
 sky130_fd_sc_hd__nor2_2 _19591_ (.A(_04243_),
    .B(_13794_),
    .Y(_04244_));
 sky130_fd_sc_hd__a21oi_1 _19592_ (.A1(_04243_),
    .A2(_13794_),
    .B1(_04244_),
    .Y(_01557_));
 sky130_vsdinv _19593_ (.A(_02560_),
    .Y(_04245_));
 sky130_fd_sc_hd__buf_1 _19594_ (.A(_04245_),
    .X(_01561_));
 sky130_fd_sc_hd__o22a_1 _19595_ (.A1(_04245_),
    .A2(_13801_),
    .B1(_12083_),
    .B2(\decoded_imm_uj[2] ),
    .X(_04246_));
 sky130_fd_sc_hd__o2bb2a_1 _19596_ (.A1_N(_04244_),
    .A2_N(_04246_),
    .B1(_04244_),
    .B2(_04246_),
    .X(_01562_));
 sky130_fd_sc_hd__o22a_1 _19597_ (.A1(_01561_),
    .A2(_02410_),
    .B1(_12083_),
    .B2(_12384_),
    .X(_01565_));
 sky130_vsdinv _19598_ (.A(_02571_),
    .Y(_04247_));
 sky130_fd_sc_hd__nor2_2 _19599_ (.A(_04247_),
    .B(_01561_),
    .Y(_04248_));
 sky130_fd_sc_hd__a21oi_1 _19600_ (.A1(_04247_),
    .A2(_01561_),
    .B1(_04248_),
    .Y(_01567_));
 sky130_fd_sc_hd__a22o_1 _19601_ (.A1(_12083_),
    .A2(\decoded_imm_uj[2] ),
    .B1(_04244_),
    .B2(_04246_),
    .X(_04249_));
 sky130_fd_sc_hd__nor2_1 _19602_ (.A(_02571_),
    .B(\decoded_imm_uj[3] ),
    .Y(_04250_));
 sky130_fd_sc_hd__a21oi_1 _19603_ (.A1(_02571_),
    .A2(\decoded_imm_uj[3] ),
    .B1(_04250_),
    .Y(_04251_));
 sky130_vsdinv _19604_ (.A(_04249_),
    .Y(_04252_));
 sky130_vsdinv _19605_ (.A(_04251_),
    .Y(_04253_));
 sky130_fd_sc_hd__o22a_1 _19606_ (.A1(_04249_),
    .A2(_04251_),
    .B1(_04252_),
    .B2(_04253_),
    .X(_01568_));
 sky130_fd_sc_hd__nand2_1 _19607_ (.A(_12082_),
    .B(_04248_),
    .Y(_04254_));
 sky130_fd_sc_hd__o21a_1 _19608_ (.A1(_02582_),
    .A2(_04248_),
    .B1(_04254_),
    .X(_01571_));
 sky130_fd_sc_hd__o22a_1 _19609_ (.A1(_04247_),
    .A2(_13808_),
    .B1(_04252_),
    .B2(_04250_),
    .X(_04255_));
 sky130_vsdinv _19610_ (.A(_04255_),
    .Y(_04256_));
 sky130_fd_sc_hd__nor2_1 _19611_ (.A(\decoded_imm_uj[4] ),
    .B(_12082_),
    .Y(_04257_));
 sky130_fd_sc_hd__a21o_1 _19612_ (.A1(\decoded_imm_uj[4] ),
    .A2(_02582_),
    .B1(_04257_),
    .X(_04258_));
 sky130_fd_sc_hd__a2bb2o_1 _19613_ (.A1_N(_04256_),
    .A2_N(_04258_),
    .B1(_04256_),
    .B2(_04258_),
    .X(_01572_));
 sky130_vsdinv _19614_ (.A(_02583_),
    .Y(_04259_));
 sky130_fd_sc_hd__nor2_2 _19615_ (.A(_04259_),
    .B(_04254_),
    .Y(_04260_));
 sky130_fd_sc_hd__a21oi_1 _19616_ (.A1(_04259_),
    .A2(_04254_),
    .B1(_04260_),
    .Y(_01575_));
 sky130_fd_sc_hd__o22a_1 _19617_ (.A1(_00367_),
    .A2(_01475_),
    .B1(_04255_),
    .B2(_04257_),
    .X(_04261_));
 sky130_fd_sc_hd__nor2_1 _19618_ (.A(_02583_),
    .B(\decoded_imm_uj[5] ),
    .Y(_04262_));
 sky130_fd_sc_hd__a21o_1 _19619_ (.A1(_02583_),
    .A2(\decoded_imm_uj[5] ),
    .B1(_04262_),
    .X(_04263_));
 sky130_fd_sc_hd__o2bb2a_1 _19620_ (.A1_N(_04261_),
    .A2_N(_04263_),
    .B1(_04261_),
    .B2(_04263_),
    .X(_01576_));
 sky130_fd_sc_hd__nand2_1 _19621_ (.A(_02584_),
    .B(_04260_),
    .Y(_04264_));
 sky130_fd_sc_hd__o21a_1 _19622_ (.A1(_12077_),
    .A2(_04260_),
    .B1(_04264_),
    .X(_01579_));
 sky130_fd_sc_hd__o22a_1 _19623_ (.A1(_04259_),
    .A2(_13819_),
    .B1(_04261_),
    .B2(_04262_),
    .X(_04265_));
 sky130_fd_sc_hd__nor2_1 _19624_ (.A(_02584_),
    .B(\decoded_imm_uj[6] ),
    .Y(_04266_));
 sky130_fd_sc_hd__a21o_1 _19625_ (.A1(_12077_),
    .A2(_13272_),
    .B1(_04266_),
    .X(_04267_));
 sky130_fd_sc_hd__o2bb2a_1 _19626_ (.A1_N(_04265_),
    .A2_N(_04267_),
    .B1(_04265_),
    .B2(_04267_),
    .X(_01580_));
 sky130_vsdinv _19627_ (.A(_02585_),
    .Y(_04268_));
 sky130_fd_sc_hd__or2_1 _19628_ (.A(_04268_),
    .B(_04264_),
    .X(_04269_));
 sky130_vsdinv _19629_ (.A(_04269_),
    .Y(_04270_));
 sky130_fd_sc_hd__a21oi_1 _19630_ (.A1(_04268_),
    .A2(_04264_),
    .B1(_04270_),
    .Y(_01583_));
 sky130_fd_sc_hd__o2bb2a_1 _19631_ (.A1_N(_12077_),
    .A2_N(_13272_),
    .B1(_04265_),
    .B2(_04266_),
    .X(_04271_));
 sky130_fd_sc_hd__nor2_1 _19632_ (.A(_02585_),
    .B(\decoded_imm_uj[7] ),
    .Y(_04272_));
 sky130_fd_sc_hd__a21o_1 _19633_ (.A1(_02585_),
    .A2(\decoded_imm_uj[7] ),
    .B1(_04272_),
    .X(_04273_));
 sky130_fd_sc_hd__o2bb2a_1 _19634_ (.A1_N(_04271_),
    .A2_N(_04273_),
    .B1(_04271_),
    .B2(_04273_),
    .X(_01584_));
 sky130_vsdinv _19635_ (.A(_02586_),
    .Y(_04274_));
 sky130_fd_sc_hd__or2_1 _19636_ (.A(_04274_),
    .B(_04269_),
    .X(_04275_));
 sky130_fd_sc_hd__o21a_1 _19637_ (.A1(_12074_),
    .A2(_04270_),
    .B1(_04275_),
    .X(_01587_));
 sky130_fd_sc_hd__o22a_1 _19638_ (.A1(_04268_),
    .A2(_13829_),
    .B1(_04271_),
    .B2(_04272_),
    .X(_04276_));
 sky130_fd_sc_hd__nor2_1 _19639_ (.A(_12074_),
    .B(\decoded_imm_uj[8] ),
    .Y(_04277_));
 sky130_fd_sc_hd__a21o_1 _19640_ (.A1(_12074_),
    .A2(\decoded_imm_uj[8] ),
    .B1(_04277_),
    .X(_04278_));
 sky130_fd_sc_hd__o2bb2a_1 _19641_ (.A1_N(_04276_),
    .A2_N(_04278_),
    .B1(_04276_),
    .B2(_04278_),
    .X(_01588_));
 sky130_vsdinv _19642_ (.A(_02587_),
    .Y(_04279_));
 sky130_fd_sc_hd__or2_1 _19643_ (.A(_04279_),
    .B(_04275_),
    .X(_04280_));
 sky130_vsdinv _19644_ (.A(_04280_),
    .Y(_04281_));
 sky130_fd_sc_hd__a21oi_1 _19645_ (.A1(_04279_),
    .A2(_04275_),
    .B1(_04281_),
    .Y(_01591_));
 sky130_fd_sc_hd__o22a_1 _19646_ (.A1(_04274_),
    .A2(_13835_),
    .B1(_04276_),
    .B2(_04277_),
    .X(_04282_));
 sky130_fd_sc_hd__nor2_1 _19647_ (.A(_02587_),
    .B(\decoded_imm_uj[9] ),
    .Y(_04283_));
 sky130_fd_sc_hd__a21o_1 _19648_ (.A1(_02587_),
    .A2(\decoded_imm_uj[9] ),
    .B1(_04283_),
    .X(_04284_));
 sky130_fd_sc_hd__o2bb2a_1 _19649_ (.A1_N(_04282_),
    .A2_N(_04284_),
    .B1(_04282_),
    .B2(_04284_),
    .X(_01592_));
 sky130_vsdinv _19650_ (.A(_02588_),
    .Y(_04285_));
 sky130_fd_sc_hd__or2_1 _19651_ (.A(_04285_),
    .B(_04280_),
    .X(_04286_));
 sky130_fd_sc_hd__o21a_1 _19652_ (.A1(_12071_),
    .A2(_04281_),
    .B1(_04286_),
    .X(_01595_));
 sky130_fd_sc_hd__o22a_1 _19653_ (.A1(_04279_),
    .A2(_13840_),
    .B1(_04282_),
    .B2(_04283_),
    .X(_04287_));
 sky130_fd_sc_hd__nor2_1 _19654_ (.A(_12071_),
    .B(\decoded_imm_uj[10] ),
    .Y(_04288_));
 sky130_fd_sc_hd__a21o_1 _19655_ (.A1(_12071_),
    .A2(\decoded_imm_uj[10] ),
    .B1(_04288_),
    .X(_04289_));
 sky130_fd_sc_hd__o2bb2a_1 _19656_ (.A1_N(_04287_),
    .A2_N(_04289_),
    .B1(_04287_),
    .B2(_04289_),
    .X(_01596_));
 sky130_vsdinv _19657_ (.A(_02589_),
    .Y(_04290_));
 sky130_fd_sc_hd__or2_1 _19658_ (.A(_04290_),
    .B(_04286_),
    .X(_04291_));
 sky130_vsdinv _19659_ (.A(_04291_),
    .Y(_04292_));
 sky130_fd_sc_hd__a21oi_1 _19660_ (.A1(_04290_),
    .A2(_04286_),
    .B1(_04292_),
    .Y(_01599_));
 sky130_fd_sc_hd__a22o_1 _19661_ (.A1(_02589_),
    .A2(\decoded_imm_uj[11] ),
    .B1(_04290_),
    .B2(_13850_),
    .X(_04293_));
 sky130_fd_sc_hd__o22a_1 _19662_ (.A1(_04285_),
    .A2(_13846_),
    .B1(_04287_),
    .B2(_04288_),
    .X(_04294_));
 sky130_fd_sc_hd__a2bb2oi_1 _19663_ (.A1_N(_04293_),
    .A2_N(_04294_),
    .B1(_04293_),
    .B2(_04294_),
    .Y(_01600_));
 sky130_vsdinv _19664_ (.A(_02561_),
    .Y(_04295_));
 sky130_fd_sc_hd__or2_1 _19665_ (.A(_04295_),
    .B(_04291_),
    .X(_04296_));
 sky130_fd_sc_hd__o21a_1 _19666_ (.A1(_02561_),
    .A2(_04292_),
    .B1(_04296_),
    .X(_01603_));
 sky130_fd_sc_hd__a22o_1 _19667_ (.A1(_02561_),
    .A2(\decoded_imm_uj[12] ),
    .B1(_04295_),
    .B2(_13857_),
    .X(_04297_));
 sky130_fd_sc_hd__o22a_1 _19668_ (.A1(_04290_),
    .A2(_13850_),
    .B1(_04293_),
    .B2(_04294_),
    .X(_04298_));
 sky130_fd_sc_hd__a2bb2oi_1 _19669_ (.A1_N(_04297_),
    .A2_N(_04298_),
    .B1(_04297_),
    .B2(_04298_),
    .Y(_01604_));
 sky130_vsdinv _19670_ (.A(_02562_),
    .Y(_04299_));
 sky130_fd_sc_hd__or2_1 _19671_ (.A(_04299_),
    .B(_04296_),
    .X(_04300_));
 sky130_vsdinv _19672_ (.A(_04300_),
    .Y(_04301_));
 sky130_fd_sc_hd__a21oi_1 _19673_ (.A1(_04299_),
    .A2(_04296_),
    .B1(_04301_),
    .Y(_01607_));
 sky130_fd_sc_hd__a22o_1 _19674_ (.A1(_02562_),
    .A2(\decoded_imm_uj[13] ),
    .B1(_04299_),
    .B2(_13865_),
    .X(_04302_));
 sky130_fd_sc_hd__o22a_1 _19675_ (.A1(_04295_),
    .A2(_13857_),
    .B1(_04297_),
    .B2(_04298_),
    .X(_04303_));
 sky130_fd_sc_hd__a2bb2oi_1 _19676_ (.A1_N(_04302_),
    .A2_N(_04303_),
    .B1(_04302_),
    .B2(_04303_),
    .Y(_01608_));
 sky130_vsdinv _19677_ (.A(_02563_),
    .Y(_04304_));
 sky130_fd_sc_hd__or2_1 _19678_ (.A(_04304_),
    .B(_04300_),
    .X(_04305_));
 sky130_fd_sc_hd__o21a_1 _19679_ (.A1(_02563_),
    .A2(_04301_),
    .B1(_04305_),
    .X(_01611_));
 sky130_fd_sc_hd__a22o_1 _19680_ (.A1(_02563_),
    .A2(\decoded_imm_uj[14] ),
    .B1(_04304_),
    .B2(_13871_),
    .X(_04306_));
 sky130_fd_sc_hd__o22a_1 _19681_ (.A1(_04299_),
    .A2(_13865_),
    .B1(_04302_),
    .B2(_04303_),
    .X(_04307_));
 sky130_fd_sc_hd__a2bb2oi_1 _19682_ (.A1_N(_04306_),
    .A2_N(_04307_),
    .B1(_04306_),
    .B2(_04307_),
    .Y(_01612_));
 sky130_vsdinv _19683_ (.A(_02564_),
    .Y(_04308_));
 sky130_fd_sc_hd__or2_1 _19684_ (.A(_04308_),
    .B(_04305_),
    .X(_04309_));
 sky130_vsdinv _19685_ (.A(_04309_),
    .Y(_04310_));
 sky130_fd_sc_hd__a21oi_1 _19686_ (.A1(_04308_),
    .A2(_04305_),
    .B1(_04310_),
    .Y(_01615_));
 sky130_fd_sc_hd__a22o_1 _19687_ (.A1(_02564_),
    .A2(\decoded_imm_uj[15] ),
    .B1(_04308_),
    .B2(_13875_),
    .X(_04311_));
 sky130_fd_sc_hd__o22a_1 _19688_ (.A1(_04304_),
    .A2(_13871_),
    .B1(_04306_),
    .B2(_04307_),
    .X(_04312_));
 sky130_fd_sc_hd__a2bb2oi_1 _19689_ (.A1_N(_04311_),
    .A2_N(_04312_),
    .B1(_04311_),
    .B2(_04312_),
    .Y(_01616_));
 sky130_vsdinv _19690_ (.A(_02565_),
    .Y(_04313_));
 sky130_fd_sc_hd__or2_1 _19691_ (.A(_04313_),
    .B(_04309_),
    .X(_04314_));
 sky130_fd_sc_hd__o21a_1 _19692_ (.A1(_02565_),
    .A2(_04310_),
    .B1(_04314_),
    .X(_01619_));
 sky130_fd_sc_hd__a22o_1 _19693_ (.A1(_02565_),
    .A2(\decoded_imm_uj[16] ),
    .B1(_04313_),
    .B2(_13883_),
    .X(_04315_));
 sky130_fd_sc_hd__o22a_1 _19694_ (.A1(_04308_),
    .A2(_13875_),
    .B1(_04311_),
    .B2(_04312_),
    .X(_04316_));
 sky130_fd_sc_hd__a2bb2oi_1 _19695_ (.A1_N(_04315_),
    .A2_N(_04316_),
    .B1(_04315_),
    .B2(_04316_),
    .Y(_01620_));
 sky130_vsdinv _19696_ (.A(_02566_),
    .Y(_04317_));
 sky130_fd_sc_hd__or2_1 _19697_ (.A(_04317_),
    .B(_04314_),
    .X(_04318_));
 sky130_vsdinv _19698_ (.A(_04318_),
    .Y(_04319_));
 sky130_fd_sc_hd__a21oi_1 _19699_ (.A1(_04317_),
    .A2(_04314_),
    .B1(_04319_),
    .Y(_01623_));
 sky130_fd_sc_hd__a22o_1 _19700_ (.A1(_02566_),
    .A2(\decoded_imm_uj[17] ),
    .B1(_04317_),
    .B2(_13888_),
    .X(_04320_));
 sky130_fd_sc_hd__o22a_1 _19701_ (.A1(_04313_),
    .A2(_13883_),
    .B1(_04315_),
    .B2(_04316_),
    .X(_04321_));
 sky130_fd_sc_hd__a2bb2oi_1 _19702_ (.A1_N(_04320_),
    .A2_N(_04321_),
    .B1(_04320_),
    .B2(_04321_),
    .Y(_01624_));
 sky130_vsdinv _19703_ (.A(_02567_),
    .Y(_04322_));
 sky130_fd_sc_hd__or2_1 _19704_ (.A(_04322_),
    .B(_04318_),
    .X(_04323_));
 sky130_fd_sc_hd__o21a_1 _19705_ (.A1(_12063_),
    .A2(_04319_),
    .B1(_04323_),
    .X(_01627_));
 sky130_fd_sc_hd__o22a_1 _19706_ (.A1(_04317_),
    .A2(_13888_),
    .B1(_04320_),
    .B2(_04321_),
    .X(_04324_));
 sky130_fd_sc_hd__nor2_1 _19707_ (.A(_12063_),
    .B(\decoded_imm_uj[18] ),
    .Y(_04325_));
 sky130_fd_sc_hd__a21o_1 _19708_ (.A1(_12063_),
    .A2(\decoded_imm_uj[18] ),
    .B1(_04325_),
    .X(_04326_));
 sky130_fd_sc_hd__o2bb2a_1 _19709_ (.A1_N(_04324_),
    .A2_N(_04326_),
    .B1(_04324_),
    .B2(_04326_),
    .X(_01628_));
 sky130_vsdinv _19710_ (.A(_02568_),
    .Y(_04327_));
 sky130_fd_sc_hd__or2_1 _19711_ (.A(_04327_),
    .B(_04323_),
    .X(_04328_));
 sky130_vsdinv _19712_ (.A(_04328_),
    .Y(_04329_));
 sky130_fd_sc_hd__a21oi_1 _19713_ (.A1(_04327_),
    .A2(_04323_),
    .B1(_04329_),
    .Y(_01631_));
 sky130_fd_sc_hd__a22o_1 _19714_ (.A1(_02568_),
    .A2(\decoded_imm_uj[19] ),
    .B1(_04327_),
    .B2(_13899_),
    .X(_04330_));
 sky130_fd_sc_hd__o22a_1 _19715_ (.A1(_04322_),
    .A2(_13894_),
    .B1(_04324_),
    .B2(_04325_),
    .X(_04331_));
 sky130_fd_sc_hd__a2bb2oi_1 _19716_ (.A1_N(_04330_),
    .A2_N(_04331_),
    .B1(_04330_),
    .B2(_04331_),
    .Y(_01632_));
 sky130_vsdinv _19717_ (.A(_02569_),
    .Y(_04332_));
 sky130_fd_sc_hd__or2_1 _19718_ (.A(_04332_),
    .B(_04328_),
    .X(_04333_));
 sky130_fd_sc_hd__o21a_1 _19719_ (.A1(_12060_),
    .A2(_04329_),
    .B1(_04333_),
    .X(_01635_));
 sky130_fd_sc_hd__o22a_1 _19720_ (.A1(_04327_),
    .A2(_13899_),
    .B1(_04330_),
    .B2(_04331_),
    .X(_04334_));
 sky130_fd_sc_hd__nor2_1 _19721_ (.A(_12060_),
    .B(\decoded_imm_uj[20] ),
    .Y(_04335_));
 sky130_fd_sc_hd__a21o_1 _19722_ (.A1(_12060_),
    .A2(_13263_),
    .B1(_04335_),
    .X(_04336_));
 sky130_fd_sc_hd__o2bb2a_1 _19723_ (.A1_N(_04334_),
    .A2_N(_04336_),
    .B1(_04334_),
    .B2(_04336_),
    .X(_01636_));
 sky130_vsdinv _19724_ (.A(_02570_),
    .Y(_04337_));
 sky130_fd_sc_hd__buf_1 _19725_ (.A(_04337_),
    .X(_04338_));
 sky130_fd_sc_hd__or2_1 _19726_ (.A(_04337_),
    .B(_04333_),
    .X(_04339_));
 sky130_vsdinv _19727_ (.A(_04339_),
    .Y(_04340_));
 sky130_fd_sc_hd__a21oi_1 _19728_ (.A1(_04338_),
    .A2(_04333_),
    .B1(_04340_),
    .Y(_01639_));
 sky130_fd_sc_hd__a22o_1 _19729_ (.A1(_02570_),
    .A2(_13259_),
    .B1(_04338_),
    .B2(_13907_),
    .X(_04341_));
 sky130_fd_sc_hd__o22a_1 _19730_ (.A1(_04332_),
    .A2(_13907_),
    .B1(_04334_),
    .B2(_04335_),
    .X(_04342_));
 sky130_fd_sc_hd__or2_1 _19731_ (.A(_04341_),
    .B(_04342_),
    .X(_04343_));
 sky130_fd_sc_hd__a21boi_1 _19732_ (.A1(_04341_),
    .A2(_04342_),
    .B1_N(_04343_),
    .Y(_01640_));
 sky130_vsdinv _19733_ (.A(_02572_),
    .Y(_04344_));
 sky130_fd_sc_hd__or2_1 _19734_ (.A(_04344_),
    .B(_04339_),
    .X(_04345_));
 sky130_fd_sc_hd__o21a_1 _19735_ (.A1(_02572_),
    .A2(_04340_),
    .B1(_04345_),
    .X(_01643_));
 sky130_fd_sc_hd__o22a_1 _19736_ (.A1(_04344_),
    .A2(_13908_),
    .B1(_02572_),
    .B2(_13259_),
    .X(_04346_));
 sky130_fd_sc_hd__o21ai_1 _19737_ (.A1(_04338_),
    .A2(_13941_),
    .B1(_04343_),
    .Y(_04347_));
 sky130_vsdinv _19738_ (.A(_04346_),
    .Y(_04348_));
 sky130_vsdinv _19739_ (.A(_04347_),
    .Y(_04349_));
 sky130_fd_sc_hd__o22a_1 _19740_ (.A1(_04346_),
    .A2(_04347_),
    .B1(_04348_),
    .B2(_04349_),
    .X(_01644_));
 sky130_vsdinv _19741_ (.A(_02573_),
    .Y(_04350_));
 sky130_fd_sc_hd__or2_1 _19742_ (.A(_04350_),
    .B(_04345_),
    .X(_04351_));
 sky130_vsdinv _19743_ (.A(_04351_),
    .Y(_04352_));
 sky130_fd_sc_hd__a21oi_1 _19744_ (.A1(_04350_),
    .A2(_04345_),
    .B1(_04352_),
    .Y(_01647_));
 sky130_fd_sc_hd__buf_1 _19745_ (.A(_13908_),
    .X(_04353_));
 sky130_fd_sc_hd__o22a_1 _19746_ (.A1(_04350_),
    .A2(_04353_),
    .B1(_02573_),
    .B2(_13260_),
    .X(_04354_));
 sky130_fd_sc_hd__or2_1 _19747_ (.A(_04343_),
    .B(_04348_),
    .X(_04355_));
 sky130_fd_sc_hd__o22a_1 _19748_ (.A1(_04338_),
    .A2(_04353_),
    .B1(_04344_),
    .B2(_04353_),
    .X(_04356_));
 sky130_fd_sc_hd__nand2_1 _19749_ (.A(_04355_),
    .B(_04356_),
    .Y(_04357_));
 sky130_fd_sc_hd__o2bb2a_1 _19750_ (.A1_N(_04354_),
    .A2_N(_04357_),
    .B1(_04354_),
    .B2(_04357_),
    .X(_01648_));
 sky130_vsdinv _19751_ (.A(_02574_),
    .Y(_04358_));
 sky130_fd_sc_hd__or2_1 _19752_ (.A(_04358_),
    .B(_04351_),
    .X(_04359_));
 sky130_fd_sc_hd__o21a_1 _19753_ (.A1(_02574_),
    .A2(_04352_),
    .B1(_04359_),
    .X(_01651_));
 sky130_fd_sc_hd__o22a_1 _19754_ (.A1(_04358_),
    .A2(_13908_),
    .B1(_02574_),
    .B2(_13259_),
    .X(_04360_));
 sky130_fd_sc_hd__a22o_1 _19755_ (.A1(_02573_),
    .A2(_13262_),
    .B1(_04354_),
    .B2(_04357_),
    .X(_04361_));
 sky130_vsdinv _19756_ (.A(_04360_),
    .Y(_04362_));
 sky130_vsdinv _19757_ (.A(_04361_),
    .Y(_04363_));
 sky130_fd_sc_hd__o22a_1 _19758_ (.A1(_04360_),
    .A2(_04361_),
    .B1(_04362_),
    .B2(_04363_),
    .X(_01652_));
 sky130_vsdinv _19759_ (.A(_02575_),
    .Y(_04364_));
 sky130_fd_sc_hd__buf_1 _19760_ (.A(_04364_),
    .X(_04365_));
 sky130_fd_sc_hd__or2_1 _19761_ (.A(_04365_),
    .B(_04359_),
    .X(_04366_));
 sky130_vsdinv _19762_ (.A(_04366_),
    .Y(_04367_));
 sky130_fd_sc_hd__a21oi_1 _19763_ (.A1(_04365_),
    .A2(_04359_),
    .B1(_04367_),
    .Y(_01655_));
 sky130_fd_sc_hd__a22o_1 _19764_ (.A1(_02575_),
    .A2(_13260_),
    .B1(_04364_),
    .B2(_13909_),
    .X(_04368_));
 sky130_vsdinv _19765_ (.A(_04354_),
    .Y(_04369_));
 sky130_fd_sc_hd__o22a_1 _19766_ (.A1(_04350_),
    .A2(_13909_),
    .B1(_04358_),
    .B2(_04353_),
    .X(_04370_));
 sky130_fd_sc_hd__o311a_1 _19767_ (.A1(_04369_),
    .A2(_04362_),
    .A3(_04355_),
    .B1(_04356_),
    .C1(_04370_),
    .X(_04371_));
 sky130_fd_sc_hd__or2_1 _19768_ (.A(_04368_),
    .B(_04371_),
    .X(_04372_));
 sky130_fd_sc_hd__a21boi_1 _19769_ (.A1(_04368_),
    .A2(_04371_),
    .B1_N(_04372_),
    .Y(_01656_));
 sky130_vsdinv _19770_ (.A(_02576_),
    .Y(_04373_));
 sky130_fd_sc_hd__or2_1 _19771_ (.A(_04373_),
    .B(_04366_),
    .X(_04374_));
 sky130_fd_sc_hd__o21a_1 _19772_ (.A1(_02576_),
    .A2(_04367_),
    .B1(_04374_),
    .X(_01659_));
 sky130_fd_sc_hd__o22a_1 _19773_ (.A1(_04373_),
    .A2(_13909_),
    .B1(_02576_),
    .B2(_13260_),
    .X(_04375_));
 sky130_fd_sc_hd__o21ai_1 _19774_ (.A1(_04365_),
    .A2(_13941_),
    .B1(_04372_),
    .Y(_04376_));
 sky130_vsdinv _19775_ (.A(_04375_),
    .Y(_04377_));
 sky130_vsdinv _19776_ (.A(_04376_),
    .Y(_04378_));
 sky130_fd_sc_hd__o22a_1 _19777_ (.A1(_04375_),
    .A2(_04376_),
    .B1(_04377_),
    .B2(_04378_),
    .X(_01660_));
 sky130_vsdinv _19778_ (.A(_02577_),
    .Y(_04379_));
 sky130_fd_sc_hd__or2_1 _19779_ (.A(_04379_),
    .B(_04374_),
    .X(_04380_));
 sky130_vsdinv _19780_ (.A(_04380_),
    .Y(_04381_));
 sky130_fd_sc_hd__a21oi_1 _19781_ (.A1(_04379_),
    .A2(_04374_),
    .B1(_04381_),
    .Y(_01663_));
 sky130_fd_sc_hd__o22a_1 _19782_ (.A1(_04379_),
    .A2(_13910_),
    .B1(_02577_),
    .B2(_13261_),
    .X(_04382_));
 sky130_fd_sc_hd__or2_1 _19783_ (.A(_04372_),
    .B(_04377_),
    .X(_04383_));
 sky130_fd_sc_hd__o22a_1 _19784_ (.A1(_04365_),
    .A2(_13911_),
    .B1(_04373_),
    .B2(_13910_),
    .X(_04384_));
 sky130_fd_sc_hd__nand2_1 _19785_ (.A(_04383_),
    .B(_04384_),
    .Y(_04385_));
 sky130_fd_sc_hd__o2bb2a_1 _19786_ (.A1_N(_04382_),
    .A2_N(_04385_),
    .B1(_04382_),
    .B2(_04385_),
    .X(_01664_));
 sky130_vsdinv _19787_ (.A(_02578_),
    .Y(_04386_));
 sky130_fd_sc_hd__or2_1 _19788_ (.A(_04386_),
    .B(_04380_),
    .X(_04387_));
 sky130_fd_sc_hd__o21a_1 _19789_ (.A1(_02578_),
    .A2(_04381_),
    .B1(_04387_),
    .X(_01667_));
 sky130_fd_sc_hd__o22a_1 _19790_ (.A1(_04386_),
    .A2(_13910_),
    .B1(_02578_),
    .B2(_13261_),
    .X(_04388_));
 sky130_fd_sc_hd__a22o_1 _19791_ (.A1(_02577_),
    .A2(_13262_),
    .B1(_04382_),
    .B2(_04385_),
    .X(_04389_));
 sky130_vsdinv _19792_ (.A(_04388_),
    .Y(_04390_));
 sky130_vsdinv _19793_ (.A(_04389_),
    .Y(_04391_));
 sky130_fd_sc_hd__o22a_1 _19794_ (.A1(_04388_),
    .A2(_04389_),
    .B1(_04390_),
    .B2(_04391_),
    .X(_01668_));
 sky130_vsdinv _19795_ (.A(_02579_),
    .Y(_04392_));
 sky130_fd_sc_hd__buf_1 _19796_ (.A(_04392_),
    .X(_04393_));
 sky130_fd_sc_hd__or2_1 _19797_ (.A(_04393_),
    .B(_04387_),
    .X(_04394_));
 sky130_vsdinv _19798_ (.A(_04394_),
    .Y(_04395_));
 sky130_fd_sc_hd__a21oi_1 _19799_ (.A1(_04393_),
    .A2(_04387_),
    .B1(_04395_),
    .Y(_01671_));
 sky130_fd_sc_hd__a22o_1 _19800_ (.A1(_02579_),
    .A2(_13261_),
    .B1(_04392_),
    .B2(_13912_),
    .X(_04396_));
 sky130_vsdinv _19801_ (.A(_04382_),
    .Y(_04397_));
 sky130_fd_sc_hd__o22a_1 _19802_ (.A1(_04379_),
    .A2(_13911_),
    .B1(_04386_),
    .B2(_13911_),
    .X(_04398_));
 sky130_fd_sc_hd__o311a_1 _19803_ (.A1(_04397_),
    .A2(_04390_),
    .A3(_04383_),
    .B1(_04384_),
    .C1(_04398_),
    .X(_04399_));
 sky130_fd_sc_hd__or2_1 _19804_ (.A(_04396_),
    .B(_04399_),
    .X(_04400_));
 sky130_vsdinv _19805_ (.A(_04400_),
    .Y(_04401_));
 sky130_fd_sc_hd__a21oi_1 _19806_ (.A1(_04396_),
    .A2(_04399_),
    .B1(_04401_),
    .Y(_01672_));
 sky130_vsdinv _19807_ (.A(_02580_),
    .Y(_04402_));
 sky130_fd_sc_hd__or2_1 _19808_ (.A(_04402_),
    .B(_04394_),
    .X(_04403_));
 sky130_fd_sc_hd__o21a_1 _19809_ (.A1(_12049_),
    .A2(_04395_),
    .B1(_04403_),
    .X(_01675_));
 sky130_fd_sc_hd__clkbuf_2 _19810_ (.A(_13912_),
    .X(_04404_));
 sky130_fd_sc_hd__o22a_1 _19811_ (.A1(_12049_),
    .A2(_13263_),
    .B1(_04402_),
    .B2(_04404_),
    .X(_04405_));
 sky130_fd_sc_hd__o21ai_1 _19812_ (.A1(_04393_),
    .A2(_04404_),
    .B1(_04400_),
    .Y(_04406_));
 sky130_fd_sc_hd__a2bb2oi_1 _19813_ (.A1_N(_04405_),
    .A2_N(_04406_),
    .B1(_04405_),
    .B2(_04406_),
    .Y(_01676_));
 sky130_vsdinv _19814_ (.A(_02581_),
    .Y(_04407_));
 sky130_fd_sc_hd__a32o_1 _19815_ (.A1(_12049_),
    .A2(_04395_),
    .A3(_04407_),
    .B1(_02581_),
    .B2(_04403_),
    .X(_01679_));
 sky130_fd_sc_hd__o21ai_1 _19816_ (.A1(_02580_),
    .A2(_13262_),
    .B1(_04401_),
    .Y(_04408_));
 sky130_fd_sc_hd__o221ai_2 _19817_ (.A1(_04393_),
    .A2(_04404_),
    .B1(_04402_),
    .B2(_04404_),
    .C1(_04408_),
    .Y(_04409_));
 sky130_fd_sc_hd__a22o_1 _19818_ (.A1(_02581_),
    .A2(_13941_),
    .B1(_04407_),
    .B2(_13263_),
    .X(_04410_));
 sky130_fd_sc_hd__a2bb2oi_1 _19819_ (.A1_N(_04409_),
    .A2_N(_04410_),
    .B1(_04409_),
    .B2(_04410_),
    .Y(_01680_));
 sky130_fd_sc_hd__or2_1 _19820_ (.A(\mem_wordsize[2] ),
    .B(\mem_wordsize[1] ),
    .X(_04411_));
 sky130_vsdinv _19821_ (.A(_04411_),
    .Y(_04412_));
 sky130_fd_sc_hd__buf_8 _19822_ (.A(_04412_),
    .X(_01683_));
 sky130_fd_sc_hd__buf_1 _19823_ (.A(_14256_),
    .X(_04413_));
 sky130_fd_sc_hd__buf_2 _19824_ (.A(_04413_),
    .X(_04414_));
 sky130_fd_sc_hd__a211o_4 _19825_ (.A1(_04414_),
    .A2(\mem_wordsize[2] ),
    .B1(_04412_),
    .C1(_00304_),
    .X(net233));
 sky130_fd_sc_hd__and2_1 _19826_ (.A(net232),
    .B(net233),
    .X(_01684_));
 sky130_fd_sc_hd__and3_1 _19827_ (.A(_12013_),
    .B(_00301_),
    .C(_01685_),
    .X(_01686_));
 sky130_fd_sc_hd__buf_1 _19828_ (.A(_04411_),
    .X(_04415_));
 sky130_fd_sc_hd__or2_2 _19829_ (.A(_13486_),
    .B(_14252_),
    .X(_04416_));
 sky130_fd_sc_hd__o211a_2 _19830_ (.A1(_13486_),
    .A2(_14147_),
    .B1(_04415_),
    .C1(_04416_),
    .X(_04417_));
 sky130_fd_sc_hd__nor2_1 _19831_ (.A(_14060_),
    .B(_04417_),
    .Y(_01687_));
 sky130_fd_sc_hd__and3_1 _19832_ (.A(_12013_),
    .B(_00301_),
    .C(_01688_),
    .X(_01689_));
 sky130_fd_sc_hd__or2_2 _19833_ (.A(_04413_),
    .B(_13487_),
    .X(_04418_));
 sky130_fd_sc_hd__buf_1 _19834_ (.A(_04418_),
    .X(_04419_));
 sky130_fd_sc_hd__o211a_2 _19835_ (.A1(_04414_),
    .A2(_13985_),
    .B1(_04415_),
    .C1(_04419_),
    .X(_04420_));
 sky130_fd_sc_hd__nor2_1 _19836_ (.A(_14060_),
    .B(_04420_),
    .Y(_01690_));
 sky130_fd_sc_hd__and3_1 _19837_ (.A(_12013_),
    .B(_00301_),
    .C(_01691_),
    .X(_01692_));
 sky130_fd_sc_hd__or2_2 _19838_ (.A(_04413_),
    .B(_14252_),
    .X(_04421_));
 sky130_fd_sc_hd__o211a_2 _19839_ (.A1(_04414_),
    .A2(_13985_),
    .B1(_04415_),
    .C1(_04421_),
    .X(_04422_));
 sky130_fd_sc_hd__nor2_1 _19840_ (.A(_14060_),
    .B(_04422_),
    .Y(_01693_));
 sky130_fd_sc_hd__and3_1 _19841_ (.A(_12012_),
    .B(_11879_),
    .C(_01694_),
    .X(_01695_));
 sky130_fd_sc_hd__or2_1 _19842_ (.A(_12358_),
    .B(net12),
    .X(_04423_));
 sky130_fd_sc_hd__buf_1 _19843_ (.A(_04423_),
    .X(_01697_));
 sky130_fd_sc_hd__inv_2 _19844_ (.A(_01697_),
    .Y(_01696_));
 sky130_fd_sc_hd__nor2_1 _19845_ (.A(_12357_),
    .B(_01696_),
    .Y(_01698_));
 sky130_fd_sc_hd__and3_2 _19846_ (.A(_12551_),
    .B(_00297_),
    .C(_13945_),
    .X(_04424_));
 sky130_fd_sc_hd__nand2_8 _19847_ (.A(_14158_),
    .B(_04424_),
    .Y(_02217_));
 sky130_vsdinv _19848_ (.A(_02217_),
    .Y(_01700_));
 sky130_fd_sc_hd__o21a_1 _19849_ (.A1(_11677_),
    .A2(\irq_mask[1] ),
    .B1(_01696_),
    .X(_01701_));
 sky130_fd_sc_hd__o22ai_1 _19850_ (.A1(_01696_),
    .A2(_04424_),
    .B1(_14158_),
    .B2(_01704_),
    .Y(_01705_));
 sky130_fd_sc_hd__and2_4 _19851_ (.A(_14039_),
    .B(_00354_),
    .X(_01706_));
 sky130_vsdinv _19852_ (.A(net33),
    .Y(_01707_));
 sky130_vsdinv _19853_ (.A(net49),
    .Y(_04425_));
 sky130_fd_sc_hd__buf_1 _19854_ (.A(_04421_),
    .X(_04426_));
 sky130_vsdinv _19855_ (.A(net63),
    .Y(_01812_));
 sky130_fd_sc_hd__buf_1 _19856_ (.A(_04416_),
    .X(_04427_));
 sky130_vsdinv _19857_ (.A(net40),
    .Y(_04428_));
 sky130_fd_sc_hd__or2_1 _19858_ (.A(_04428_),
    .B(_04419_),
    .X(_04429_));
 sky130_fd_sc_hd__o221a_1 _19859_ (.A1(_04425_),
    .A2(_04426_),
    .B1(_01812_),
    .B2(_04427_),
    .C1(_04429_),
    .X(_01708_));
 sky130_vsdinv _19860_ (.A(_01710_),
    .Y(_04430_));
 sky130_fd_sc_hd__o22a_1 _19861_ (.A1(_14165_),
    .A2(_01709_),
    .B1(_14148_),
    .B2(_04430_),
    .X(_01711_));
 sky130_fd_sc_hd__buf_1 _19862_ (.A(_11741_),
    .X(_04431_));
 sky130_fd_sc_hd__buf_1 _19863_ (.A(_04431_),
    .X(_04432_));
 sky130_fd_sc_hd__buf_1 _19864_ (.A(_13344_),
    .X(_04433_));
 sky130_fd_sc_hd__or2_1 _19865_ (.A(_12147_),
    .B(_13337_),
    .X(_04434_));
 sky130_fd_sc_hd__o221a_1 _19866_ (.A1(_12115_),
    .A2(_04432_),
    .B1(_04433_),
    .B2(_12437_),
    .C1(_04434_),
    .X(_01715_));
 sky130_fd_sc_hd__buf_1 _19867_ (.A(_13300_),
    .X(_04435_));
 sky130_fd_sc_hd__buf_1 _19868_ (.A(_13307_),
    .X(_04436_));
 sky130_fd_sc_hd__o21ai_2 _19869_ (.A1(instr_setq),
    .A2(instr_getq),
    .B1(\cpuregs_rs1[0] ),
    .Y(_04437_));
 sky130_fd_sc_hd__o221a_1 _19870_ (.A1(_04435_),
    .A2(_14201_),
    .B1(_12360_),
    .B2(_04436_),
    .C1(_04437_),
    .X(_01718_));
 sky130_fd_sc_hd__buf_2 _19871_ (.A(_12280_),
    .X(_04438_));
 sky130_fd_sc_hd__o2bb2a_1 _19872_ (.A1_N(_12367_),
    .A2_N(_01713_),
    .B1(_04438_),
    .B2(_01719_),
    .X(_04439_));
 sky130_fd_sc_hd__clkbuf_4 _19873_ (.A(_11733_),
    .X(_04440_));
 sky130_fd_sc_hd__a221o_1 _19874_ (.A1(\decoded_imm[0] ),
    .A2(_13781_),
    .B1(_13278_),
    .B2(_14251_),
    .C1(_04440_),
    .X(_04441_));
 sky130_fd_sc_hd__o211ai_2 _19875_ (.A1(_14040_),
    .A2(_01712_),
    .B1(_04439_),
    .C1(_04441_),
    .Y(_01720_));
 sky130_vsdinv _19876_ (.A(net44),
    .Y(_01721_));
 sky130_vsdinv _19877_ (.A(net50),
    .Y(_04442_));
 sky130_vsdinv _19878_ (.A(net64),
    .Y(_01826_));
 sky130_vsdinv _19879_ (.A(net41),
    .Y(_04443_));
 sky130_fd_sc_hd__or2_1 _19880_ (.A(_04443_),
    .B(_04419_),
    .X(_04444_));
 sky130_fd_sc_hd__o221a_1 _19881_ (.A1(_04442_),
    .A2(_04426_),
    .B1(_01826_),
    .B2(_04427_),
    .C1(_04444_),
    .X(_01722_));
 sky130_vsdinv _19882_ (.A(_01724_),
    .Y(_04445_));
 sky130_fd_sc_hd__o22a_1 _19883_ (.A1(_14165_),
    .A2(_01723_),
    .B1(_14148_),
    .B2(_04445_),
    .X(_01725_));
 sky130_fd_sc_hd__or2_1 _19884_ (.A(_12114_),
    .B(_04431_),
    .X(_04446_));
 sky130_fd_sc_hd__o221a_1 _19885_ (.A1(_12146_),
    .A2(_13337_),
    .B1(_04433_),
    .B2(_12436_),
    .C1(_04446_),
    .X(_01729_));
 sky130_fd_sc_hd__clkbuf_2 _19886_ (.A(_11745_),
    .X(_04447_));
 sky130_fd_sc_hd__clkbuf_2 _19887_ (.A(_04447_),
    .X(_04448_));
 sky130_fd_sc_hd__buf_1 _19888_ (.A(_04448_),
    .X(_04449_));
 sky130_fd_sc_hd__nand2_1 _19889_ (.A(_04449_),
    .B(\cpuregs_rs1[1] ),
    .Y(_04450_));
 sky130_fd_sc_hd__o221a_1 _19890_ (.A1(_04435_),
    .A2(_14200_),
    .B1(_12357_),
    .B2(_04436_),
    .C1(_04450_),
    .X(_01731_));
 sky130_fd_sc_hd__a22o_1 _19891_ (.A1(\reg_pc[1] ),
    .A2(\decoded_imm[1] ),
    .B1(_14254_),
    .B2(_13790_),
    .X(_04451_));
 sky130_fd_sc_hd__or3_1 _19892_ (.A(_13277_),
    .B(_14251_),
    .C(_04451_),
    .X(_04452_));
 sky130_fd_sc_hd__o21ai_1 _19893_ (.A1(_13278_),
    .A2(_14251_),
    .B1(_04451_),
    .Y(_04453_));
 sky130_fd_sc_hd__buf_1 _19894_ (.A(_11560_),
    .X(_04454_));
 sky130_fd_sc_hd__clkbuf_4 _19895_ (.A(_04454_),
    .X(_04455_));
 sky130_fd_sc_hd__buf_1 _19896_ (.A(_12365_),
    .X(_04456_));
 sky130_fd_sc_hd__buf_2 _19897_ (.A(_11570_),
    .X(_04457_));
 sky130_fd_sc_hd__buf_1 _19898_ (.A(_04457_),
    .X(_04458_));
 sky130_fd_sc_hd__o2bb2a_1 _19899_ (.A1_N(_04456_),
    .A2_N(_01727_),
    .B1(_04458_),
    .B2(_01732_),
    .X(_04459_));
 sky130_fd_sc_hd__o21ai_1 _19900_ (.A1(_04455_),
    .A2(_01726_),
    .B1(_04459_),
    .Y(_04460_));
 sky130_fd_sc_hd__a31o_1 _19901_ (.A1(_14153_),
    .A2(_04452_),
    .A3(_04453_),
    .B1(_04460_),
    .X(_01733_));
 sky130_vsdinv _19902_ (.A(net55),
    .Y(_01734_));
 sky130_vsdinv _19903_ (.A(net51),
    .Y(_04461_));
 sky130_vsdinv _19904_ (.A(net34),
    .Y(_01839_));
 sky130_vsdinv _19905_ (.A(net42),
    .Y(_04462_));
 sky130_fd_sc_hd__or2_1 _19906_ (.A(_04462_),
    .B(_04419_),
    .X(_04463_));
 sky130_fd_sc_hd__o221a_1 _19907_ (.A1(_04461_),
    .A2(_04426_),
    .B1(_01839_),
    .B2(_04427_),
    .C1(_04463_),
    .X(_01735_));
 sky130_vsdinv _19908_ (.A(_01737_),
    .Y(_04464_));
 sky130_fd_sc_hd__o22a_1 _19909_ (.A1(_14165_),
    .A2(_01736_),
    .B1(_14148_),
    .B2(_04464_),
    .X(_01738_));
 sky130_fd_sc_hd__or2_1 _19910_ (.A(_12145_),
    .B(_13337_),
    .X(_04465_));
 sky130_fd_sc_hd__o221a_1 _19911_ (.A1(_12113_),
    .A2(_04432_),
    .B1(_04433_),
    .B2(_12435_),
    .C1(_04465_),
    .X(_01742_));
 sky130_vsdinv _19912_ (.A(\timer[2] ),
    .Y(_04466_));
 sky130_fd_sc_hd__nand2_1 _19913_ (.A(_04449_),
    .B(\cpuregs_rs1[2] ),
    .Y(_04467_));
 sky130_fd_sc_hd__o221a_1 _19914_ (.A1(_04435_),
    .A2(_04466_),
    .B1(_12354_),
    .B2(_04436_),
    .C1(_04467_),
    .X(_01744_));
 sky130_fd_sc_hd__clkbuf_1 _19915_ (.A(_12366_),
    .X(_04468_));
 sky130_fd_sc_hd__o2bb2a_1 _19916_ (.A1_N(_04468_),
    .A2_N(_01740_),
    .B1(_04438_),
    .B2(_01745_),
    .X(_04469_));
 sky130_fd_sc_hd__o21ai_1 _19917_ (.A1(_14254_),
    .A2(_13790_),
    .B1(_04452_),
    .Y(_04470_));
 sky130_fd_sc_hd__nor2_1 _19918_ (.A(\reg_pc[2] ),
    .B(_14260_),
    .Y(_04471_));
 sky130_fd_sc_hd__a21oi_1 _19919_ (.A1(\reg_pc[2] ),
    .A2(_14260_),
    .B1(_04471_),
    .Y(_04472_));
 sky130_vsdinv _19920_ (.A(_04470_),
    .Y(_04473_));
 sky130_vsdinv _19921_ (.A(_04472_),
    .Y(_04474_));
 sky130_fd_sc_hd__a221o_1 _19922_ (.A1(_04470_),
    .A2(_04472_),
    .B1(_04473_),
    .B2(_04474_),
    .C1(_04440_),
    .X(_04475_));
 sky130_fd_sc_hd__o211ai_1 _19923_ (.A1(_14040_),
    .A2(_01739_),
    .B1(_04469_),
    .C1(_04475_),
    .Y(_01746_));
 sky130_vsdinv _19924_ (.A(net58),
    .Y(_01747_));
 sky130_vsdinv _19925_ (.A(net52),
    .Y(_04476_));
 sky130_vsdinv _19926_ (.A(net35),
    .Y(_01852_));
 sky130_vsdinv _19927_ (.A(net43),
    .Y(_04477_));
 sky130_fd_sc_hd__buf_1 _19928_ (.A(_04418_),
    .X(_04478_));
 sky130_fd_sc_hd__or2_1 _19929_ (.A(_04477_),
    .B(_04478_),
    .X(_04479_));
 sky130_fd_sc_hd__o221a_1 _19930_ (.A1(_04476_),
    .A2(_04426_),
    .B1(_01852_),
    .B2(_04427_),
    .C1(_04479_),
    .X(_01748_));
 sky130_fd_sc_hd__buf_1 _19931_ (.A(_14164_),
    .X(_04480_));
 sky130_fd_sc_hd__buf_1 _19932_ (.A(_14147_),
    .X(_04481_));
 sky130_vsdinv _19933_ (.A(_01750_),
    .Y(_04482_));
 sky130_fd_sc_hd__o22a_1 _19934_ (.A1(_04480_),
    .A2(_01749_),
    .B1(_04481_),
    .B2(_04482_),
    .X(_01751_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _19935_ (.A(_11742_),
    .X(_04483_));
 sky130_fd_sc_hd__buf_1 _19936_ (.A(_04483_),
    .X(_04484_));
 sky130_fd_sc_hd__or2_1 _19937_ (.A(_12144_),
    .B(_04484_),
    .X(_04485_));
 sky130_fd_sc_hd__o221a_1 _19938_ (.A1(_12112_),
    .A2(_04432_),
    .B1(_04433_),
    .B2(_12434_),
    .C1(_04485_),
    .X(_01755_));
 sky130_fd_sc_hd__clkbuf_2 _19939_ (.A(_04447_),
    .X(_04486_));
 sky130_fd_sc_hd__buf_2 _19940_ (.A(_04486_),
    .X(_04487_));
 sky130_fd_sc_hd__clkbuf_2 _19941_ (.A(instr_timer),
    .X(_04488_));
 sky130_fd_sc_hd__buf_1 _19942_ (.A(_04488_),
    .X(_04489_));
 sky130_fd_sc_hd__clkbuf_2 _19943_ (.A(instr_maskirq),
    .X(_04490_));
 sky130_fd_sc_hd__buf_1 _19944_ (.A(_04490_),
    .X(_04491_));
 sky130_fd_sc_hd__a22o_1 _19945_ (.A1(_04489_),
    .A2(\timer[3] ),
    .B1(\irq_mask[3] ),
    .B2(_04491_),
    .X(_04492_));
 sky130_fd_sc_hd__a21oi_2 _19946_ (.A1(_04487_),
    .A2(\cpuregs_rs1[3] ),
    .B1(_04492_),
    .Y(_01757_));
 sky130_fd_sc_hd__o2bb2a_1 _19947_ (.A1_N(_04468_),
    .A2_N(_01753_),
    .B1(_14160_),
    .B2(_01758_),
    .X(_04493_));
 sky130_fd_sc_hd__o22a_2 _19948_ (.A1(_02073_),
    .A2(_13797_),
    .B1(_04473_),
    .B2(_04471_),
    .X(_04494_));
 sky130_vsdinv _19949_ (.A(_04494_),
    .Y(_04495_));
 sky130_fd_sc_hd__nor2_2 _19950_ (.A(\reg_pc[3] ),
    .B(_14268_),
    .Y(_04496_));
 sky130_fd_sc_hd__a21oi_1 _19951_ (.A1(\reg_pc[3] ),
    .A2(_14268_),
    .B1(_04496_),
    .Y(_04497_));
 sky130_vsdinv _19952_ (.A(_04497_),
    .Y(_04498_));
 sky130_fd_sc_hd__a221o_1 _19953_ (.A1(_04495_),
    .A2(_04497_),
    .B1(_04494_),
    .B2(_04498_),
    .C1(_04440_),
    .X(_04499_));
 sky130_fd_sc_hd__o211ai_1 _19954_ (.A1(_04455_),
    .A2(_01752_),
    .B1(_04493_),
    .C1(_04499_),
    .Y(_01759_));
 sky130_vsdinv _19955_ (.A(net59),
    .Y(_01760_));
 sky130_vsdinv _19956_ (.A(net53),
    .Y(_04500_));
 sky130_fd_sc_hd__buf_1 _19957_ (.A(_04421_),
    .X(_04501_));
 sky130_vsdinv _19958_ (.A(net36),
    .Y(_01865_));
 sky130_fd_sc_hd__buf_1 _19959_ (.A(_04416_),
    .X(_04502_));
 sky130_vsdinv _19960_ (.A(net464),
    .Y(_04503_));
 sky130_fd_sc_hd__or2_1 _19961_ (.A(_04503_),
    .B(_04478_),
    .X(_04504_));
 sky130_fd_sc_hd__o221a_1 _19962_ (.A1(_04500_),
    .A2(_04501_),
    .B1(_01865_),
    .B2(_04502_),
    .C1(_04504_),
    .X(_01761_));
 sky130_vsdinv _19963_ (.A(_01763_),
    .Y(_04505_));
 sky130_fd_sc_hd__o22a_1 _19964_ (.A1(_04480_),
    .A2(_01762_),
    .B1(_04481_),
    .B2(_04505_),
    .X(_01764_));
 sky130_fd_sc_hd__buf_1 _19965_ (.A(_13344_),
    .X(_04506_));
 sky130_fd_sc_hd__or2_1 _19966_ (.A(_12143_),
    .B(_04484_),
    .X(_04507_));
 sky130_fd_sc_hd__o221a_1 _19967_ (.A1(_12111_),
    .A2(_04432_),
    .B1(_04506_),
    .B2(_12433_),
    .C1(_04507_),
    .X(_01768_));
 sky130_fd_sc_hd__a22o_1 _19968_ (.A1(_04489_),
    .A2(_14202_),
    .B1(\irq_mask[4] ),
    .B2(_04491_),
    .X(_04508_));
 sky130_fd_sc_hd__a21oi_2 _19969_ (.A1(_04487_),
    .A2(\cpuregs_rs1[4] ),
    .B1(_04508_),
    .Y(_01770_));
 sky130_fd_sc_hd__o22ai_4 _19970_ (.A1(_14265_),
    .A2(_13805_),
    .B1(_04494_),
    .B2(_04496_),
    .Y(_04509_));
 sky130_fd_sc_hd__o22a_1 _19971_ (.A1(_14271_),
    .A2(_13812_),
    .B1(_12081_),
    .B2(\decoded_imm[4] ),
    .X(_04510_));
 sky130_fd_sc_hd__or2_1 _19972_ (.A(_04509_),
    .B(_04510_),
    .X(_04511_));
 sky130_fd_sc_hd__nand2_1 _19973_ (.A(_04509_),
    .B(_04510_),
    .Y(_04512_));
 sky130_fd_sc_hd__buf_1 _19974_ (.A(_04454_),
    .X(_04513_));
 sky130_fd_sc_hd__o2bb2a_1 _19975_ (.A1_N(_04456_),
    .A2_N(_01766_),
    .B1(_04458_),
    .B2(_01771_),
    .X(_04514_));
 sky130_fd_sc_hd__o21ai_1 _19976_ (.A1(_04513_),
    .A2(_01765_),
    .B1(_04514_),
    .Y(_04515_));
 sky130_fd_sc_hd__a31o_1 _19977_ (.A1(_14153_),
    .A2(_04511_),
    .A3(_04512_),
    .B1(_04515_),
    .X(_01772_));
 sky130_vsdinv _19978_ (.A(net60),
    .Y(_01773_));
 sky130_vsdinv _19979_ (.A(net54),
    .Y(_04516_));
 sky130_vsdinv _19980_ (.A(net37),
    .Y(_01878_));
 sky130_vsdinv _19981_ (.A(net46),
    .Y(_04517_));
 sky130_fd_sc_hd__or2_1 _19982_ (.A(_04517_),
    .B(_04478_),
    .X(_04518_));
 sky130_fd_sc_hd__o221a_1 _19983_ (.A1(_04516_),
    .A2(_04501_),
    .B1(_01878_),
    .B2(_04502_),
    .C1(_04518_),
    .X(_01774_));
 sky130_vsdinv _19984_ (.A(_01776_),
    .Y(_04519_));
 sky130_fd_sc_hd__o22a_1 _19985_ (.A1(_04480_),
    .A2(_01775_),
    .B1(_04481_),
    .B2(_04519_),
    .X(_01777_));
 sky130_fd_sc_hd__buf_1 _19986_ (.A(_04431_),
    .X(_04520_));
 sky130_fd_sc_hd__or2_1 _19987_ (.A(_12142_),
    .B(_04484_),
    .X(_04521_));
 sky130_fd_sc_hd__o221a_1 _19988_ (.A1(_12110_),
    .A2(_04520_),
    .B1(_04506_),
    .B2(_12432_),
    .C1(_04521_),
    .X(_01781_));
 sky130_fd_sc_hd__nand2_1 _19989_ (.A(_04449_),
    .B(\cpuregs_rs1[5] ),
    .Y(_04522_));
 sky130_fd_sc_hd__o221a_1 _19990_ (.A1(_04435_),
    .A2(_14204_),
    .B1(_11637_),
    .B2(_04436_),
    .C1(_04522_),
    .X(_01783_));
 sky130_fd_sc_hd__buf_1 _19991_ (.A(_04456_),
    .X(_04523_));
 sky130_fd_sc_hd__nor2_1 _19992_ (.A(\reg_pc[5] ),
    .B(_14280_),
    .Y(_04524_));
 sky130_fd_sc_hd__a21oi_2 _19993_ (.A1(\reg_pc[5] ),
    .A2(_14280_),
    .B1(_04524_),
    .Y(_04525_));
 sky130_fd_sc_hd__o21ai_1 _19994_ (.A1(_14271_),
    .A2(_13812_),
    .B1(_04512_),
    .Y(_04526_));
 sky130_fd_sc_hd__or2_1 _19995_ (.A(_04525_),
    .B(_04526_),
    .X(_04527_));
 sky130_fd_sc_hd__a21oi_1 _19996_ (.A1(_04525_),
    .A2(_04526_),
    .B1(_14159_),
    .Y(_04528_));
 sky130_fd_sc_hd__buf_2 _19997_ (.A(_04458_),
    .X(_04529_));
 sky130_fd_sc_hd__o22ai_2 _19998_ (.A1(_14039_),
    .A2(_01778_),
    .B1(_04529_),
    .B2(_01784_),
    .Y(_04530_));
 sky130_fd_sc_hd__a221o_1 _19999_ (.A1(_04523_),
    .A2(_01779_),
    .B1(_04527_),
    .B2(_04528_),
    .C1(_04530_),
    .X(_01785_));
 sky130_vsdinv _20000_ (.A(net61),
    .Y(_01786_));
 sky130_vsdinv _20001_ (.A(net56),
    .Y(_04531_));
 sky130_vsdinv _20002_ (.A(net38),
    .Y(_01891_));
 sky130_vsdinv _20003_ (.A(net47),
    .Y(_04532_));
 sky130_fd_sc_hd__or2_1 _20004_ (.A(_04532_),
    .B(_04478_),
    .X(_04533_));
 sky130_fd_sc_hd__o221a_1 _20005_ (.A1(_04531_),
    .A2(_04501_),
    .B1(_01891_),
    .B2(_04502_),
    .C1(_04533_),
    .X(_01787_));
 sky130_vsdinv _20006_ (.A(_01789_),
    .Y(_04534_));
 sky130_fd_sc_hd__o22a_1 _20007_ (.A1(_04480_),
    .A2(_01788_),
    .B1(_04481_),
    .B2(_04534_),
    .X(_01790_));
 sky130_fd_sc_hd__or2_1 _20008_ (.A(_12141_),
    .B(_04484_),
    .X(_04535_));
 sky130_fd_sc_hd__o221a_1 _20009_ (.A1(_12109_),
    .A2(_04520_),
    .B1(_04506_),
    .B2(_12431_),
    .C1(_04535_),
    .X(_01794_));
 sky130_fd_sc_hd__a22o_1 _20010_ (.A1(_04489_),
    .A2(\timer[6] ),
    .B1(\irq_mask[6] ),
    .B2(_04491_),
    .X(_04536_));
 sky130_fd_sc_hd__a21oi_2 _20011_ (.A1(_04487_),
    .A2(\cpuregs_rs1[6] ),
    .B1(_04536_),
    .Y(_01796_));
 sky130_fd_sc_hd__o32a_1 _20012_ (.A1(_14271_),
    .A2(_13811_),
    .A3(_04524_),
    .B1(_14276_),
    .B2(_13818_),
    .X(_04537_));
 sky130_vsdinv _20013_ (.A(_04537_),
    .Y(_04538_));
 sky130_fd_sc_hd__a31o_1 _20014_ (.A1(_04510_),
    .A2(_04525_),
    .A3(_04509_),
    .B1(_04538_),
    .X(_04539_));
 sky130_fd_sc_hd__o22a_1 _20015_ (.A1(_04075_),
    .A2(_13824_),
    .B1(_12076_),
    .B2(\decoded_imm[6] ),
    .X(_04540_));
 sky130_fd_sc_hd__or2_1 _20016_ (.A(_04539_),
    .B(_04540_),
    .X(_04541_));
 sky130_fd_sc_hd__nand2_1 _20017_ (.A(_04539_),
    .B(_04540_),
    .Y(_04542_));
 sky130_fd_sc_hd__o2bb2a_1 _20018_ (.A1_N(_04456_),
    .A2_N(_01792_),
    .B1(_04458_),
    .B2(_01797_),
    .X(_04543_));
 sky130_fd_sc_hd__o21ai_1 _20019_ (.A1(_04513_),
    .A2(_01791_),
    .B1(_04543_),
    .Y(_04544_));
 sky130_fd_sc_hd__a31o_1 _20020_ (.A1(_14153_),
    .A2(_04541_),
    .A3(_04542_),
    .B1(_04544_),
    .X(_01798_));
 sky130_vsdinv _20021_ (.A(net62),
    .Y(_01799_));
 sky130_vsdinv _20022_ (.A(net57),
    .Y(_04545_));
 sky130_vsdinv _20023_ (.A(net39),
    .Y(_01904_));
 sky130_vsdinv _20024_ (.A(net48),
    .Y(_04546_));
 sky130_fd_sc_hd__or2_1 _20025_ (.A(_04546_),
    .B(_04418_),
    .X(_04547_));
 sky130_fd_sc_hd__o221a_1 _20026_ (.A1(_04545_),
    .A2(_04501_),
    .B1(_01904_),
    .B2(_04502_),
    .C1(_04547_),
    .X(_01800_));
 sky130_vsdinv _20027_ (.A(_01802_),
    .Y(_04548_));
 sky130_fd_sc_hd__o22a_1 _20028_ (.A1(_14164_),
    .A2(_01801_),
    .B1(_14147_),
    .B2(_04548_),
    .X(_01803_));
 sky130_fd_sc_hd__buf_1 _20029_ (.A(_04483_),
    .X(_04549_));
 sky130_fd_sc_hd__or2_1 _20030_ (.A(_12140_),
    .B(_04549_),
    .X(_04550_));
 sky130_fd_sc_hd__o221a_1 _20031_ (.A1(_12108_),
    .A2(_04520_),
    .B1(_04506_),
    .B2(_12430_),
    .C1(_04550_),
    .X(_01807_));
 sky130_fd_sc_hd__buf_1 _20032_ (.A(_13300_),
    .X(_04551_));
 sky130_fd_sc_hd__buf_1 _20033_ (.A(_13307_),
    .X(_04552_));
 sky130_fd_sc_hd__nand2_1 _20034_ (.A(_04449_),
    .B(\cpuregs_rs1[7] ),
    .Y(_04553_));
 sky130_fd_sc_hd__o221a_1 _20035_ (.A1(_04551_),
    .A2(_14206_),
    .B1(_11638_),
    .B2(_04552_),
    .C1(_04553_),
    .X(_01809_));
 sky130_fd_sc_hd__nor2_1 _20036_ (.A(\reg_pc[7] ),
    .B(_04081_),
    .Y(_04554_));
 sky130_fd_sc_hd__a21oi_2 _20037_ (.A1(\reg_pc[7] ),
    .A2(_04081_),
    .B1(_04554_),
    .Y(_04555_));
 sky130_fd_sc_hd__o21ai_1 _20038_ (.A1(_04075_),
    .A2(_13825_),
    .B1(_04542_),
    .Y(_04556_));
 sky130_fd_sc_hd__or2_1 _20039_ (.A(_04555_),
    .B(_04556_),
    .X(_04557_));
 sky130_fd_sc_hd__a21oi_1 _20040_ (.A1(_04555_),
    .A2(_04556_),
    .B1(_14159_),
    .Y(_04558_));
 sky130_fd_sc_hd__o22ai_4 _20041_ (.A1(_04438_),
    .A2(_01810_),
    .B1(_14039_),
    .B2(_01804_),
    .Y(_04559_));
 sky130_fd_sc_hd__a221o_1 _20042_ (.A1(_04523_),
    .A2(_01805_),
    .B1(_04557_),
    .B2(_04558_),
    .C1(_04559_),
    .X(_01811_));
 sky130_fd_sc_hd__clkbuf_2 _20043_ (.A(\mem_wordsize[2] ),
    .X(_04560_));
 sky130_fd_sc_hd__clkbuf_2 _20044_ (.A(_04560_),
    .X(_04561_));
 sky130_fd_sc_hd__nand2_1 _20045_ (.A(_04561_),
    .B(_01813_),
    .Y(_01814_));
 sky130_fd_sc_hd__nor2_8 _20046_ (.A(latched_is_lb),
    .B(latched_is_lh),
    .Y(_01816_));
 sky130_vsdinv _20047_ (.A(latched_is_lb),
    .Y(_04562_));
 sky130_fd_sc_hd__buf_1 _20048_ (.A(_04562_),
    .X(_04563_));
 sky130_fd_sc_hd__buf_1 _20049_ (.A(_01804_),
    .X(_04564_));
 sky130_vsdinv _20050_ (.A(latched_is_lh),
    .Y(_04565_));
 sky130_fd_sc_hd__buf_1 _20051_ (.A(_04565_),
    .X(_04566_));
 sky130_fd_sc_hd__o22a_1 _20052_ (.A1(_04563_),
    .A2(_04564_),
    .B1(_04566_),
    .B2(_01815_),
    .X(_01817_));
 sky130_fd_sc_hd__buf_1 _20053_ (.A(_13344_),
    .X(_04567_));
 sky130_fd_sc_hd__or2_1 _20054_ (.A(_12139_),
    .B(_04549_),
    .X(_04568_));
 sky130_fd_sc_hd__o221a_1 _20055_ (.A1(_12107_),
    .A2(_04520_),
    .B1(_04567_),
    .B2(_12429_),
    .C1(_04568_),
    .X(_01821_));
 sky130_fd_sc_hd__a22o_1 _20056_ (.A1(_04489_),
    .A2(\timer[8] ),
    .B1(\irq_mask[8] ),
    .B2(_04491_),
    .X(_04569_));
 sky130_fd_sc_hd__a21oi_4 _20057_ (.A1(_04487_),
    .A2(\cpuregs_rs1[8] ),
    .B1(_04569_),
    .Y(_01823_));
 sky130_fd_sc_hd__buf_1 _20058_ (.A(_11726_),
    .X(_04570_));
 sky130_fd_sc_hd__o32a_1 _20059_ (.A1(_04075_),
    .A2(_13824_),
    .A3(_04554_),
    .B1(_04080_),
    .B2(_13828_),
    .X(_04571_));
 sky130_vsdinv _20060_ (.A(_04571_),
    .Y(_04572_));
 sky130_fd_sc_hd__a31o_1 _20061_ (.A1(_04540_),
    .A2(_04555_),
    .A3(_04539_),
    .B1(_04572_),
    .X(_04573_));
 sky130_fd_sc_hd__o22a_1 _20062_ (.A1(_04086_),
    .A2(_13832_),
    .B1(\reg_pc[8] ),
    .B2(\decoded_imm[8] ),
    .X(_04574_));
 sky130_fd_sc_hd__or2_1 _20063_ (.A(_04573_),
    .B(_04574_),
    .X(_04575_));
 sky130_fd_sc_hd__nand2_1 _20064_ (.A(_04573_),
    .B(_04574_),
    .Y(_04576_));
 sky130_fd_sc_hd__clkbuf_2 _20065_ (.A(_12365_),
    .X(_04577_));
 sky130_fd_sc_hd__buf_1 _20066_ (.A(_04577_),
    .X(_04578_));
 sky130_fd_sc_hd__buf_1 _20067_ (.A(_12302_),
    .X(_04579_));
 sky130_fd_sc_hd__o2bb2a_1 _20068_ (.A1_N(_04578_),
    .A2_N(_01819_),
    .B1(_04579_),
    .B2(_01824_),
    .X(_04580_));
 sky130_fd_sc_hd__o21ai_1 _20069_ (.A1(_04513_),
    .A2(_01818_),
    .B1(_04580_),
    .Y(_04581_));
 sky130_fd_sc_hd__a31o_1 _20070_ (.A1(_04570_),
    .A2(_04575_),
    .A3(_04576_),
    .B1(_04581_),
    .X(_01825_));
 sky130_fd_sc_hd__nand2_1 _20071_ (.A(_04561_),
    .B(_01827_),
    .Y(_01828_));
 sky130_fd_sc_hd__o22a_1 _20072_ (.A1(_04563_),
    .A2(_04564_),
    .B1(_04566_),
    .B2(_01829_),
    .X(_01830_));
 sky130_fd_sc_hd__clkbuf_2 _20073_ (.A(_04431_),
    .X(_04582_));
 sky130_fd_sc_hd__or2_1 _20074_ (.A(_12138_),
    .B(_04549_),
    .X(_04583_));
 sky130_fd_sc_hd__o221a_1 _20075_ (.A1(_12106_),
    .A2(_04582_),
    .B1(_04567_),
    .B2(_12428_),
    .C1(_04583_),
    .X(_01834_));
 sky130_fd_sc_hd__buf_1 _20076_ (.A(_04447_),
    .X(_04584_));
 sky130_fd_sc_hd__nand2_1 _20077_ (.A(_04584_),
    .B(\cpuregs_rs1[9] ),
    .Y(_04585_));
 sky130_fd_sc_hd__o221a_1 _20078_ (.A1(_04551_),
    .A2(_14208_),
    .B1(_11656_),
    .B2(_04552_),
    .C1(_04585_),
    .X(_01836_));
 sky130_fd_sc_hd__nor2_1 _20079_ (.A(\reg_pc[9] ),
    .B(_04098_),
    .Y(_04586_));
 sky130_fd_sc_hd__a21oi_2 _20080_ (.A1(\reg_pc[9] ),
    .A2(_04098_),
    .B1(_04586_),
    .Y(_04587_));
 sky130_fd_sc_hd__o21ai_1 _20081_ (.A1(_04086_),
    .A2(_13833_),
    .B1(_04576_),
    .Y(_04588_));
 sky130_fd_sc_hd__or2_1 _20082_ (.A(_04587_),
    .B(_04588_),
    .X(_04589_));
 sky130_fd_sc_hd__a21oi_1 _20083_ (.A1(_04587_),
    .A2(_04588_),
    .B1(_14159_),
    .Y(_04590_));
 sky130_fd_sc_hd__clkbuf_4 _20084_ (.A(_04454_),
    .X(_04591_));
 sky130_fd_sc_hd__o22ai_4 _20085_ (.A1(_04591_),
    .A2(_01831_),
    .B1(_04529_),
    .B2(_01837_),
    .Y(_04592_));
 sky130_fd_sc_hd__a221o_1 _20086_ (.A1(_04523_),
    .A2(_01832_),
    .B1(_04589_),
    .B2(_04590_),
    .C1(_04592_),
    .X(_01838_));
 sky130_fd_sc_hd__nand2_1 _20087_ (.A(_04561_),
    .B(_01840_),
    .Y(_01841_));
 sky130_fd_sc_hd__o22a_1 _20088_ (.A1(_04563_),
    .A2(_04564_),
    .B1(_04566_),
    .B2(_01842_),
    .X(_01843_));
 sky130_fd_sc_hd__or2_1 _20089_ (.A(_12137_),
    .B(_04549_),
    .X(_04593_));
 sky130_fd_sc_hd__o221a_1 _20090_ (.A1(_12105_),
    .A2(_04582_),
    .B1(_04567_),
    .B2(_12427_),
    .C1(_04593_),
    .X(_01847_));
 sky130_fd_sc_hd__clkbuf_4 _20091_ (.A(_04448_),
    .X(_04594_));
 sky130_fd_sc_hd__buf_1 _20092_ (.A(_04488_),
    .X(_04595_));
 sky130_fd_sc_hd__buf_1 _20093_ (.A(_04490_),
    .X(_04596_));
 sky130_fd_sc_hd__a22o_1 _20094_ (.A1(_04595_),
    .A2(\timer[10] ),
    .B1(\irq_mask[10] ),
    .B2(_04596_),
    .X(_04597_));
 sky130_fd_sc_hd__a21oi_4 _20095_ (.A1(_04594_),
    .A2(\cpuregs_rs1[10] ),
    .B1(_04597_),
    .Y(_01849_));
 sky130_fd_sc_hd__o22a_1 _20096_ (.A1(_04102_),
    .A2(_13843_),
    .B1(\reg_pc[10] ),
    .B2(\decoded_imm[10] ),
    .X(_04598_));
 sky130_fd_sc_hd__o32a_1 _20097_ (.A1(_04086_),
    .A2(_13831_),
    .A3(_04586_),
    .B1(_04095_),
    .B2(_13839_),
    .X(_04599_));
 sky130_vsdinv _20098_ (.A(_04599_),
    .Y(_04600_));
 sky130_fd_sc_hd__a31o_1 _20099_ (.A1(_04574_),
    .A2(_04587_),
    .A3(_04573_),
    .B1(_04600_),
    .X(_04601_));
 sky130_fd_sc_hd__or2_1 _20100_ (.A(_04598_),
    .B(_04601_),
    .X(_04602_));
 sky130_fd_sc_hd__nand2_1 _20101_ (.A(_04598_),
    .B(_04601_),
    .Y(_04603_));
 sky130_fd_sc_hd__o2bb2a_1 _20102_ (.A1_N(_04578_),
    .A2_N(_01845_),
    .B1(_04579_),
    .B2(_01850_),
    .X(_04604_));
 sky130_fd_sc_hd__o21ai_2 _20103_ (.A1(_04513_),
    .A2(_01844_),
    .B1(_04604_),
    .Y(_04605_));
 sky130_fd_sc_hd__a31o_1 _20104_ (.A1(_04570_),
    .A2(_04602_),
    .A3(_04603_),
    .B1(_04605_),
    .X(_01851_));
 sky130_fd_sc_hd__nand2_1 _20105_ (.A(_04561_),
    .B(_01853_),
    .Y(_01854_));
 sky130_fd_sc_hd__o22a_1 _20106_ (.A1(_04563_),
    .A2(_04564_),
    .B1(_04566_),
    .B2(_01855_),
    .X(_01856_));
 sky130_fd_sc_hd__buf_1 _20107_ (.A(_04483_),
    .X(_04606_));
 sky130_fd_sc_hd__or2_1 _20108_ (.A(_12136_),
    .B(_04606_),
    .X(_04607_));
 sky130_fd_sc_hd__o221a_1 _20109_ (.A1(_12104_),
    .A2(_04582_),
    .B1(_04567_),
    .B2(_12426_),
    .C1(_04607_),
    .X(_01860_));
 sky130_fd_sc_hd__nand2_1 _20110_ (.A(_04584_),
    .B(\cpuregs_rs1[11] ),
    .Y(_04608_));
 sky130_fd_sc_hd__o221a_2 _20111_ (.A1(_04551_),
    .A2(_14210_),
    .B1(_11657_),
    .B2(_04552_),
    .C1(_04608_),
    .X(_01862_));
 sky130_fd_sc_hd__o22a_1 _20112_ (.A1(_04109_),
    .A2(_13848_),
    .B1(\reg_pc[11] ),
    .B2(\decoded_imm[11] ),
    .X(_04609_));
 sky130_fd_sc_hd__o21ai_1 _20113_ (.A1(_04102_),
    .A2(_13843_),
    .B1(_04603_),
    .Y(_04610_));
 sky130_fd_sc_hd__nand2_1 _20114_ (.A(_04609_),
    .B(_04610_),
    .Y(_04611_));
 sky130_fd_sc_hd__or2_1 _20115_ (.A(_04609_),
    .B(_04610_),
    .X(_04612_));
 sky130_fd_sc_hd__clkbuf_2 _20116_ (.A(_04454_),
    .X(_04613_));
 sky130_fd_sc_hd__o2bb2a_1 _20117_ (.A1_N(_04578_),
    .A2_N(_01858_),
    .B1(_04579_),
    .B2(_01863_),
    .X(_04614_));
 sky130_fd_sc_hd__o21ai_2 _20118_ (.A1(_04613_),
    .A2(_01857_),
    .B1(_04614_),
    .Y(_04615_));
 sky130_fd_sc_hd__a31o_1 _20119_ (.A1(_04570_),
    .A2(_04611_),
    .A3(_04612_),
    .B1(_04615_),
    .X(_01864_));
 sky130_fd_sc_hd__buf_1 _20120_ (.A(_04560_),
    .X(_04616_));
 sky130_fd_sc_hd__nand2_1 _20121_ (.A(_04616_),
    .B(_01866_),
    .Y(_01867_));
 sky130_fd_sc_hd__buf_1 _20122_ (.A(_04562_),
    .X(_04617_));
 sky130_fd_sc_hd__buf_1 _20123_ (.A(_01804_),
    .X(_04618_));
 sky130_fd_sc_hd__clkbuf_2 _20124_ (.A(_04565_),
    .X(_04619_));
 sky130_fd_sc_hd__o22a_1 _20125_ (.A1(_04617_),
    .A2(_04618_),
    .B1(_04619_),
    .B2(_01868_),
    .X(_01869_));
 sky130_fd_sc_hd__clkbuf_2 _20126_ (.A(_11743_),
    .X(_04620_));
 sky130_fd_sc_hd__clkbuf_2 _20127_ (.A(_04620_),
    .X(_04621_));
 sky130_fd_sc_hd__or2_1 _20128_ (.A(_12135_),
    .B(_04606_),
    .X(_04622_));
 sky130_fd_sc_hd__o221a_1 _20129_ (.A1(_12103_),
    .A2(_04582_),
    .B1(_04621_),
    .B2(_12425_),
    .C1(_04622_),
    .X(_01873_));
 sky130_fd_sc_hd__a22o_1 _20130_ (.A1(_04595_),
    .A2(\timer[12] ),
    .B1(\irq_mask[12] ),
    .B2(_04596_),
    .X(_04623_));
 sky130_fd_sc_hd__a21oi_4 _20131_ (.A1(_04594_),
    .A2(\cpuregs_rs1[12] ),
    .B1(_04623_),
    .Y(_01875_));
 sky130_fd_sc_hd__o22a_1 _20132_ (.A1(_04114_),
    .A2(_13854_),
    .B1(\reg_pc[12] ),
    .B2(\decoded_imm[12] ),
    .X(_04624_));
 sky130_fd_sc_hd__o21ai_1 _20133_ (.A1(_04109_),
    .A2(_13848_),
    .B1(_04611_),
    .Y(_04625_));
 sky130_fd_sc_hd__or2_1 _20134_ (.A(_04624_),
    .B(_04625_),
    .X(_04626_));
 sky130_fd_sc_hd__nand2_1 _20135_ (.A(_04624_),
    .B(_04625_),
    .Y(_04627_));
 sky130_fd_sc_hd__o2bb2a_1 _20136_ (.A1_N(_04578_),
    .A2_N(_01871_),
    .B1(_04579_),
    .B2(_01876_),
    .X(_04628_));
 sky130_fd_sc_hd__o21ai_2 _20137_ (.A1(_04613_),
    .A2(_01870_),
    .B1(_04628_),
    .Y(_04629_));
 sky130_fd_sc_hd__a31o_1 _20138_ (.A1(_04570_),
    .A2(_04626_),
    .A3(_04627_),
    .B1(_04629_),
    .X(_01877_));
 sky130_fd_sc_hd__nand2_1 _20139_ (.A(_04616_),
    .B(_01879_),
    .Y(_01880_));
 sky130_fd_sc_hd__o22a_1 _20140_ (.A1(_04617_),
    .A2(_04618_),
    .B1(_04619_),
    .B2(_01881_),
    .X(_01882_));
 sky130_fd_sc_hd__buf_2 _20141_ (.A(_11741_),
    .X(_04630_));
 sky130_fd_sc_hd__buf_1 _20142_ (.A(_04630_),
    .X(_04631_));
 sky130_fd_sc_hd__or2_1 _20143_ (.A(_12134_),
    .B(_04606_),
    .X(_04632_));
 sky130_fd_sc_hd__o221a_1 _20144_ (.A1(_12102_),
    .A2(_04631_),
    .B1(_04621_),
    .B2(_12424_),
    .C1(_04632_),
    .X(_01886_));
 sky130_fd_sc_hd__nand2_1 _20145_ (.A(_04584_),
    .B(\cpuregs_rs1[13] ),
    .Y(_04633_));
 sky130_fd_sc_hd__o221a_2 _20146_ (.A1(_04551_),
    .A2(_14212_),
    .B1(_11644_),
    .B2(_04552_),
    .C1(_04633_),
    .X(_01888_));
 sky130_fd_sc_hd__buf_1 _20147_ (.A(_14152_),
    .X(_04634_));
 sky130_fd_sc_hd__o22a_1 _20148_ (.A1(_04120_),
    .A2(_13863_),
    .B1(\reg_pc[13] ),
    .B2(\decoded_imm[13] ),
    .X(_04635_));
 sky130_fd_sc_hd__o21ai_1 _20149_ (.A1(_04114_),
    .A2(_13854_),
    .B1(_04627_),
    .Y(_04636_));
 sky130_fd_sc_hd__nand2_1 _20150_ (.A(_04635_),
    .B(_04636_),
    .Y(_04637_));
 sky130_fd_sc_hd__or2_1 _20151_ (.A(_04635_),
    .B(_04636_),
    .X(_04638_));
 sky130_fd_sc_hd__buf_1 _20152_ (.A(_04577_),
    .X(_04639_));
 sky130_fd_sc_hd__buf_1 _20153_ (.A(_04457_),
    .X(_04640_));
 sky130_fd_sc_hd__o2bb2a_1 _20154_ (.A1_N(_04639_),
    .A2_N(_01884_),
    .B1(_04640_),
    .B2(_01889_),
    .X(_04641_));
 sky130_fd_sc_hd__o21ai_2 _20155_ (.A1(_04613_),
    .A2(_01883_),
    .B1(_04641_),
    .Y(_04642_));
 sky130_fd_sc_hd__a31o_1 _20156_ (.A1(_04634_),
    .A2(_04637_),
    .A3(_04638_),
    .B1(_04642_),
    .X(_01890_));
 sky130_fd_sc_hd__nand2_1 _20157_ (.A(_04616_),
    .B(_01892_),
    .Y(_01893_));
 sky130_fd_sc_hd__o22a_1 _20158_ (.A1(_04617_),
    .A2(_04618_),
    .B1(_04619_),
    .B2(_01894_),
    .X(_01895_));
 sky130_fd_sc_hd__or2_1 _20159_ (.A(_12133_),
    .B(_04606_),
    .X(_04643_));
 sky130_fd_sc_hd__o221a_1 _20160_ (.A1(_12101_),
    .A2(_04631_),
    .B1(_04621_),
    .B2(_12423_),
    .C1(_04643_),
    .X(_01899_));
 sky130_fd_sc_hd__a22o_1 _20161_ (.A1(_04595_),
    .A2(\timer[14] ),
    .B1(\irq_mask[14] ),
    .B2(_04596_),
    .X(_04644_));
 sky130_fd_sc_hd__a21oi_4 _20162_ (.A1(_04594_),
    .A2(\cpuregs_rs1[14] ),
    .B1(_04644_),
    .Y(_01901_));
 sky130_fd_sc_hd__o22a_1 _20163_ (.A1(_04127_),
    .A2(_13868_),
    .B1(\reg_pc[14] ),
    .B2(\decoded_imm[14] ),
    .X(_04645_));
 sky130_fd_sc_hd__o21ai_1 _20164_ (.A1(_04120_),
    .A2(_13863_),
    .B1(_04637_),
    .Y(_04646_));
 sky130_fd_sc_hd__or2_1 _20165_ (.A(_04645_),
    .B(_04646_),
    .X(_04647_));
 sky130_fd_sc_hd__nand2_1 _20166_ (.A(_04645_),
    .B(_04646_),
    .Y(_04648_));
 sky130_fd_sc_hd__o2bb2a_1 _20167_ (.A1_N(_04639_),
    .A2_N(_01897_),
    .B1(_04640_),
    .B2(_01902_),
    .X(_04649_));
 sky130_fd_sc_hd__o21ai_2 _20168_ (.A1(_04613_),
    .A2(_01896_),
    .B1(_04649_),
    .Y(_04650_));
 sky130_fd_sc_hd__a31o_1 _20169_ (.A1(_04634_),
    .A2(_04647_),
    .A3(_04648_),
    .B1(_04650_),
    .X(_01903_));
 sky130_fd_sc_hd__nand2_1 _20170_ (.A(_04616_),
    .B(_01905_),
    .Y(_01906_));
 sky130_fd_sc_hd__o22a_4 _20171_ (.A1(_04617_),
    .A2(_04618_),
    .B1(_04619_),
    .B2(_01907_),
    .X(_01908_));
 sky130_fd_sc_hd__buf_2 _20172_ (.A(_11742_),
    .X(_04651_));
 sky130_fd_sc_hd__buf_1 _20173_ (.A(_04651_),
    .X(_04652_));
 sky130_fd_sc_hd__or2_1 _20174_ (.A(_12132_),
    .B(_04652_),
    .X(_04653_));
 sky130_fd_sc_hd__o221a_1 _20175_ (.A1(_12100_),
    .A2(_04631_),
    .B1(_04621_),
    .B2(_12422_),
    .C1(_04653_),
    .X(_01912_));
 sky130_fd_sc_hd__clkbuf_2 _20176_ (.A(_13300_),
    .X(_04654_));
 sky130_fd_sc_hd__clkbuf_2 _20177_ (.A(_13307_),
    .X(_04655_));
 sky130_fd_sc_hd__nand2_1 _20178_ (.A(_04584_),
    .B(\cpuregs_rs1[15] ),
    .Y(_04656_));
 sky130_fd_sc_hd__o221a_2 _20179_ (.A1(_04654_),
    .A2(_14214_),
    .B1(_11645_),
    .B2(_04655_),
    .C1(_04656_),
    .X(_01914_));
 sky130_fd_sc_hd__o22a_1 _20180_ (.A1(_04133_),
    .A2(_13873_),
    .B1(\reg_pc[15] ),
    .B2(\decoded_imm[15] ),
    .X(_04657_));
 sky130_fd_sc_hd__o21ai_1 _20181_ (.A1(_04127_),
    .A2(_13868_),
    .B1(_04648_),
    .Y(_04658_));
 sky130_fd_sc_hd__nand2_1 _20182_ (.A(_04657_),
    .B(_04658_),
    .Y(_04659_));
 sky130_fd_sc_hd__or2_1 _20183_ (.A(_04657_),
    .B(_04658_),
    .X(_04660_));
 sky130_fd_sc_hd__buf_4 _20184_ (.A(_14038_),
    .X(_04661_));
 sky130_fd_sc_hd__o2bb2a_1 _20185_ (.A1_N(_04639_),
    .A2_N(_01910_),
    .B1(_04640_),
    .B2(_01915_),
    .X(_04662_));
 sky130_fd_sc_hd__o21ai_4 _20186_ (.A1(_04661_),
    .A2(_01909_),
    .B1(_04662_),
    .Y(_04663_));
 sky130_fd_sc_hd__a31o_1 _20187_ (.A1(_04634_),
    .A2(_04659_),
    .A3(_04660_),
    .B1(_04663_),
    .X(_01916_));
 sky130_fd_sc_hd__buf_1 _20188_ (.A(_04415_),
    .X(_04664_));
 sky130_fd_sc_hd__buf_1 _20189_ (.A(_04664_),
    .X(_04665_));
 sky130_fd_sc_hd__or2_1 _20190_ (.A(_04428_),
    .B(_04665_),
    .X(_01917_));
 sky130_fd_sc_hd__buf_1 _20191_ (.A(_04620_),
    .X(_04666_));
 sky130_fd_sc_hd__or2_1 _20192_ (.A(_12131_),
    .B(_04652_),
    .X(_04667_));
 sky130_fd_sc_hd__o221a_1 _20193_ (.A1(_12099_),
    .A2(_04631_),
    .B1(_04666_),
    .B2(_12421_),
    .C1(_04667_),
    .X(_01921_));
 sky130_fd_sc_hd__a22o_1 _20194_ (.A1(_04595_),
    .A2(\timer[16] ),
    .B1(\irq_mask[16] ),
    .B2(_04596_),
    .X(_04668_));
 sky130_fd_sc_hd__a21oi_4 _20195_ (.A1(_04594_),
    .A2(\cpuregs_rs1[16] ),
    .B1(_04668_),
    .Y(_01923_));
 sky130_fd_sc_hd__o21ai_1 _20196_ (.A1(_04133_),
    .A2(_13873_),
    .B1(_04659_),
    .Y(_04669_));
 sky130_fd_sc_hd__o22a_1 _20197_ (.A1(_04139_),
    .A2(_13880_),
    .B1(\reg_pc[16] ),
    .B2(\decoded_imm[16] ),
    .X(_04670_));
 sky130_fd_sc_hd__or2_1 _20198_ (.A(_04669_),
    .B(_04670_),
    .X(_04671_));
 sky130_fd_sc_hd__nand2_1 _20199_ (.A(_04669_),
    .B(_04670_),
    .Y(_04672_));
 sky130_fd_sc_hd__o2bb2a_1 _20200_ (.A1_N(_04639_),
    .A2_N(_01919_),
    .B1(_04640_),
    .B2(_01924_),
    .X(_04673_));
 sky130_fd_sc_hd__o21ai_4 _20201_ (.A1(_04661_),
    .A2(_01918_),
    .B1(_04673_),
    .Y(_04674_));
 sky130_fd_sc_hd__a31o_1 _20202_ (.A1(_04634_),
    .A2(_04671_),
    .A3(_04672_),
    .B1(_04674_),
    .X(_01925_));
 sky130_fd_sc_hd__or2_1 _20203_ (.A(_04443_),
    .B(_04665_),
    .X(_01926_));
 sky130_fd_sc_hd__buf_1 _20204_ (.A(_04630_),
    .X(_04675_));
 sky130_fd_sc_hd__or2_1 _20205_ (.A(_12130_),
    .B(_04652_),
    .X(_04676_));
 sky130_fd_sc_hd__o221a_1 _20206_ (.A1(_12098_),
    .A2(_04675_),
    .B1(_04666_),
    .B2(_12420_),
    .C1(_04676_),
    .X(_01930_));
 sky130_fd_sc_hd__clkbuf_4 _20207_ (.A(_04448_),
    .X(_04677_));
 sky130_fd_sc_hd__buf_1 _20208_ (.A(_04488_),
    .X(_04678_));
 sky130_fd_sc_hd__buf_1 _20209_ (.A(_04490_),
    .X(_04679_));
 sky130_fd_sc_hd__a22o_1 _20210_ (.A1(_04678_),
    .A2(\timer[17] ),
    .B1(\irq_mask[17] ),
    .B2(_04679_),
    .X(_04680_));
 sky130_fd_sc_hd__a21oi_4 _20211_ (.A1(_04677_),
    .A2(\cpuregs_rs1[17] ),
    .B1(_04680_),
    .Y(_01932_));
 sky130_fd_sc_hd__nor2_2 _20212_ (.A(\reg_pc[17] ),
    .B(_04148_),
    .Y(_04681_));
 sky130_fd_sc_hd__a21oi_4 _20213_ (.A1(\reg_pc[17] ),
    .A2(_04148_),
    .B1(_04681_),
    .Y(_04682_));
 sky130_fd_sc_hd__o21ai_2 _20214_ (.A1(_04139_),
    .A2(_13881_),
    .B1(_04672_),
    .Y(_04683_));
 sky130_fd_sc_hd__or2_1 _20215_ (.A(_04682_),
    .B(_04683_),
    .X(_04684_));
 sky130_fd_sc_hd__a21oi_1 _20216_ (.A1(_04682_),
    .A2(_04683_),
    .B1(_14061_),
    .Y(_04685_));
 sky130_fd_sc_hd__o22ai_2 _20217_ (.A1(_04591_),
    .A2(_01927_),
    .B1(_04529_),
    .B2(_01933_),
    .Y(_04686_));
 sky130_fd_sc_hd__a221o_2 _20218_ (.A1(_04523_),
    .A2(_01928_),
    .B1(_04684_),
    .B2(_04685_),
    .C1(_04686_),
    .X(_01934_));
 sky130_fd_sc_hd__or2_1 _20219_ (.A(_04462_),
    .B(_04665_),
    .X(_01935_));
 sky130_fd_sc_hd__or2_1 _20220_ (.A(_12129_),
    .B(_04652_),
    .X(_04687_));
 sky130_fd_sc_hd__o221a_1 _20221_ (.A1(_12097_),
    .A2(_04675_),
    .B1(_04666_),
    .B2(_12419_),
    .C1(_04687_),
    .X(_01939_));
 sky130_fd_sc_hd__buf_1 _20222_ (.A(_04447_),
    .X(_04688_));
 sky130_fd_sc_hd__nand2_1 _20223_ (.A(_04688_),
    .B(\cpuregs_rs1[18] ),
    .Y(_04689_));
 sky130_fd_sc_hd__o221a_2 _20224_ (.A1(_04654_),
    .A2(_14170_),
    .B1(_12312_),
    .B2(_04655_),
    .C1(_04689_),
    .X(_01941_));
 sky130_fd_sc_hd__buf_1 _20225_ (.A(_14152_),
    .X(_04690_));
 sky130_fd_sc_hd__o22a_1 _20226_ (.A1(_04153_),
    .A2(_13892_),
    .B1(\reg_pc[18] ),
    .B2(\decoded_imm[18] ),
    .X(_04691_));
 sky130_fd_sc_hd__o32a_1 _20227_ (.A1(_04139_),
    .A2(_13879_),
    .A3(_04681_),
    .B1(_04146_),
    .B2(_13887_),
    .X(_04692_));
 sky130_vsdinv _20228_ (.A(_04692_),
    .Y(_04693_));
 sky130_fd_sc_hd__a31o_1 _20229_ (.A1(_04670_),
    .A2(_04682_),
    .A3(_04669_),
    .B1(_04693_),
    .X(_04694_));
 sky130_fd_sc_hd__or2_1 _20230_ (.A(_04691_),
    .B(_04694_),
    .X(_04695_));
 sky130_fd_sc_hd__nand2_1 _20231_ (.A(_04691_),
    .B(_04694_),
    .Y(_04696_));
 sky130_fd_sc_hd__clkbuf_1 _20232_ (.A(_04577_),
    .X(_04697_));
 sky130_fd_sc_hd__buf_1 _20233_ (.A(_04457_),
    .X(_04698_));
 sky130_fd_sc_hd__o2bb2a_1 _20234_ (.A1_N(_04697_),
    .A2_N(_01937_),
    .B1(_04698_),
    .B2(_01942_),
    .X(_04699_));
 sky130_fd_sc_hd__o21ai_4 _20235_ (.A1(_04661_),
    .A2(_01936_),
    .B1(_04699_),
    .Y(_04700_));
 sky130_fd_sc_hd__a31o_1 _20236_ (.A1(_04690_),
    .A2(_04695_),
    .A3(_04696_),
    .B1(_04700_),
    .X(_01943_));
 sky130_fd_sc_hd__or2_1 _20237_ (.A(_04477_),
    .B(_04665_),
    .X(_01944_));
 sky130_fd_sc_hd__buf_1 _20238_ (.A(_04651_),
    .X(_04701_));
 sky130_fd_sc_hd__or2_1 _20239_ (.A(_12128_),
    .B(_04701_),
    .X(_04702_));
 sky130_fd_sc_hd__o221a_1 _20240_ (.A1(_12096_),
    .A2(_04675_),
    .B1(_04666_),
    .B2(_12418_),
    .C1(_04702_),
    .X(_01948_));
 sky130_fd_sc_hd__a22o_1 _20241_ (.A1(_04678_),
    .A2(\timer[19] ),
    .B1(\irq_mask[19] ),
    .B2(_04679_),
    .X(_04703_));
 sky130_fd_sc_hd__a21oi_4 _20242_ (.A1(_04677_),
    .A2(\cpuregs_rs1[19] ),
    .B1(_04703_),
    .Y(_01950_));
 sky130_fd_sc_hd__o22a_1 _20243_ (.A1(_04161_),
    .A2(_13897_),
    .B1(\reg_pc[19] ),
    .B2(\decoded_imm[19] ),
    .X(_04704_));
 sky130_fd_sc_hd__o21ai_1 _20244_ (.A1(_04153_),
    .A2(_13892_),
    .B1(_04696_),
    .Y(_04705_));
 sky130_fd_sc_hd__nand2_1 _20245_ (.A(_04704_),
    .B(_04705_),
    .Y(_04706_));
 sky130_fd_sc_hd__or2_1 _20246_ (.A(_04704_),
    .B(_04705_),
    .X(_04707_));
 sky130_fd_sc_hd__o2bb2a_1 _20247_ (.A1_N(_04697_),
    .A2_N(_01946_),
    .B1(_04698_),
    .B2(_01951_),
    .X(_04708_));
 sky130_fd_sc_hd__o21ai_4 _20248_ (.A1(_04661_),
    .A2(_01945_),
    .B1(_04708_),
    .Y(_04709_));
 sky130_fd_sc_hd__a31o_1 _20249_ (.A1(_04690_),
    .A2(_04706_),
    .A3(_04707_),
    .B1(_04709_),
    .X(_01952_));
 sky130_fd_sc_hd__buf_1 _20250_ (.A(_04664_),
    .X(_04710_));
 sky130_fd_sc_hd__or2_1 _20251_ (.A(_04503_),
    .B(_04710_),
    .X(_01953_));
 sky130_fd_sc_hd__buf_1 _20252_ (.A(_04620_),
    .X(_04711_));
 sky130_fd_sc_hd__or2_1 _20253_ (.A(_12127_),
    .B(_04701_),
    .X(_04712_));
 sky130_fd_sc_hd__o221a_1 _20254_ (.A1(_12095_),
    .A2(_04675_),
    .B1(_04711_),
    .B2(_12417_),
    .C1(_04712_),
    .X(_01957_));
 sky130_fd_sc_hd__nand2_1 _20255_ (.A(_04688_),
    .B(\cpuregs_rs1[20] ),
    .Y(_04713_));
 sky130_fd_sc_hd__o221a_2 _20256_ (.A1(_04654_),
    .A2(_14216_),
    .B1(_11662_),
    .B2(_04655_),
    .C1(_04713_),
    .X(_01959_));
 sky130_fd_sc_hd__o22a_1 _20257_ (.A1(_04166_),
    .A2(_14230_),
    .B1(\reg_pc[20] ),
    .B2(\decoded_imm[20] ),
    .X(_04714_));
 sky130_fd_sc_hd__o21ai_1 _20258_ (.A1(_04161_),
    .A2(_13897_),
    .B1(_04706_),
    .Y(_04715_));
 sky130_fd_sc_hd__or2_1 _20259_ (.A(_04714_),
    .B(_04715_),
    .X(_04716_));
 sky130_fd_sc_hd__nand2_1 _20260_ (.A(_04714_),
    .B(_04715_),
    .Y(_04717_));
 sky130_fd_sc_hd__buf_4 _20261_ (.A(_14038_),
    .X(_04718_));
 sky130_fd_sc_hd__o2bb2a_1 _20262_ (.A1_N(_04697_),
    .A2_N(_01955_),
    .B1(_04698_),
    .B2(_01960_),
    .X(_04719_));
 sky130_fd_sc_hd__o21ai_4 _20263_ (.A1(_04718_),
    .A2(_01954_),
    .B1(_04719_),
    .Y(_04720_));
 sky130_fd_sc_hd__a31o_1 _20264_ (.A1(_04690_),
    .A2(_04716_),
    .A3(_04717_),
    .B1(_04720_),
    .X(_01961_));
 sky130_fd_sc_hd__or2_1 _20265_ (.A(_04517_),
    .B(_04710_),
    .X(_01962_));
 sky130_fd_sc_hd__buf_1 _20266_ (.A(_04630_),
    .X(_04721_));
 sky130_fd_sc_hd__or2_1 _20267_ (.A(_12126_),
    .B(_04701_),
    .X(_04722_));
 sky130_fd_sc_hd__o221a_1 _20268_ (.A1(_12094_),
    .A2(_04721_),
    .B1(_04711_),
    .B2(_12416_),
    .C1(_04722_),
    .X(_01966_));
 sky130_fd_sc_hd__a22o_1 _20269_ (.A1(_04678_),
    .A2(\timer[21] ),
    .B1(\irq_mask[21] ),
    .B2(_04679_),
    .X(_04723_));
 sky130_fd_sc_hd__a21oi_4 _20270_ (.A1(_04677_),
    .A2(\cpuregs_rs1[21] ),
    .B1(_04723_),
    .Y(_01968_));
 sky130_fd_sc_hd__o22a_1 _20271_ (.A1(_04172_),
    .A2(_14232_),
    .B1(\reg_pc[21] ),
    .B2(\decoded_imm[21] ),
    .X(_04724_));
 sky130_fd_sc_hd__o21ai_1 _20272_ (.A1(_04166_),
    .A2(_14231_),
    .B1(_04717_),
    .Y(_04725_));
 sky130_fd_sc_hd__nand2_1 _20273_ (.A(_04724_),
    .B(_04725_),
    .Y(_04726_));
 sky130_fd_sc_hd__or2_1 _20274_ (.A(_04724_),
    .B(_04725_),
    .X(_04727_));
 sky130_fd_sc_hd__o2bb2a_1 _20275_ (.A1_N(_04697_),
    .A2_N(_01964_),
    .B1(_04698_),
    .B2(_01969_),
    .X(_04728_));
 sky130_fd_sc_hd__o21ai_4 _20276_ (.A1(_04718_),
    .A2(_01963_),
    .B1(_04728_),
    .Y(_04729_));
 sky130_fd_sc_hd__a31o_1 _20277_ (.A1(_04690_),
    .A2(_04726_),
    .A3(_04727_),
    .B1(_04729_),
    .X(_01970_));
 sky130_fd_sc_hd__or2_1 _20278_ (.A(_04532_),
    .B(_04710_),
    .X(_01971_));
 sky130_fd_sc_hd__or2_1 _20279_ (.A(_12125_),
    .B(_04701_),
    .X(_04730_));
 sky130_fd_sc_hd__o221a_1 _20280_ (.A1(_12093_),
    .A2(_04721_),
    .B1(_04711_),
    .B2(_12415_),
    .C1(_04730_),
    .X(_01975_));
 sky130_fd_sc_hd__nand2_1 _20281_ (.A(_04688_),
    .B(\cpuregs_rs1[22] ),
    .Y(_04731_));
 sky130_fd_sc_hd__o221a_2 _20282_ (.A1(_04654_),
    .A2(_14218_),
    .B1(_11663_),
    .B2(_04655_),
    .C1(_04731_),
    .X(_01977_));
 sky130_fd_sc_hd__clkbuf_2 _20283_ (.A(_14152_),
    .X(_04732_));
 sky130_fd_sc_hd__o22a_1 _20284_ (.A1(_04178_),
    .A2(_14234_),
    .B1(\reg_pc[22] ),
    .B2(\decoded_imm[22] ),
    .X(_04733_));
 sky130_fd_sc_hd__o21ai_1 _20285_ (.A1(_04172_),
    .A2(_14233_),
    .B1(_04726_),
    .Y(_04734_));
 sky130_fd_sc_hd__or2_1 _20286_ (.A(_04733_),
    .B(_04734_),
    .X(_04735_));
 sky130_fd_sc_hd__nand2_1 _20287_ (.A(_04733_),
    .B(_04734_),
    .Y(_04736_));
 sky130_fd_sc_hd__buf_1 _20288_ (.A(_04577_),
    .X(_04737_));
 sky130_fd_sc_hd__buf_1 _20289_ (.A(_04457_),
    .X(_04738_));
 sky130_fd_sc_hd__o2bb2a_1 _20290_ (.A1_N(_04737_),
    .A2_N(_01973_),
    .B1(_04738_),
    .B2(_01978_),
    .X(_04739_));
 sky130_fd_sc_hd__o21ai_4 _20291_ (.A1(_04718_),
    .A2(_01972_),
    .B1(_04739_),
    .Y(_04740_));
 sky130_fd_sc_hd__a31o_1 _20292_ (.A1(_04732_),
    .A2(_04735_),
    .A3(_04736_),
    .B1(_04740_),
    .X(_01979_));
 sky130_fd_sc_hd__or2_1 _20293_ (.A(_04546_),
    .B(_04710_),
    .X(_01980_));
 sky130_fd_sc_hd__buf_1 _20294_ (.A(_04651_),
    .X(_04741_));
 sky130_fd_sc_hd__or2_1 _20295_ (.A(_12124_),
    .B(_04741_),
    .X(_04742_));
 sky130_fd_sc_hd__o221a_1 _20296_ (.A1(_12092_),
    .A2(_04721_),
    .B1(_04711_),
    .B2(_12414_),
    .C1(_04742_),
    .X(_01984_));
 sky130_fd_sc_hd__a22o_1 _20297_ (.A1(_04678_),
    .A2(\timer[23] ),
    .B1(\irq_mask[23] ),
    .B2(_04679_),
    .X(_04743_));
 sky130_fd_sc_hd__a21oi_4 _20298_ (.A1(_04677_),
    .A2(\cpuregs_rs1[23] ),
    .B1(_04743_),
    .Y(_01986_));
 sky130_fd_sc_hd__o22a_1 _20299_ (.A1(_04184_),
    .A2(_14236_),
    .B1(\reg_pc[23] ),
    .B2(\decoded_imm[23] ),
    .X(_04744_));
 sky130_fd_sc_hd__o21ai_1 _20300_ (.A1(_04178_),
    .A2(_14235_),
    .B1(_04736_),
    .Y(_04745_));
 sky130_fd_sc_hd__nand2_1 _20301_ (.A(_04744_),
    .B(_04745_),
    .Y(_04746_));
 sky130_fd_sc_hd__or2_1 _20302_ (.A(_04744_),
    .B(_04745_),
    .X(_04747_));
 sky130_fd_sc_hd__o2bb2a_1 _20303_ (.A1_N(_04737_),
    .A2_N(_01982_),
    .B1(_04738_),
    .B2(_01987_),
    .X(_04748_));
 sky130_fd_sc_hd__o21ai_4 _20304_ (.A1(_04718_),
    .A2(_01981_),
    .B1(_04748_),
    .Y(_04749_));
 sky130_fd_sc_hd__a31o_1 _20305_ (.A1(_04732_),
    .A2(_04746_),
    .A3(_04747_),
    .B1(_04749_),
    .X(_01988_));
 sky130_fd_sc_hd__buf_1 _20306_ (.A(_04664_),
    .X(_04750_));
 sky130_fd_sc_hd__or2_1 _20307_ (.A(_04425_),
    .B(_04750_),
    .X(_01989_));
 sky130_fd_sc_hd__buf_1 _20308_ (.A(_04620_),
    .X(_04751_));
 sky130_fd_sc_hd__or2_1 _20309_ (.A(_12123_),
    .B(_04741_),
    .X(_04752_));
 sky130_fd_sc_hd__o221a_1 _20310_ (.A1(_12091_),
    .A2(_04721_),
    .B1(_04751_),
    .B2(_12413_),
    .C1(_04752_),
    .X(_01993_));
 sky130_fd_sc_hd__buf_1 _20311_ (.A(_13299_),
    .X(_04753_));
 sky130_fd_sc_hd__clkbuf_2 _20312_ (.A(_11815_),
    .X(_04754_));
 sky130_fd_sc_hd__nand2_1 _20313_ (.A(_04688_),
    .B(\cpuregs_rs1[24] ),
    .Y(_04755_));
 sky130_fd_sc_hd__o221a_2 _20314_ (.A1(_04753_),
    .A2(_14220_),
    .B1(_11631_),
    .B2(_04754_),
    .C1(_04755_),
    .X(_01995_));
 sky130_fd_sc_hd__o21ai_2 _20315_ (.A1(_04184_),
    .A2(_14237_),
    .B1(_04746_),
    .Y(_04756_));
 sky130_fd_sc_hd__o22a_1 _20316_ (.A1(_04190_),
    .A2(_14239_),
    .B1(\reg_pc[24] ),
    .B2(_13925_),
    .X(_04757_));
 sky130_fd_sc_hd__or2_1 _20317_ (.A(_04756_),
    .B(_04757_),
    .X(_04758_));
 sky130_fd_sc_hd__nand2_1 _20318_ (.A(_04756_),
    .B(_04757_),
    .Y(_04759_));
 sky130_fd_sc_hd__clkbuf_4 _20319_ (.A(_14038_),
    .X(_04760_));
 sky130_fd_sc_hd__o2bb2a_1 _20320_ (.A1_N(_04737_),
    .A2_N(_01991_),
    .B1(_04738_),
    .B2(_01996_),
    .X(_04761_));
 sky130_fd_sc_hd__o21ai_4 _20321_ (.A1(_04760_),
    .A2(_01990_),
    .B1(_04761_),
    .Y(_04762_));
 sky130_fd_sc_hd__a31o_1 _20322_ (.A1(_04732_),
    .A2(_04758_),
    .A3(_04759_),
    .B1(_04762_),
    .X(_01997_));
 sky130_fd_sc_hd__or2_1 _20323_ (.A(_04442_),
    .B(_04750_),
    .X(_01998_));
 sky130_fd_sc_hd__clkbuf_2 _20324_ (.A(_04630_),
    .X(_04763_));
 sky130_fd_sc_hd__or2_1 _20325_ (.A(_12122_),
    .B(_04741_),
    .X(_04764_));
 sky130_fd_sc_hd__o221a_1 _20326_ (.A1(_12090_),
    .A2(_04763_),
    .B1(_04751_),
    .B2(_12412_),
    .C1(_04764_),
    .X(_02002_));
 sky130_fd_sc_hd__clkbuf_4 _20327_ (.A(_04448_),
    .X(_04765_));
 sky130_fd_sc_hd__buf_1 _20328_ (.A(_04488_),
    .X(_04766_));
 sky130_fd_sc_hd__buf_1 _20329_ (.A(_04490_),
    .X(_04767_));
 sky130_fd_sc_hd__a22o_1 _20330_ (.A1(_04766_),
    .A2(\timer[25] ),
    .B1(\irq_mask[25] ),
    .B2(_04767_),
    .X(_04768_));
 sky130_fd_sc_hd__a21oi_4 _20331_ (.A1(_04765_),
    .A2(\cpuregs_rs1[25] ),
    .B1(_04768_),
    .Y(_02004_));
 sky130_fd_sc_hd__nor2_1 _20332_ (.A(\reg_pc[25] ),
    .B(\decoded_imm[25] ),
    .Y(_04769_));
 sky130_fd_sc_hd__a21oi_2 _20333_ (.A1(\reg_pc[25] ),
    .A2(_13927_),
    .B1(_04769_),
    .Y(_04770_));
 sky130_fd_sc_hd__o21ai_1 _20334_ (.A1(_04190_),
    .A2(_14240_),
    .B1(_04759_),
    .Y(_04771_));
 sky130_fd_sc_hd__or2_1 _20335_ (.A(_04770_),
    .B(_04771_),
    .X(_04772_));
 sky130_fd_sc_hd__a21oi_1 _20336_ (.A1(_04770_),
    .A2(_04771_),
    .B1(_14061_),
    .Y(_04773_));
 sky130_fd_sc_hd__o22ai_4 _20337_ (.A1(_04591_),
    .A2(_01999_),
    .B1(_04529_),
    .B2(_02005_),
    .Y(_04774_));
 sky130_fd_sc_hd__a221o_1 _20338_ (.A1(_12367_),
    .A2(_02000_),
    .B1(_04772_),
    .B2(_04773_),
    .C1(_04774_),
    .X(_02006_));
 sky130_fd_sc_hd__or2_1 _20339_ (.A(_04461_),
    .B(_04750_),
    .X(_02007_));
 sky130_fd_sc_hd__or2_1 _20340_ (.A(_12121_),
    .B(_04741_),
    .X(_04775_));
 sky130_fd_sc_hd__o221a_1 _20341_ (.A1(_12089_),
    .A2(_04763_),
    .B1(_04751_),
    .B2(_12411_),
    .C1(_04775_),
    .X(_02011_));
 sky130_fd_sc_hd__nand2_1 _20342_ (.A(_04486_),
    .B(\cpuregs_rs1[26] ),
    .Y(_04776_));
 sky130_fd_sc_hd__o221a_2 _20343_ (.A1(_04753_),
    .A2(_14169_),
    .B1(_11632_),
    .B2(_04754_),
    .C1(_04776_),
    .X(_02013_));
 sky130_fd_sc_hd__o32a_1 _20344_ (.A1(_04189_),
    .A2(_14239_),
    .A3(_04769_),
    .B1(_04194_),
    .B2(_14241_),
    .X(_04777_));
 sky130_vsdinv _20345_ (.A(_04777_),
    .Y(_04778_));
 sky130_fd_sc_hd__a31o_1 _20346_ (.A1(_04757_),
    .A2(_04770_),
    .A3(_04756_),
    .B1(_04778_),
    .X(_04779_));
 sky130_fd_sc_hd__o22a_1 _20347_ (.A1(_04200_),
    .A2(_14242_),
    .B1(\reg_pc[26] ),
    .B2(_13931_),
    .X(_04780_));
 sky130_fd_sc_hd__or2_1 _20348_ (.A(_04779_),
    .B(_04780_),
    .X(_04781_));
 sky130_fd_sc_hd__nand2_1 _20349_ (.A(_04779_),
    .B(_04780_),
    .Y(_04782_));
 sky130_fd_sc_hd__o2bb2a_1 _20350_ (.A1_N(_04737_),
    .A2_N(_02009_),
    .B1(_04738_),
    .B2(_02014_),
    .X(_04783_));
 sky130_fd_sc_hd__o21ai_4 _20351_ (.A1(_04760_),
    .A2(_02008_),
    .B1(_04783_),
    .Y(_04784_));
 sky130_fd_sc_hd__a31o_1 _20352_ (.A1(_04732_),
    .A2(_04781_),
    .A3(_04782_),
    .B1(_04784_),
    .X(_02015_));
 sky130_fd_sc_hd__or2_1 _20353_ (.A(_04476_),
    .B(_04750_),
    .X(_02016_));
 sky130_fd_sc_hd__buf_1 _20354_ (.A(_04651_),
    .X(_04785_));
 sky130_fd_sc_hd__or2_1 _20355_ (.A(_12120_),
    .B(_04785_),
    .X(_04786_));
 sky130_fd_sc_hd__o221a_1 _20356_ (.A1(_12088_),
    .A2(_04763_),
    .B1(_04751_),
    .B2(_12410_),
    .C1(_04786_),
    .X(_02020_));
 sky130_fd_sc_hd__a22o_1 _20357_ (.A1(_04766_),
    .A2(\timer[27] ),
    .B1(\irq_mask[27] ),
    .B2(_04767_),
    .X(_04787_));
 sky130_fd_sc_hd__a21oi_4 _20358_ (.A1(_04765_),
    .A2(\cpuregs_rs1[27] ),
    .B1(_04787_),
    .Y(_02022_));
 sky130_fd_sc_hd__nor2_1 _20359_ (.A(\reg_pc[27] ),
    .B(\decoded_imm[27] ),
    .Y(_04788_));
 sky130_fd_sc_hd__a21oi_2 _20360_ (.A1(\reg_pc[27] ),
    .A2(_13933_),
    .B1(_04788_),
    .Y(_04789_));
 sky130_fd_sc_hd__o21ai_1 _20361_ (.A1(_04200_),
    .A2(_14243_),
    .B1(_04782_),
    .Y(_04790_));
 sky130_fd_sc_hd__or2_1 _20362_ (.A(_04789_),
    .B(_04790_),
    .X(_04791_));
 sky130_fd_sc_hd__a21oi_1 _20363_ (.A1(_04789_),
    .A2(_04790_),
    .B1(_14061_),
    .Y(_04792_));
 sky130_fd_sc_hd__o22ai_4 _20364_ (.A1(_04591_),
    .A2(_02017_),
    .B1(_04438_),
    .B2(_02023_),
    .Y(_04793_));
 sky130_fd_sc_hd__a221o_1 _20365_ (.A1(_12367_),
    .A2(_02018_),
    .B1(_04791_),
    .B2(_04792_),
    .C1(_04793_),
    .X(_02024_));
 sky130_fd_sc_hd__buf_1 _20366_ (.A(_04664_),
    .X(_04794_));
 sky130_fd_sc_hd__or2_1 _20367_ (.A(_04500_),
    .B(_04794_),
    .X(_02025_));
 sky130_fd_sc_hd__clkbuf_2 _20368_ (.A(_11743_),
    .X(_04795_));
 sky130_fd_sc_hd__or2_1 _20369_ (.A(_12119_),
    .B(_04785_),
    .X(_04796_));
 sky130_fd_sc_hd__o221a_1 _20370_ (.A1(_12087_),
    .A2(_04763_),
    .B1(_04795_),
    .B2(_12409_),
    .C1(_04796_),
    .X(_02029_));
 sky130_fd_sc_hd__nand2_1 _20371_ (.A(_04486_),
    .B(\cpuregs_rs1[28] ),
    .Y(_04797_));
 sky130_fd_sc_hd__o221a_1 _20372_ (.A1(_04753_),
    .A2(_14222_),
    .B1(_11650_),
    .B2(_04754_),
    .C1(_04797_),
    .X(_02031_));
 sky130_fd_sc_hd__o2bb2a_1 _20373_ (.A1_N(_04468_),
    .A2_N(_02027_),
    .B1(_14160_),
    .B2(_02032_),
    .X(_04798_));
 sky130_fd_sc_hd__o32a_1 _20374_ (.A1(_04199_),
    .A2(_14242_),
    .A3(_04788_),
    .B1(_04208_),
    .B2(_14244_),
    .X(_04799_));
 sky130_vsdinv _20375_ (.A(_04799_),
    .Y(_04800_));
 sky130_fd_sc_hd__a31o_1 _20376_ (.A1(_04780_),
    .A2(_04789_),
    .A3(_04779_),
    .B1(_04800_),
    .X(_04801_));
 sky130_fd_sc_hd__nor2_1 _20377_ (.A(_12052_),
    .B(\decoded_imm[28] ),
    .Y(_04802_));
 sky130_fd_sc_hd__a21oi_2 _20378_ (.A1(_12052_),
    .A2(_13935_),
    .B1(_04802_),
    .Y(_04803_));
 sky130_vsdinv _20379_ (.A(_04801_),
    .Y(_04804_));
 sky130_vsdinv _20380_ (.A(_04803_),
    .Y(_04805_));
 sky130_fd_sc_hd__a221o_4 _20381_ (.A1(_04801_),
    .A2(_04803_),
    .B1(_04804_),
    .B2(_04805_),
    .C1(_04440_),
    .X(_04806_));
 sky130_fd_sc_hd__o211ai_4 _20382_ (.A1(_04455_),
    .A2(_02026_),
    .B1(_04798_),
    .C1(_04806_),
    .Y(_02033_));
 sky130_fd_sc_hd__or2_1 _20383_ (.A(_04516_),
    .B(_04794_),
    .X(_02034_));
 sky130_fd_sc_hd__or2_1 _20384_ (.A(_12118_),
    .B(_04785_),
    .X(_04807_));
 sky130_fd_sc_hd__o221a_1 _20385_ (.A1(_12086_),
    .A2(_13334_),
    .B1(_04795_),
    .B2(_12408_),
    .C1(_04807_),
    .X(_02038_));
 sky130_fd_sc_hd__a22o_1 _20386_ (.A1(_04766_),
    .A2(\timer[29] ),
    .B1(\irq_mask[29] ),
    .B2(_04767_),
    .X(_04808_));
 sky130_fd_sc_hd__a21oi_4 _20387_ (.A1(_04765_),
    .A2(\cpuregs_rs1[29] ),
    .B1(_04808_),
    .Y(_02040_));
 sky130_fd_sc_hd__o2bb2a_1 _20388_ (.A1_N(_04468_),
    .A2_N(_02036_),
    .B1(_14160_),
    .B2(_02041_),
    .X(_04809_));
 sky130_fd_sc_hd__o22a_2 _20389_ (.A1(_04212_),
    .A2(_14246_),
    .B1(_04804_),
    .B2(_04802_),
    .X(_04810_));
 sky130_vsdinv _20390_ (.A(_04810_),
    .Y(_04811_));
 sky130_fd_sc_hd__nor2_2 _20391_ (.A(\reg_pc[29] ),
    .B(\decoded_imm[29] ),
    .Y(_04812_));
 sky130_fd_sc_hd__a21oi_2 _20392_ (.A1(\reg_pc[29] ),
    .A2(_13937_),
    .B1(_04812_),
    .Y(_04813_));
 sky130_vsdinv _20393_ (.A(_04813_),
    .Y(_04814_));
 sky130_fd_sc_hd__a221o_2 _20394_ (.A1(_04811_),
    .A2(_04813_),
    .B1(_04810_),
    .B2(_04814_),
    .C1(_11734_),
    .X(_04815_));
 sky130_fd_sc_hd__o211ai_4 _20395_ (.A1(_04455_),
    .A2(_02035_),
    .B1(_04809_),
    .C1(_04815_),
    .Y(_02042_));
 sky130_fd_sc_hd__or2_1 _20396_ (.A(_04531_),
    .B(_04794_),
    .X(_02043_));
 sky130_fd_sc_hd__or2_1 _20397_ (.A(_12117_),
    .B(_04785_),
    .X(_04816_));
 sky130_fd_sc_hd__o221a_1 _20398_ (.A1(_12085_),
    .A2(_13334_),
    .B1(_04795_),
    .B2(_12407_),
    .C1(_04816_),
    .X(_02047_));
 sky130_fd_sc_hd__nand2_1 _20399_ (.A(_04486_),
    .B(\cpuregs_rs1[30] ),
    .Y(_04817_));
 sky130_fd_sc_hd__o221a_2 _20400_ (.A1(_04753_),
    .A2(_14224_),
    .B1(_11651_),
    .B2(_04754_),
    .C1(_04817_),
    .X(_02049_));
 sky130_fd_sc_hd__o22a_1 _20401_ (.A1(_04227_),
    .A2(_14248_),
    .B1(_12048_),
    .B2(\decoded_imm[30] ),
    .X(_04818_));
 sky130_fd_sc_hd__o22ai_2 _20402_ (.A1(_04222_),
    .A2(_14247_),
    .B1(_04810_),
    .B2(_04812_),
    .Y(_04819_));
 sky130_fd_sc_hd__or2_1 _20403_ (.A(_04818_),
    .B(_04819_),
    .X(_04820_));
 sky130_fd_sc_hd__nand2_1 _20404_ (.A(_04818_),
    .B(_04819_),
    .Y(_04821_));
 sky130_fd_sc_hd__o2bb2a_1 _20405_ (.A1_N(_12366_),
    .A2_N(_02045_),
    .B1(_11572_),
    .B2(_02050_),
    .X(_04822_));
 sky130_fd_sc_hd__o21ai_2 _20406_ (.A1(_04760_),
    .A2(_02044_),
    .B1(_04822_),
    .Y(_04823_));
 sky130_fd_sc_hd__a31o_1 _20407_ (.A1(_11726_),
    .A2(_04820_),
    .A3(_04821_),
    .B1(_04823_),
    .X(_02051_));
 sky130_fd_sc_hd__or2_1 _20408_ (.A(_04545_),
    .B(_04794_),
    .X(_02052_));
 sky130_fd_sc_hd__or2_1 _20409_ (.A(_12116_),
    .B(_04483_),
    .X(_04824_));
 sky130_fd_sc_hd__o221a_1 _20410_ (.A1(_12211_),
    .A2(_13334_),
    .B1(_04795_),
    .B2(_12502_),
    .C1(_04824_),
    .X(_02056_));
 sky130_fd_sc_hd__a22o_1 _20411_ (.A1(_04766_),
    .A2(\timer[31] ),
    .B1(\irq_mask[31] ),
    .B2(_04767_),
    .X(_04825_));
 sky130_fd_sc_hd__a21oi_4 _20412_ (.A1(_04765_),
    .A2(\cpuregs_rs1[31] ),
    .B1(_04825_),
    .Y(_02058_));
 sky130_fd_sc_hd__o21ai_1 _20413_ (.A1(_04227_),
    .A2(_14249_),
    .B1(_04821_),
    .Y(_04826_));
 sky130_fd_sc_hd__a221o_1 _20414_ (.A1(_12046_),
    .A2(_13939_),
    .B1(_04232_),
    .B2(\decoded_imm[31] ),
    .C1(_04826_),
    .X(_04827_));
 sky130_fd_sc_hd__o221ai_1 _20415_ (.A1(_12046_),
    .A2(\decoded_imm[31] ),
    .B1(_04232_),
    .B2(_13940_),
    .C1(_04826_),
    .Y(_04828_));
 sky130_fd_sc_hd__o2bb2a_1 _20416_ (.A1_N(_12366_),
    .A2_N(_02054_),
    .B1(_11572_),
    .B2(_02059_),
    .X(_04829_));
 sky130_fd_sc_hd__o21ai_2 _20417_ (.A1(_04760_),
    .A2(_02053_),
    .B1(_04829_),
    .Y(_04830_));
 sky130_fd_sc_hd__a31o_1 _20418_ (.A1(_11726_),
    .A2(_04827_),
    .A3(_04828_),
    .B1(_04830_),
    .X(_02060_));
 sky130_fd_sc_hd__or2_1 _20419_ (.A(\decoded_rd[4] ),
    .B(net410),
    .X(_02061_));
 sky130_vsdinv _20420_ (.A(_13991_),
    .Y(_02062_));
 sky130_fd_sc_hd__o21ai_1 _20421_ (.A1(_14062_),
    .A2(_02064_),
    .B1(_14161_),
    .Y(_02065_));
 sky130_fd_sc_hd__nor3_1 _20422_ (.A(_11673_),
    .B(_02410_),
    .C(_00308_),
    .Y(_02066_));
 sky130_fd_sc_hd__clkbuf_1 _20423_ (.A(_01706_),
    .X(_02067_));
 sky130_fd_sc_hd__nor2_1 _20424_ (.A(_11982_),
    .B(_14157_),
    .Y(_04831_));
 sky130_fd_sc_hd__o211ai_1 _20425_ (.A1(_14062_),
    .A2(_04831_),
    .B1(_14161_),
    .C1(_14040_),
    .Y(_02068_));
 sky130_fd_sc_hd__clkbuf_4 _20426_ (.A(_11779_),
    .X(_04832_));
 sky130_fd_sc_hd__or2_1 _20427_ (.A(_11575_),
    .B(_12559_),
    .X(_04833_));
 sky130_fd_sc_hd__and3_4 _20428_ (.A(_04832_),
    .B(_11777_),
    .C(_04833_),
    .X(_02069_));
 sky130_vsdinv _20429_ (.A(_04833_),
    .Y(_04834_));
 sky130_fd_sc_hd__clkbuf_2 _20430_ (.A(_04834_),
    .X(_04835_));
 sky130_fd_sc_hd__clkbuf_2 _20431_ (.A(_04835_),
    .X(_04836_));
 sky130_fd_sc_hd__buf_2 _20432_ (.A(_11775_),
    .X(_04837_));
 sky130_fd_sc_hd__a22o_1 _20433_ (.A1(_02070_),
    .A2(_04836_),
    .B1(_04837_),
    .B2(_13781_),
    .X(_04838_));
 sky130_fd_sc_hd__a31o_1 _20434_ (.A1(_12360_),
    .A2(\irq_pending[0] ),
    .A3(_11771_),
    .B1(_04838_),
    .X(_02071_));
 sky130_fd_sc_hd__clkbuf_2 _20435_ (.A(_04834_),
    .X(_04839_));
 sky130_fd_sc_hd__buf_1 _20436_ (.A(_04839_),
    .X(_04840_));
 sky130_fd_sc_hd__and3_1 _20437_ (.A(_12357_),
    .B(_12358_),
    .C(_11771_),
    .X(_04841_));
 sky130_fd_sc_hd__a221o_1 _20438_ (.A1(_01465_),
    .A2(_04840_),
    .B1(_11785_),
    .B2(\reg_next_pc[1] ),
    .C1(_04841_),
    .X(_02072_));
 sky130_fd_sc_hd__and3_1 _20439_ (.A(_12354_),
    .B(_12355_),
    .C(_11771_),
    .X(_04842_));
 sky130_fd_sc_hd__a221o_1 _20440_ (.A1(_00293_),
    .A2(_04840_),
    .B1(_11785_),
    .B2(\reg_next_pc[2] ),
    .C1(_04842_),
    .X(_02074_));
 sky130_fd_sc_hd__nor2_2 _20441_ (.A(_14265_),
    .B(_14258_),
    .Y(_04843_));
 sky130_fd_sc_hd__a21oi_2 _20442_ (.A1(_14265_),
    .A2(_02073_),
    .B1(_04843_),
    .Y(_02075_));
 sky130_fd_sc_hd__buf_1 _20443_ (.A(_04837_),
    .X(_04844_));
 sky130_fd_sc_hd__nor3_4 _20444_ (.A(_11873_),
    .B(_11622_),
    .C(_04832_),
    .Y(_04845_));
 sky130_fd_sc_hd__a221o_1 _20445_ (.A1(_01468_),
    .A2(_04840_),
    .B1(_04844_),
    .B2(\reg_next_pc[3] ),
    .C1(_04845_),
    .X(_02076_));
 sky130_fd_sc_hd__nand2_2 _20446_ (.A(\reg_pc[4] ),
    .B(_04843_),
    .Y(_04846_));
 sky130_fd_sc_hd__o21a_1 _20447_ (.A1(_12081_),
    .A2(_04843_),
    .B1(_04846_),
    .X(_02077_));
 sky130_fd_sc_hd__nor3_4 _20448_ (.A(_11872_),
    .B(_11639_),
    .C(_04832_),
    .Y(_04847_));
 sky130_fd_sc_hd__a221o_1 _20449_ (.A1(_01472_),
    .A2(_04840_),
    .B1(_04844_),
    .B2(\reg_next_pc[4] ),
    .C1(_04847_),
    .X(_02078_));
 sky130_fd_sc_hd__nor2_2 _20450_ (.A(_14276_),
    .B(_04846_),
    .Y(_04848_));
 sky130_fd_sc_hd__a21oi_1 _20451_ (.A1(_14276_),
    .A2(_04846_),
    .B1(_04848_),
    .Y(_02079_));
 sky130_fd_sc_hd__buf_1 _20452_ (.A(_04839_),
    .X(_04849_));
 sky130_fd_sc_hd__buf_1 _20453_ (.A(_11770_),
    .X(_04850_));
 sky130_fd_sc_hd__buf_1 _20454_ (.A(_04850_),
    .X(_04851_));
 sky130_fd_sc_hd__and3_2 _20455_ (.A(_11637_),
    .B(_12346_),
    .C(_04851_),
    .X(_04852_));
 sky130_fd_sc_hd__a221o_1 _20456_ (.A1(_01476_),
    .A2(_04849_),
    .B1(_04844_),
    .B2(\reg_next_pc[5] ),
    .C1(_04852_),
    .X(_02080_));
 sky130_fd_sc_hd__nand2_1 _20457_ (.A(\reg_pc[6] ),
    .B(_04848_),
    .Y(_04853_));
 sky130_fd_sc_hd__o21a_1 _20458_ (.A1(_12076_),
    .A2(_04848_),
    .B1(_04853_),
    .X(_02081_));
 sky130_fd_sc_hd__nor3_4 _20459_ (.A(_11870_),
    .B(_11640_),
    .C(_04832_),
    .Y(_04854_));
 sky130_fd_sc_hd__a221o_1 _20460_ (.A1(_01479_),
    .A2(_04849_),
    .B1(_04844_),
    .B2(\reg_next_pc[6] ),
    .C1(_04854_),
    .X(_02082_));
 sky130_fd_sc_hd__or2_1 _20461_ (.A(_04080_),
    .B(_04853_),
    .X(_04855_));
 sky130_vsdinv _20462_ (.A(_04855_),
    .Y(_04856_));
 sky130_fd_sc_hd__a21oi_1 _20463_ (.A1(_04080_),
    .A2(_04853_),
    .B1(_04856_),
    .Y(_02083_));
 sky130_fd_sc_hd__buf_1 _20464_ (.A(_04837_),
    .X(_04857_));
 sky130_fd_sc_hd__and3_1 _20465_ (.A(_11638_),
    .B(_12342_),
    .C(_04851_),
    .X(_04858_));
 sky130_fd_sc_hd__a221o_1 _20466_ (.A1(_01482_),
    .A2(_04849_),
    .B1(_04857_),
    .B2(\reg_next_pc[7] ),
    .C1(_04858_),
    .X(_02084_));
 sky130_fd_sc_hd__or2_2 _20467_ (.A(_04085_),
    .B(_04855_),
    .X(_04859_));
 sky130_fd_sc_hd__o21a_1 _20468_ (.A1(\reg_pc[8] ),
    .A2(_04856_),
    .B1(_04859_),
    .X(_02085_));
 sky130_fd_sc_hd__buf_4 _20469_ (.A(_11780_),
    .X(_04860_));
 sky130_fd_sc_hd__nor3_4 _20470_ (.A(_11866_),
    .B(_11658_),
    .C(_04860_),
    .Y(_04861_));
 sky130_fd_sc_hd__a221o_1 _20471_ (.A1(_01485_),
    .A2(_04849_),
    .B1(_04857_),
    .B2(\reg_next_pc[8] ),
    .C1(_04861_),
    .X(_02086_));
 sky130_fd_sc_hd__or2_1 _20472_ (.A(_04095_),
    .B(_04859_),
    .X(_04862_));
 sky130_vsdinv _20473_ (.A(_04862_),
    .Y(_04863_));
 sky130_fd_sc_hd__a21oi_2 _20474_ (.A1(_04095_),
    .A2(_04859_),
    .B1(_04863_),
    .Y(_02087_));
 sky130_fd_sc_hd__buf_1 _20475_ (.A(_04839_),
    .X(_04864_));
 sky130_fd_sc_hd__and3_1 _20476_ (.A(_11656_),
    .B(_12336_),
    .C(_04851_),
    .X(_04865_));
 sky130_fd_sc_hd__a221o_1 _20477_ (.A1(_01488_),
    .A2(_04864_),
    .B1(_04857_),
    .B2(\reg_next_pc[9] ),
    .C1(_04865_),
    .X(_02088_));
 sky130_fd_sc_hd__or2_1 _20478_ (.A(_04102_),
    .B(_04862_),
    .X(_04866_));
 sky130_fd_sc_hd__o21a_1 _20479_ (.A1(\reg_pc[10] ),
    .A2(_04863_),
    .B1(_04866_),
    .X(_02089_));
 sky130_fd_sc_hd__nor3_4 _20480_ (.A(_11864_),
    .B(_11659_),
    .C(_04860_),
    .Y(_04867_));
 sky130_fd_sc_hd__a221o_1 _20481_ (.A1(_01491_),
    .A2(_04864_),
    .B1(_04857_),
    .B2(\reg_next_pc[10] ),
    .C1(_04867_),
    .X(_02090_));
 sky130_fd_sc_hd__or2_1 _20482_ (.A(_04108_),
    .B(_04866_),
    .X(_04868_));
 sky130_vsdinv _20483_ (.A(_04868_),
    .Y(_04869_));
 sky130_fd_sc_hd__a21oi_1 _20484_ (.A1(_04109_),
    .A2(_04866_),
    .B1(_04869_),
    .Y(_02091_));
 sky130_fd_sc_hd__clkbuf_4 _20485_ (.A(_11775_),
    .X(_04870_));
 sky130_fd_sc_hd__buf_1 _20486_ (.A(_04870_),
    .X(_04871_));
 sky130_fd_sc_hd__and3_1 _20487_ (.A(_11657_),
    .B(_12332_),
    .C(_04851_),
    .X(_04872_));
 sky130_fd_sc_hd__a221o_1 _20488_ (.A1(_01494_),
    .A2(_04864_),
    .B1(_04871_),
    .B2(\reg_next_pc[11] ),
    .C1(_04872_),
    .X(_02092_));
 sky130_fd_sc_hd__or2_1 _20489_ (.A(_04114_),
    .B(_04868_),
    .X(_04873_));
 sky130_fd_sc_hd__o21a_1 _20490_ (.A1(\reg_pc[12] ),
    .A2(_04869_),
    .B1(_04873_),
    .X(_02093_));
 sky130_fd_sc_hd__nor3_4 _20491_ (.A(_11861_),
    .B(_11646_),
    .C(_04860_),
    .Y(_04874_));
 sky130_fd_sc_hd__a221o_1 _20492_ (.A1(_01497_),
    .A2(_04864_),
    .B1(_04871_),
    .B2(\reg_next_pc[12] ),
    .C1(_04874_),
    .X(_02094_));
 sky130_fd_sc_hd__or2_1 _20493_ (.A(_04119_),
    .B(_04873_),
    .X(_04875_));
 sky130_vsdinv _20494_ (.A(_04875_),
    .Y(_04876_));
 sky130_fd_sc_hd__a21oi_1 _20495_ (.A1(_04120_),
    .A2(_04873_),
    .B1(_04876_),
    .Y(_02095_));
 sky130_fd_sc_hd__clkbuf_2 _20496_ (.A(_04839_),
    .X(_04877_));
 sky130_fd_sc_hd__buf_1 _20497_ (.A(_04850_),
    .X(_04878_));
 sky130_fd_sc_hd__and3_1 _20498_ (.A(_11644_),
    .B(_12326_),
    .C(_04878_),
    .X(_04879_));
 sky130_fd_sc_hd__a221o_1 _20499_ (.A1(_01500_),
    .A2(_04877_),
    .B1(_04871_),
    .B2(\reg_next_pc[13] ),
    .C1(_04879_),
    .X(_02096_));
 sky130_fd_sc_hd__or2_1 _20500_ (.A(_04127_),
    .B(_04875_),
    .X(_04880_));
 sky130_fd_sc_hd__o21a_1 _20501_ (.A1(\reg_pc[14] ),
    .A2(_04876_),
    .B1(_04880_),
    .X(_02097_));
 sky130_fd_sc_hd__nor3_4 _20502_ (.A(_11858_),
    .B(_11647_),
    .C(_04860_),
    .Y(_04881_));
 sky130_fd_sc_hd__a221o_1 _20503_ (.A1(_01503_),
    .A2(_04877_),
    .B1(_04871_),
    .B2(\reg_next_pc[14] ),
    .C1(_04881_),
    .X(_02098_));
 sky130_fd_sc_hd__or2_1 _20504_ (.A(_04132_),
    .B(_04880_),
    .X(_04882_));
 sky130_vsdinv _20505_ (.A(_04882_),
    .Y(_04883_));
 sky130_fd_sc_hd__a21oi_1 _20506_ (.A1(_04133_),
    .A2(_04880_),
    .B1(_04883_),
    .Y(_02099_));
 sky130_fd_sc_hd__buf_1 _20507_ (.A(_04870_),
    .X(_04884_));
 sky130_fd_sc_hd__and3_1 _20508_ (.A(_11645_),
    .B(_12322_),
    .C(_04878_),
    .X(_04885_));
 sky130_fd_sc_hd__a221o_1 _20509_ (.A1(_01506_),
    .A2(_04877_),
    .B1(_04884_),
    .B2(\reg_next_pc[15] ),
    .C1(_04885_),
    .X(_02100_));
 sky130_fd_sc_hd__or2_2 _20510_ (.A(_04138_),
    .B(_04882_),
    .X(_04886_));
 sky130_fd_sc_hd__o21a_1 _20511_ (.A1(\reg_pc[16] ),
    .A2(_04883_),
    .B1(_04886_),
    .X(_02101_));
 sky130_fd_sc_hd__buf_4 _20512_ (.A(_11779_),
    .X(_04887_));
 sky130_fd_sc_hd__nor3_4 _20513_ (.A(_11853_),
    .B(_11627_),
    .C(_04887_),
    .Y(_04888_));
 sky130_fd_sc_hd__a221o_1 _20514_ (.A1(_01509_),
    .A2(_04877_),
    .B1(_04884_),
    .B2(\reg_next_pc[16] ),
    .C1(_04888_),
    .X(_02102_));
 sky130_fd_sc_hd__or2_1 _20515_ (.A(_04146_),
    .B(_04886_),
    .X(_04889_));
 sky130_vsdinv _20516_ (.A(_04889_),
    .Y(_04890_));
 sky130_fd_sc_hd__a21oi_1 _20517_ (.A1(_04146_),
    .A2(_04886_),
    .B1(_04890_),
    .Y(_02103_));
 sky130_fd_sc_hd__clkbuf_2 _20518_ (.A(_04835_),
    .X(_04891_));
 sky130_fd_sc_hd__nor3_4 _20519_ (.A(_11852_),
    .B(_11625_),
    .C(_04887_),
    .Y(_04892_));
 sky130_fd_sc_hd__a221o_1 _20520_ (.A1(_01512_),
    .A2(_04891_),
    .B1(_04884_),
    .B2(\reg_next_pc[17] ),
    .C1(_04892_),
    .X(_02104_));
 sky130_fd_sc_hd__or2_1 _20521_ (.A(_04153_),
    .B(_04889_),
    .X(_04893_));
 sky130_fd_sc_hd__o21a_1 _20522_ (.A1(\reg_pc[18] ),
    .A2(_04890_),
    .B1(_04893_),
    .X(_02105_));
 sky130_fd_sc_hd__and3_1 _20523_ (.A(_12312_),
    .B(_12313_),
    .C(_04878_),
    .X(_04894_));
 sky130_fd_sc_hd__a221o_1 _20524_ (.A1(_01515_),
    .A2(_04891_),
    .B1(_04884_),
    .B2(\reg_next_pc[18] ),
    .C1(_04894_),
    .X(_02106_));
 sky130_fd_sc_hd__or2_1 _20525_ (.A(_04160_),
    .B(_04893_),
    .X(_04895_));
 sky130_vsdinv _20526_ (.A(_04895_),
    .Y(_04896_));
 sky130_fd_sc_hd__a21oi_1 _20527_ (.A1(_04161_),
    .A2(_04893_),
    .B1(_04896_),
    .Y(_02107_));
 sky130_fd_sc_hd__buf_1 _20528_ (.A(_04870_),
    .X(_04897_));
 sky130_fd_sc_hd__nor3_4 _20529_ (.A(_11846_),
    .B(_11626_),
    .C(_04887_),
    .Y(_04898_));
 sky130_fd_sc_hd__a221o_1 _20530_ (.A1(_01518_),
    .A2(_04891_),
    .B1(_04897_),
    .B2(\reg_next_pc[19] ),
    .C1(_04898_),
    .X(_02108_));
 sky130_fd_sc_hd__or2_1 _20531_ (.A(_04166_),
    .B(_04895_),
    .X(_04899_));
 sky130_fd_sc_hd__o21a_1 _20532_ (.A1(\reg_pc[20] ),
    .A2(_04896_),
    .B1(_04899_),
    .X(_02109_));
 sky130_fd_sc_hd__and3_1 _20533_ (.A(_11662_),
    .B(_12306_),
    .C(_04878_),
    .X(_04900_));
 sky130_fd_sc_hd__a221o_1 _20534_ (.A1(_01521_),
    .A2(_04891_),
    .B1(_04897_),
    .B2(\reg_next_pc[20] ),
    .C1(_04900_),
    .X(_02110_));
 sky130_fd_sc_hd__or2_1 _20535_ (.A(_04171_),
    .B(_04899_),
    .X(_04901_));
 sky130_vsdinv _20536_ (.A(_04901_),
    .Y(_04902_));
 sky130_fd_sc_hd__a21oi_1 _20537_ (.A1(_04172_),
    .A2(_04899_),
    .B1(_04902_),
    .Y(_02111_));
 sky130_fd_sc_hd__clkbuf_2 _20538_ (.A(_04835_),
    .X(_04903_));
 sky130_fd_sc_hd__nor3_4 _20539_ (.A(_11845_),
    .B(_11664_),
    .C(_04887_),
    .Y(_04904_));
 sky130_fd_sc_hd__a221o_1 _20540_ (.A1(_01524_),
    .A2(_04903_),
    .B1(_04897_),
    .B2(\reg_next_pc[21] ),
    .C1(_04904_),
    .X(_02112_));
 sky130_fd_sc_hd__or2_1 _20541_ (.A(_04178_),
    .B(_04901_),
    .X(_04905_));
 sky130_fd_sc_hd__o21a_1 _20542_ (.A1(\reg_pc[22] ),
    .A2(_04902_),
    .B1(_04905_),
    .X(_02113_));
 sky130_fd_sc_hd__buf_1 _20543_ (.A(_04850_),
    .X(_04906_));
 sky130_fd_sc_hd__and3_1 _20544_ (.A(_11663_),
    .B(_12301_),
    .C(_04906_),
    .X(_04907_));
 sky130_fd_sc_hd__a221o_1 _20545_ (.A1(_01527_),
    .A2(_04903_),
    .B1(_04897_),
    .B2(\reg_next_pc[22] ),
    .C1(_04907_),
    .X(_02114_));
 sky130_fd_sc_hd__or2_1 _20546_ (.A(_04183_),
    .B(_04905_),
    .X(_04908_));
 sky130_vsdinv _20547_ (.A(_04908_),
    .Y(_04909_));
 sky130_fd_sc_hd__a21oi_1 _20548_ (.A1(_04184_),
    .A2(_04905_),
    .B1(_04909_),
    .Y(_02115_));
 sky130_fd_sc_hd__clkbuf_2 _20549_ (.A(_04870_),
    .X(_04910_));
 sky130_fd_sc_hd__buf_4 _20550_ (.A(_11779_),
    .X(_04911_));
 sky130_fd_sc_hd__nor3_4 _20551_ (.A(_11839_),
    .B(_11665_),
    .C(_04911_),
    .Y(_04912_));
 sky130_fd_sc_hd__a221o_1 _20552_ (.A1(_01530_),
    .A2(_04903_),
    .B1(_04910_),
    .B2(\reg_next_pc[23] ),
    .C1(_04912_),
    .X(_02116_));
 sky130_fd_sc_hd__or2_2 _20553_ (.A(_04190_),
    .B(_04908_),
    .X(_04913_));
 sky130_fd_sc_hd__o21a_1 _20554_ (.A1(\reg_pc[24] ),
    .A2(_04909_),
    .B1(_04913_),
    .X(_02117_));
 sky130_fd_sc_hd__and3_1 _20555_ (.A(_11631_),
    .B(_12293_),
    .C(_04906_),
    .X(_04914_));
 sky130_fd_sc_hd__a221o_1 _20556_ (.A1(_01533_),
    .A2(_04903_),
    .B1(_04910_),
    .B2(\reg_next_pc[24] ),
    .C1(_04914_),
    .X(_02118_));
 sky130_fd_sc_hd__or2_1 _20557_ (.A(_04194_),
    .B(_04913_),
    .X(_04915_));
 sky130_vsdinv _20558_ (.A(_04915_),
    .Y(_04916_));
 sky130_fd_sc_hd__a21oi_1 _20559_ (.A1(_04194_),
    .A2(_04913_),
    .B1(_04916_),
    .Y(_02119_));
 sky130_fd_sc_hd__buf_1 _20560_ (.A(_04835_),
    .X(_04917_));
 sky130_fd_sc_hd__nor3_4 _20561_ (.A(_11838_),
    .B(_11633_),
    .C(_04911_),
    .Y(_04918_));
 sky130_fd_sc_hd__a221o_1 _20562_ (.A1(_01536_),
    .A2(_04917_),
    .B1(_04910_),
    .B2(\reg_next_pc[25] ),
    .C1(_04918_),
    .X(_02120_));
 sky130_fd_sc_hd__or2_1 _20563_ (.A(_04200_),
    .B(_04915_),
    .X(_04919_));
 sky130_fd_sc_hd__o21a_1 _20564_ (.A1(\reg_pc[26] ),
    .A2(_04916_),
    .B1(_04919_),
    .X(_02121_));
 sky130_fd_sc_hd__and3_1 _20565_ (.A(_11632_),
    .B(_12290_),
    .C(_04906_),
    .X(_04920_));
 sky130_fd_sc_hd__a221o_1 _20566_ (.A1(_01539_),
    .A2(_04917_),
    .B1(_04910_),
    .B2(\reg_next_pc[26] ),
    .C1(_04920_),
    .X(_02122_));
 sky130_fd_sc_hd__or2_1 _20567_ (.A(_04208_),
    .B(_04919_),
    .X(_04921_));
 sky130_vsdinv _20568_ (.A(_04921_),
    .Y(_04922_));
 sky130_fd_sc_hd__a21oi_1 _20569_ (.A1(_04208_),
    .A2(_04919_),
    .B1(_04922_),
    .Y(_02123_));
 sky130_fd_sc_hd__buf_1 _20570_ (.A(_11784_),
    .X(_04923_));
 sky130_fd_sc_hd__nor3_4 _20571_ (.A(_11834_),
    .B(_11634_),
    .C(_04911_),
    .Y(_04924_));
 sky130_fd_sc_hd__a221o_1 _20572_ (.A1(_01542_),
    .A2(_04917_),
    .B1(_04923_),
    .B2(\reg_next_pc[27] ),
    .C1(_04924_),
    .X(_02124_));
 sky130_fd_sc_hd__or2_2 _20573_ (.A(_04212_),
    .B(_04921_),
    .X(_04925_));
 sky130_fd_sc_hd__o21a_1 _20574_ (.A1(_12052_),
    .A2(_04922_),
    .B1(_04925_),
    .X(_02125_));
 sky130_fd_sc_hd__and3_1 _20575_ (.A(_11650_),
    .B(_12284_),
    .C(_04906_),
    .X(_04926_));
 sky130_fd_sc_hd__a221o_1 _20576_ (.A1(_01545_),
    .A2(_04917_),
    .B1(_04923_),
    .B2(\reg_next_pc[28] ),
    .C1(_04926_),
    .X(_02126_));
 sky130_fd_sc_hd__or2_1 _20577_ (.A(_04222_),
    .B(_04925_),
    .X(_04927_));
 sky130_vsdinv _20578_ (.A(_04927_),
    .Y(_04928_));
 sky130_fd_sc_hd__a21oi_1 _20579_ (.A1(_04222_),
    .A2(_04925_),
    .B1(_04928_),
    .Y(_02127_));
 sky130_fd_sc_hd__nor3_4 _20580_ (.A(_11833_),
    .B(_11652_),
    .C(_04911_),
    .Y(_04929_));
 sky130_fd_sc_hd__a221o_1 _20581_ (.A1(_01548_),
    .A2(_04836_),
    .B1(_04923_),
    .B2(\reg_next_pc[29] ),
    .C1(_04929_),
    .X(_02128_));
 sky130_fd_sc_hd__or2_1 _20582_ (.A(_04227_),
    .B(_04927_),
    .X(_04930_));
 sky130_fd_sc_hd__o21a_1 _20583_ (.A1(_12048_),
    .A2(_04928_),
    .B1(_04930_),
    .X(_02129_));
 sky130_fd_sc_hd__and3_1 _20584_ (.A(_11651_),
    .B(_12279_),
    .C(_04850_),
    .X(_04931_));
 sky130_fd_sc_hd__a221o_1 _20585_ (.A1(_01551_),
    .A2(_04836_),
    .B1(_04923_),
    .B2(\reg_next_pc[30] ),
    .C1(_04931_),
    .X(_02130_));
 sky130_fd_sc_hd__a32o_1 _20586_ (.A1(_12048_),
    .A2(_04928_),
    .A3(_04232_),
    .B1(_12046_),
    .B2(_04930_),
    .X(_02131_));
 sky130_fd_sc_hd__nor3_4 _20587_ (.A(_11814_),
    .B(_11653_),
    .C(_11780_),
    .Y(_04932_));
 sky130_fd_sc_hd__a221o_1 _20588_ (.A1(_01554_),
    .A2(_04836_),
    .B1(_04837_),
    .B2(\reg_next_pc[31] ),
    .C1(_04932_),
    .X(_02132_));
 sky130_fd_sc_hd__or2_4 _20589_ (.A(instr_xor),
    .B(instr_xori),
    .X(_04933_));
 sky130_fd_sc_hd__clkbuf_2 _20590_ (.A(_04933_),
    .X(_04934_));
 sky130_fd_sc_hd__or3_2 _20591_ (.A(is_compare),
    .B(_04934_),
    .C(_11756_),
    .X(_04935_));
 sky130_fd_sc_hd__nor2_8 _20592_ (.A(instr_and),
    .B(instr_andi),
    .Y(_04936_));
 sky130_fd_sc_hd__clkbuf_2 _20593_ (.A(_04936_),
    .X(_04937_));
 sky130_fd_sc_hd__buf_1 _20594_ (.A(_04937_),
    .X(_04938_));
 sky130_fd_sc_hd__nor2_8 _20595_ (.A(instr_or),
    .B(instr_ori),
    .Y(_04939_));
 sky130_fd_sc_hd__clkbuf_2 _20596_ (.A(_04939_),
    .X(_04940_));
 sky130_fd_sc_hd__or2_4 _20597_ (.A(instr_sll),
    .B(instr_slli),
    .X(_04941_));
 sky130_fd_sc_hd__buf_2 _20598_ (.A(_04941_),
    .X(_04942_));
 sky130_vsdinv _20599_ (.A(_04942_),
    .Y(_04943_));
 sky130_fd_sc_hd__and4b_4 _20600_ (.A_N(_04935_),
    .B(_04938_),
    .C(_04940_),
    .D(_04943_),
    .X(_02133_));
 sky130_fd_sc_hd__clkbuf_2 _20601_ (.A(_04933_),
    .X(_04944_));
 sky130_fd_sc_hd__clkbuf_2 _20602_ (.A(_11756_),
    .X(_04945_));
 sky130_fd_sc_hd__clkbuf_2 _20603_ (.A(_04945_),
    .X(_04946_));
 sky130_vsdinv _20604_ (.A(is_compare),
    .Y(_04947_));
 sky130_fd_sc_hd__nor2_1 _20605_ (.A(_12744_),
    .B(_13488_),
    .Y(_04948_));
 sky130_fd_sc_hd__buf_1 _20606_ (.A(_14069_),
    .X(_04949_));
 sky130_vsdinv _20607_ (.A(\alu_shl[0] ),
    .Y(_04950_));
 sky130_fd_sc_hd__o32a_1 _20608_ (.A1(_04949_),
    .A2(_14252_),
    .A3(_04937_),
    .B1(_04950_),
    .B2(_04943_),
    .X(_04951_));
 sky130_fd_sc_hd__o221ai_2 _20609_ (.A1(_00343_),
    .A2(_04947_),
    .B1(_04940_),
    .B2(_04948_),
    .C1(_04951_),
    .Y(_04952_));
 sky130_fd_sc_hd__a221o_1 _20610_ (.A1(_02591_),
    .A2(_04944_),
    .B1(\alu_shr[0] ),
    .B2(_04946_),
    .C1(_04952_),
    .X(_02134_));
 sky130_fd_sc_hd__clkbuf_2 _20611_ (.A(_11756_),
    .X(_04953_));
 sky130_fd_sc_hd__buf_1 _20612_ (.A(_04953_),
    .X(_04954_));
 sky130_fd_sc_hd__clkbuf_2 _20613_ (.A(_04941_),
    .X(_04955_));
 sky130_fd_sc_hd__buf_1 _20614_ (.A(_04955_),
    .X(_04956_));
 sky130_fd_sc_hd__a22o_1 _20615_ (.A1(\alu_shl[1] ),
    .A2(_04956_),
    .B1(_14113_),
    .B2(_04944_),
    .X(_04957_));
 sky130_fd_sc_hd__o32a_1 _20616_ (.A1(_13966_),
    .A2(_04414_),
    .A3(_04938_),
    .B1(_14112_),
    .B2(_04940_),
    .X(_04958_));
 sky130_vsdinv _20617_ (.A(_04958_),
    .Y(_04959_));
 sky130_fd_sc_hd__a211o_1 _20618_ (.A1(\alu_shr[1] ),
    .A2(_04954_),
    .B1(_04957_),
    .C1(_04959_),
    .X(_02135_));
 sky130_fd_sc_hd__a22o_1 _20619_ (.A1(\alu_shl[2] ),
    .A2(_04956_),
    .B1(_14122_),
    .B2(_04944_),
    .X(_04960_));
 sky130_fd_sc_hd__o32a_1 _20620_ (.A1(_13962_),
    .A2(_14266_),
    .A3(_04938_),
    .B1(_14121_),
    .B2(_04940_),
    .X(_04961_));
 sky130_vsdinv _20621_ (.A(_04961_),
    .Y(_04962_));
 sky130_fd_sc_hd__a211o_1 _20622_ (.A1(\alu_shr[2] ),
    .A2(_04954_),
    .B1(_04960_),
    .C1(_04962_),
    .X(_02136_));
 sky130_fd_sc_hd__a22o_1 _20623_ (.A1(\alu_shl[3] ),
    .A2(_04956_),
    .B1(_14115_),
    .B2(_04944_),
    .X(_04963_));
 sky130_fd_sc_hd__clkbuf_2 _20624_ (.A(_04939_),
    .X(_04964_));
 sky130_fd_sc_hd__buf_1 _20625_ (.A(_04964_),
    .X(_04965_));
 sky130_fd_sc_hd__o32a_1 _20626_ (.A1(_13957_),
    .A2(_14272_),
    .A3(_04938_),
    .B1(_14114_),
    .B2(_04965_),
    .X(_04966_));
 sky130_vsdinv _20627_ (.A(_04966_),
    .Y(_04967_));
 sky130_fd_sc_hd__a211o_1 _20628_ (.A1(\alu_shr[3] ),
    .A2(_04954_),
    .B1(_04963_),
    .C1(_04967_),
    .X(_02137_));
 sky130_fd_sc_hd__buf_1 _20629_ (.A(_04934_),
    .X(_04968_));
 sky130_fd_sc_hd__a22o_1 _20630_ (.A1(\alu_shl[4] ),
    .A2(_04956_),
    .B1(_14118_),
    .B2(_04968_),
    .X(_04969_));
 sky130_fd_sc_hd__buf_1 _20631_ (.A(_04937_),
    .X(_04970_));
 sky130_fd_sc_hd__o32a_1 _20632_ (.A1(_13953_),
    .A2(_14278_),
    .A3(_04970_),
    .B1(_14117_),
    .B2(_04965_),
    .X(_04971_));
 sky130_vsdinv _20633_ (.A(_04971_),
    .Y(_04972_));
 sky130_fd_sc_hd__a211o_1 _20634_ (.A1(\alu_shr[4] ),
    .A2(_04954_),
    .B1(_04969_),
    .C1(_04972_),
    .X(_02138_));
 sky130_fd_sc_hd__buf_1 _20635_ (.A(_04953_),
    .X(_04973_));
 sky130_fd_sc_hd__clkbuf_2 _20636_ (.A(_04942_),
    .X(_04974_));
 sky130_fd_sc_hd__buf_1 _20637_ (.A(_04974_),
    .X(_04975_));
 sky130_fd_sc_hd__a22o_1 _20638_ (.A1(\alu_shl[5] ),
    .A2(_04975_),
    .B1(_14109_),
    .B2(_04968_),
    .X(_04976_));
 sky130_fd_sc_hd__inv_2 _20639_ (.A(_12732_),
    .Y(_02330_));
 sky130_fd_sc_hd__o32a_1 _20640_ (.A1(_02330_),
    .A2(_04076_),
    .A3(_04970_),
    .B1(_14108_),
    .B2(_04965_),
    .X(_04977_));
 sky130_vsdinv _20641_ (.A(_04977_),
    .Y(_04978_));
 sky130_fd_sc_hd__a211o_1 _20642_ (.A1(\alu_shr[5] ),
    .A2(_04973_),
    .B1(_04976_),
    .C1(_04978_),
    .X(_02139_));
 sky130_fd_sc_hd__a22o_1 _20643_ (.A1(\alu_shl[6] ),
    .A2(_04975_),
    .B1(_14120_),
    .B2(_04968_),
    .X(_04979_));
 sky130_vsdinv _20644_ (.A(_12730_),
    .Y(_04980_));
 sky130_fd_sc_hd__buf_1 _20645_ (.A(_04980_),
    .X(_02333_));
 sky130_fd_sc_hd__o32a_1 _20646_ (.A1(_02333_),
    .A2(_04078_),
    .A3(_04970_),
    .B1(_14119_),
    .B2(_04965_),
    .X(_04981_));
 sky130_vsdinv _20647_ (.A(_04981_),
    .Y(_04982_));
 sky130_fd_sc_hd__a211o_1 _20648_ (.A1(\alu_shr[6] ),
    .A2(_04973_),
    .B1(_04979_),
    .C1(_04982_),
    .X(_02140_));
 sky130_fd_sc_hd__a22o_1 _20649_ (.A1(\alu_shl[7] ),
    .A2(_04975_),
    .B1(_14111_),
    .B2(_04968_),
    .X(_04983_));
 sky130_fd_sc_hd__inv_2 _20650_ (.A(_12727_),
    .Y(_02336_));
 sky130_fd_sc_hd__buf_1 _20651_ (.A(_04964_),
    .X(_04984_));
 sky130_fd_sc_hd__o32a_1 _20652_ (.A1(_02336_),
    .A2(_04087_),
    .A3(_04970_),
    .B1(_14110_),
    .B2(_04984_),
    .X(_04985_));
 sky130_vsdinv _20653_ (.A(_04985_),
    .Y(_04986_));
 sky130_fd_sc_hd__a211o_1 _20654_ (.A1(\alu_shr[7] ),
    .A2(_04973_),
    .B1(_04983_),
    .C1(_04986_),
    .X(_02141_));
 sky130_fd_sc_hd__buf_1 _20655_ (.A(_04934_),
    .X(_04987_));
 sky130_fd_sc_hd__a22o_1 _20656_ (.A1(\alu_shl[8] ),
    .A2(_04975_),
    .B1(_14136_),
    .B2(_04987_),
    .X(_04988_));
 sky130_fd_sc_hd__inv_2 _20657_ (.A(net368),
    .Y(_02339_));
 sky130_fd_sc_hd__buf_1 _20658_ (.A(_04937_),
    .X(_04989_));
 sky130_fd_sc_hd__o32a_1 _20659_ (.A1(_02339_),
    .A2(_04092_),
    .A3(_04989_),
    .B1(_14135_),
    .B2(_04984_),
    .X(_04990_));
 sky130_vsdinv _20660_ (.A(_04990_),
    .Y(_04991_));
 sky130_fd_sc_hd__a211o_1 _20661_ (.A1(\alu_shr[8] ),
    .A2(_04973_),
    .B1(_04988_),
    .C1(_04991_),
    .X(_02142_));
 sky130_fd_sc_hd__buf_1 _20662_ (.A(_04953_),
    .X(_04992_));
 sky130_fd_sc_hd__buf_1 _20663_ (.A(_04974_),
    .X(_04993_));
 sky130_fd_sc_hd__a22o_1 _20664_ (.A1(\alu_shl[9] ),
    .A2(_04993_),
    .B1(_14138_),
    .B2(_04987_),
    .X(_04994_));
 sky130_fd_sc_hd__inv_2 _20665_ (.A(_12723_),
    .Y(_02342_));
 sky130_fd_sc_hd__o32a_1 _20666_ (.A1(_02342_),
    .A2(_04105_),
    .A3(_04989_),
    .B1(_14137_),
    .B2(_04984_),
    .X(_04995_));
 sky130_vsdinv _20667_ (.A(_04995_),
    .Y(_04996_));
 sky130_fd_sc_hd__a211o_1 _20668_ (.A1(\alu_shr[9] ),
    .A2(_04992_),
    .B1(_04994_),
    .C1(_04996_),
    .X(_02143_));
 sky130_fd_sc_hd__a22o_1 _20669_ (.A1(\alu_shl[10] ),
    .A2(_04993_),
    .B1(_14140_),
    .B2(_04987_),
    .X(_04997_));
 sky130_fd_sc_hd__inv_2 _20670_ (.A(net339),
    .Y(_02345_));
 sky130_fd_sc_hd__o32a_1 _20671_ (.A1(_02345_),
    .A2(_04112_),
    .A3(_04989_),
    .B1(_14139_),
    .B2(_04984_),
    .X(_04998_));
 sky130_vsdinv _20672_ (.A(_04998_),
    .Y(_04999_));
 sky130_fd_sc_hd__a211o_1 _20673_ (.A1(\alu_shr[10] ),
    .A2(_04992_),
    .B1(_04997_),
    .C1(_04999_),
    .X(_02144_));
 sky130_fd_sc_hd__a22o_1 _20674_ (.A1(\alu_shl[11] ),
    .A2(_04993_),
    .B1(_14134_),
    .B2(_04987_),
    .X(_05000_));
 sky130_fd_sc_hd__inv_2 _20675_ (.A(_12719_),
    .Y(_02348_));
 sky130_fd_sc_hd__buf_1 _20676_ (.A(_04964_),
    .X(_05001_));
 sky130_fd_sc_hd__o32a_1 _20677_ (.A1(_02348_),
    .A2(_04117_),
    .A3(_04989_),
    .B1(_14133_),
    .B2(_05001_),
    .X(_05002_));
 sky130_vsdinv _20678_ (.A(_05002_),
    .Y(_05003_));
 sky130_fd_sc_hd__a211o_1 _20679_ (.A1(\alu_shr[11] ),
    .A2(_04992_),
    .B1(_05000_),
    .C1(_05003_),
    .X(_02145_));
 sky130_fd_sc_hd__buf_1 _20680_ (.A(_04934_),
    .X(_05004_));
 sky130_fd_sc_hd__a22o_1 _20681_ (.A1(\alu_shl[12] ),
    .A2(_04993_),
    .B1(_14127_),
    .B2(_05004_),
    .X(_05005_));
 sky130_fd_sc_hd__inv_2 _20682_ (.A(net341),
    .Y(_02351_));
 sky130_fd_sc_hd__clkbuf_2 _20683_ (.A(_04936_),
    .X(_05006_));
 sky130_fd_sc_hd__clkbuf_2 _20684_ (.A(_05006_),
    .X(_05007_));
 sky130_fd_sc_hd__o32a_1 _20685_ (.A1(_02351_),
    .A2(_04125_),
    .A3(_05007_),
    .B1(_14126_),
    .B2(_05001_),
    .X(_05008_));
 sky130_vsdinv _20686_ (.A(_05008_),
    .Y(_05009_));
 sky130_fd_sc_hd__a211o_1 _20687_ (.A1(\alu_shr[12] ),
    .A2(_04992_),
    .B1(_05005_),
    .C1(_05009_),
    .X(_02146_));
 sky130_fd_sc_hd__clkbuf_2 _20688_ (.A(_04953_),
    .X(_05010_));
 sky130_fd_sc_hd__clkbuf_2 _20689_ (.A(_04974_),
    .X(_05011_));
 sky130_fd_sc_hd__a22o_1 _20690_ (.A1(\alu_shl[13] ),
    .A2(_05011_),
    .B1(_14129_),
    .B2(_05004_),
    .X(_05012_));
 sky130_fd_sc_hd__inv_2 _20691_ (.A(_12715_),
    .Y(_02354_));
 sky130_fd_sc_hd__o32a_1 _20692_ (.A1(_02354_),
    .A2(_04130_),
    .A3(_05007_),
    .B1(_14128_),
    .B2(_05001_),
    .X(_05013_));
 sky130_vsdinv _20693_ (.A(_05013_),
    .Y(_05014_));
 sky130_fd_sc_hd__a211o_1 _20694_ (.A1(\alu_shr[13] ),
    .A2(_05010_),
    .B1(_05012_),
    .C1(_05014_),
    .X(_02147_));
 sky130_fd_sc_hd__a22o_1 _20695_ (.A1(\alu_shl[14] ),
    .A2(_05011_),
    .B1(_14131_),
    .B2(_05004_),
    .X(_05015_));
 sky130_fd_sc_hd__inv_2 _20696_ (.A(_12714_),
    .Y(_02357_));
 sky130_fd_sc_hd__o32a_1 _20697_ (.A1(_02357_),
    .A2(_04136_),
    .A3(_05007_),
    .B1(_14130_),
    .B2(_05001_),
    .X(_05016_));
 sky130_vsdinv _20698_ (.A(_05016_),
    .Y(_05017_));
 sky130_fd_sc_hd__a211o_1 _20699_ (.A1(\alu_shr[14] ),
    .A2(_05010_),
    .B1(_05015_),
    .C1(_05017_),
    .X(_02148_));
 sky130_fd_sc_hd__a22o_1 _20700_ (.A1(\alu_shl[15] ),
    .A2(_05011_),
    .B1(_14125_),
    .B2(_05004_),
    .X(_05018_));
 sky130_fd_sc_hd__inv_2 _20701_ (.A(_12710_),
    .Y(_02360_));
 sky130_fd_sc_hd__clkbuf_2 _20702_ (.A(_04939_),
    .X(_05019_));
 sky130_fd_sc_hd__clkbuf_2 _20703_ (.A(_05019_),
    .X(_05020_));
 sky130_fd_sc_hd__o32a_1 _20704_ (.A1(_02360_),
    .A2(_04140_),
    .A3(_05007_),
    .B1(_14124_),
    .B2(_05020_),
    .X(_05021_));
 sky130_vsdinv _20705_ (.A(_05021_),
    .Y(_05022_));
 sky130_fd_sc_hd__a211o_1 _20706_ (.A1(\alu_shr[15] ),
    .A2(_05010_),
    .B1(_05018_),
    .C1(_05022_),
    .X(_02149_));
 sky130_fd_sc_hd__buf_2 _20707_ (.A(_04933_),
    .X(_05023_));
 sky130_fd_sc_hd__buf_1 _20708_ (.A(_05023_),
    .X(_05024_));
 sky130_fd_sc_hd__a22o_1 _20709_ (.A1(\alu_shl[16] ),
    .A2(_05011_),
    .B1(_14081_),
    .B2(_05024_),
    .X(_05025_));
 sky130_fd_sc_hd__inv_2 _20710_ (.A(net345),
    .Y(_02363_));
 sky130_fd_sc_hd__buf_1 _20711_ (.A(_05006_),
    .X(_05026_));
 sky130_fd_sc_hd__o32a_1 _20712_ (.A1(_02363_),
    .A2(_04142_),
    .A3(_05026_),
    .B1(_14080_),
    .B2(_05020_),
    .X(_05027_));
 sky130_vsdinv _20713_ (.A(_05027_),
    .Y(_05028_));
 sky130_fd_sc_hd__a211o_1 _20714_ (.A1(\alu_shr[16] ),
    .A2(_05010_),
    .B1(_05025_),
    .C1(_05028_),
    .X(_02150_));
 sky130_fd_sc_hd__buf_1 _20715_ (.A(_04945_),
    .X(_05029_));
 sky130_fd_sc_hd__buf_1 _20716_ (.A(_04974_),
    .X(_05030_));
 sky130_fd_sc_hd__a22o_1 _20717_ (.A1(\alu_shl[17] ),
    .A2(_05030_),
    .B1(_14085_),
    .B2(_05024_),
    .X(_05031_));
 sky130_fd_sc_hd__inv_2 _20718_ (.A(_12706_),
    .Y(_02366_));
 sky130_fd_sc_hd__o32a_1 _20719_ (.A1(_02366_),
    .A2(_04157_),
    .A3(_05026_),
    .B1(_14084_),
    .B2(_05020_),
    .X(_05032_));
 sky130_vsdinv _20720_ (.A(_05032_),
    .Y(_05033_));
 sky130_fd_sc_hd__a211o_1 _20721_ (.A1(\alu_shr[17] ),
    .A2(_05029_),
    .B1(_05031_),
    .C1(_05033_),
    .X(_02151_));
 sky130_fd_sc_hd__a22o_1 _20722_ (.A1(\alu_shl[18] ),
    .A2(_05030_),
    .B1(_14083_),
    .B2(_05024_),
    .X(_05034_));
 sky130_fd_sc_hd__inv_2 _20723_ (.A(_12705_),
    .Y(_02369_));
 sky130_fd_sc_hd__o32a_1 _20724_ (.A1(_02369_),
    .A2(_04155_),
    .A3(_05026_),
    .B1(_14082_),
    .B2(_05020_),
    .X(_05035_));
 sky130_vsdinv _20725_ (.A(_05035_),
    .Y(_05036_));
 sky130_fd_sc_hd__a211o_1 _20726_ (.A1(\alu_shr[18] ),
    .A2(_05029_),
    .B1(_05034_),
    .C1(_05036_),
    .X(_02152_));
 sky130_fd_sc_hd__a22o_1 _20727_ (.A1(\alu_shl[19] ),
    .A2(_05030_),
    .B1(_14087_),
    .B2(_05024_),
    .X(_05037_));
 sky130_fd_sc_hd__inv_2 _20728_ (.A(net348),
    .Y(_02372_));
 sky130_fd_sc_hd__clkbuf_2 _20729_ (.A(_05019_),
    .X(_05038_));
 sky130_fd_sc_hd__o32a_1 _20730_ (.A1(_02372_),
    .A2(_04163_),
    .A3(_05026_),
    .B1(_14086_),
    .B2(_05038_),
    .X(_05039_));
 sky130_vsdinv _20731_ (.A(_05039_),
    .Y(_05040_));
 sky130_fd_sc_hd__a211o_1 _20732_ (.A1(\alu_shr[19] ),
    .A2(_05029_),
    .B1(_05037_),
    .C1(_05040_),
    .X(_02153_));
 sky130_fd_sc_hd__buf_1 _20733_ (.A(_05023_),
    .X(_05041_));
 sky130_fd_sc_hd__a22o_1 _20734_ (.A1(\alu_shl[20] ),
    .A2(_05030_),
    .B1(_14078_),
    .B2(_05041_),
    .X(_05042_));
 sky130_fd_sc_hd__inv_2 _20735_ (.A(_12701_),
    .Y(_02375_));
 sky130_fd_sc_hd__buf_1 _20736_ (.A(_05006_),
    .X(_05043_));
 sky130_fd_sc_hd__o32a_1 _20737_ (.A1(_02375_),
    .A2(_04168_),
    .A3(_05043_),
    .B1(_14077_),
    .B2(_05038_),
    .X(_05044_));
 sky130_vsdinv _20738_ (.A(_05044_),
    .Y(_05045_));
 sky130_fd_sc_hd__a211o_1 _20739_ (.A1(\alu_shr[20] ),
    .A2(_05029_),
    .B1(_05042_),
    .C1(_05045_),
    .X(_02154_));
 sky130_fd_sc_hd__buf_1 _20740_ (.A(_04945_),
    .X(_05046_));
 sky130_fd_sc_hd__buf_1 _20741_ (.A(_04942_),
    .X(_05047_));
 sky130_fd_sc_hd__a22o_1 _20742_ (.A1(\alu_shl[21] ),
    .A2(_05047_),
    .B1(_14074_),
    .B2(_05041_),
    .X(_05048_));
 sky130_fd_sc_hd__inv_2 _20743_ (.A(_12700_),
    .Y(_02378_));
 sky130_fd_sc_hd__o32a_1 _20744_ (.A1(_02378_),
    .A2(_04175_),
    .A3(_05043_),
    .B1(_14073_),
    .B2(_05038_),
    .X(_05049_));
 sky130_vsdinv _20745_ (.A(_05049_),
    .Y(_05050_));
 sky130_fd_sc_hd__a211o_1 _20746_ (.A1(\alu_shr[21] ),
    .A2(_05046_),
    .B1(_05048_),
    .C1(_05050_),
    .X(_02155_));
 sky130_fd_sc_hd__a22o_1 _20747_ (.A1(\alu_shl[22] ),
    .A2(_05047_),
    .B1(_14076_),
    .B2(_05041_),
    .X(_05051_));
 sky130_fd_sc_hd__inv_2 _20748_ (.A(_12699_),
    .Y(_02381_));
 sky130_fd_sc_hd__o32a_1 _20749_ (.A1(_02381_),
    .A2(_04180_),
    .A3(_05043_),
    .B1(_14075_),
    .B2(_05038_),
    .X(_05052_));
 sky130_vsdinv _20750_ (.A(_05052_),
    .Y(_05053_));
 sky130_fd_sc_hd__a211o_1 _20751_ (.A1(\alu_shr[22] ),
    .A2(_05046_),
    .B1(_05051_),
    .C1(_05053_),
    .X(_02156_));
 sky130_fd_sc_hd__a22o_1 _20752_ (.A1(\alu_shl[23] ),
    .A2(_05047_),
    .B1(_14072_),
    .B2(_05041_),
    .X(_05054_));
 sky130_fd_sc_hd__inv_2 _20753_ (.A(_12697_),
    .Y(_02384_));
 sky130_fd_sc_hd__buf_1 _20754_ (.A(_05019_),
    .X(_05055_));
 sky130_fd_sc_hd__o32a_1 _20755_ (.A1(_02384_),
    .A2(_04186_),
    .A3(_05043_),
    .B1(_14071_),
    .B2(_05055_),
    .X(_05056_));
 sky130_vsdinv _20756_ (.A(_05056_),
    .Y(_05057_));
 sky130_fd_sc_hd__a211o_1 _20757_ (.A1(\alu_shr[23] ),
    .A2(_05046_),
    .B1(_05054_),
    .C1(_05057_),
    .X(_02157_));
 sky130_fd_sc_hd__buf_1 _20758_ (.A(_05023_),
    .X(_05058_));
 sky130_fd_sc_hd__a22o_1 _20759_ (.A1(\alu_shl[24] ),
    .A2(_05047_),
    .B1(_14105_),
    .B2(_05058_),
    .X(_05059_));
 sky130_fd_sc_hd__inv_2 _20760_ (.A(net354),
    .Y(_02387_));
 sky130_fd_sc_hd__buf_1 _20761_ (.A(_05006_),
    .X(_05060_));
 sky130_fd_sc_hd__o32a_1 _20762_ (.A1(_02387_),
    .A2(_04192_),
    .A3(_05060_),
    .B1(_14104_),
    .B2(_05055_),
    .X(_05061_));
 sky130_vsdinv _20763_ (.A(_05061_),
    .Y(_05062_));
 sky130_fd_sc_hd__a211o_1 _20764_ (.A1(\alu_shr[24] ),
    .A2(_05046_),
    .B1(_05059_),
    .C1(_05062_),
    .X(_02158_));
 sky130_fd_sc_hd__buf_1 _20765_ (.A(_04945_),
    .X(_05063_));
 sky130_fd_sc_hd__buf_1 _20766_ (.A(_04942_),
    .X(_05064_));
 sky130_fd_sc_hd__a22o_1 _20767_ (.A1(\alu_shl[25] ),
    .A2(_05064_),
    .B1(_14103_),
    .B2(_05058_),
    .X(_05065_));
 sky130_fd_sc_hd__inv_2 _20768_ (.A(net355),
    .Y(_02390_));
 sky130_fd_sc_hd__o32a_1 _20769_ (.A1(_02390_),
    .A2(_04202_),
    .A3(_05060_),
    .B1(_14102_),
    .B2(_05055_),
    .X(_05066_));
 sky130_vsdinv _20770_ (.A(_05066_),
    .Y(_05067_));
 sky130_fd_sc_hd__a211o_1 _20771_ (.A1(\alu_shr[25] ),
    .A2(_05063_),
    .B1(_05065_),
    .C1(_05067_),
    .X(_02159_));
 sky130_fd_sc_hd__a22o_1 _20772_ (.A1(\alu_shl[26] ),
    .A2(_05064_),
    .B1(_14101_),
    .B2(_05058_),
    .X(_05068_));
 sky130_fd_sc_hd__inv_2 _20773_ (.A(net356),
    .Y(_02393_));
 sky130_fd_sc_hd__o32a_1 _20774_ (.A1(_02393_),
    .A2(_04206_),
    .A3(_05060_),
    .B1(_14100_),
    .B2(_05055_),
    .X(_05069_));
 sky130_vsdinv _20775_ (.A(_05069_),
    .Y(_05070_));
 sky130_fd_sc_hd__a211o_1 _20776_ (.A1(\alu_shr[26] ),
    .A2(_05063_),
    .B1(_05068_),
    .C1(_05070_),
    .X(_02160_));
 sky130_fd_sc_hd__a22o_1 _20777_ (.A1(\alu_shl[27] ),
    .A2(_05064_),
    .B1(_14099_),
    .B2(_05058_),
    .X(_05071_));
 sky130_fd_sc_hd__inv_2 _20778_ (.A(net357),
    .Y(_02396_));
 sky130_fd_sc_hd__clkbuf_2 _20779_ (.A(_05019_),
    .X(_05072_));
 sky130_fd_sc_hd__o32a_1 _20780_ (.A1(_02396_),
    .A2(_04214_),
    .A3(_05060_),
    .B1(_14098_),
    .B2(_05072_),
    .X(_05073_));
 sky130_vsdinv _20781_ (.A(_05073_),
    .Y(_05074_));
 sky130_fd_sc_hd__a211o_1 _20782_ (.A1(\alu_shr[27] ),
    .A2(_05063_),
    .B1(_05071_),
    .C1(_05074_),
    .X(_02161_));
 sky130_fd_sc_hd__buf_1 _20783_ (.A(_05023_),
    .X(_05075_));
 sky130_fd_sc_hd__a22o_1 _20784_ (.A1(\alu_shl[28] ),
    .A2(_05064_),
    .B1(_14092_),
    .B2(_05075_),
    .X(_05076_));
 sky130_fd_sc_hd__inv_2 _20785_ (.A(net358),
    .Y(_02399_));
 sky130_fd_sc_hd__clkbuf_2 _20786_ (.A(_04936_),
    .X(_05077_));
 sky130_fd_sc_hd__o32a_1 _20787_ (.A1(_02399_),
    .A2(_04223_),
    .A3(_05077_),
    .B1(_14091_),
    .B2(_05072_),
    .X(_05078_));
 sky130_vsdinv _20788_ (.A(_05078_),
    .Y(_05079_));
 sky130_fd_sc_hd__a211o_1 _20789_ (.A1(\alu_shr[28] ),
    .A2(_05063_),
    .B1(_05076_),
    .C1(_05079_),
    .X(_02162_));
 sky130_fd_sc_hd__a22o_1 _20790_ (.A1(\alu_shl[29] ),
    .A2(_04955_),
    .B1(_14090_),
    .B2(_05075_),
    .X(_05080_));
 sky130_fd_sc_hd__inv_2 _20791_ (.A(net359),
    .Y(_02402_));
 sky130_fd_sc_hd__o32a_1 _20792_ (.A1(_02402_),
    .A2(_04230_),
    .A3(_05077_),
    .B1(_14089_),
    .B2(_05072_),
    .X(_05081_));
 sky130_vsdinv _20793_ (.A(_05081_),
    .Y(_05082_));
 sky130_fd_sc_hd__a211o_1 _20794_ (.A1(\alu_shr[29] ),
    .A2(_04946_),
    .B1(_05080_),
    .C1(_05082_),
    .X(_02163_));
 sky130_fd_sc_hd__a22o_1 _20795_ (.A1(\alu_shl[30] ),
    .A2(_04955_),
    .B1(_14096_),
    .B2(_05075_),
    .X(_05083_));
 sky130_vsdinv _20796_ (.A(_12686_),
    .Y(_05084_));
 sky130_fd_sc_hd__buf_1 _20797_ (.A(_05084_),
    .X(_02405_));
 sky130_fd_sc_hd__o32a_1 _20798_ (.A1(_02405_),
    .A2(_04233_),
    .A3(_05077_),
    .B1(_14095_),
    .B2(_05072_),
    .X(_05085_));
 sky130_vsdinv _20799_ (.A(_05085_),
    .Y(_05086_));
 sky130_fd_sc_hd__a211o_1 _20800_ (.A1(\alu_shr[30] ),
    .A2(_04946_),
    .B1(_05083_),
    .C1(_05086_),
    .X(_02164_));
 sky130_fd_sc_hd__a22o_1 _20801_ (.A1(\alu_shl[31] ),
    .A2(_04955_),
    .B1(_14094_),
    .B2(_05075_),
    .X(_05087_));
 sky130_fd_sc_hd__o32a_1 _20802_ (.A1(_11683_),
    .A2(_11713_),
    .A3(_05077_),
    .B1(_14093_),
    .B2(_04964_),
    .X(_05088_));
 sky130_vsdinv _20803_ (.A(_05088_),
    .Y(_05089_));
 sky130_fd_sc_hd__a211o_1 _20804_ (.A1(\alu_shr[31] ),
    .A2(_04946_),
    .B1(_05087_),
    .C1(_05089_),
    .X(_02165_));
 sky130_fd_sc_hd__and3_1 _20805_ (.A(_11597_),
    .B(_12012_),
    .C(_00289_),
    .X(_02166_));
 sky130_vsdinv _20806_ (.A(_04417_),
    .Y(net234));
 sky130_vsdinv _20807_ (.A(_04420_),
    .Y(net235));
 sky130_vsdinv _20808_ (.A(_04422_),
    .Y(net236));
 sky130_fd_sc_hd__buf_1 _20809_ (.A(\mem_wordsize[1] ),
    .X(_05090_));
 sky130_fd_sc_hd__buf_1 _20810_ (.A(_04560_),
    .X(_05091_));
 sky130_fd_sc_hd__a22o_1 _20811_ (.A1(_12745_),
    .A2(_05090_),
    .B1(_12725_),
    .B2(_05091_),
    .X(_02167_));
 sky130_fd_sc_hd__a22o_1 _20812_ (.A1(_12743_),
    .A2(_05090_),
    .B1(_12724_),
    .B2(_05091_),
    .X(_02168_));
 sky130_fd_sc_hd__a22o_1 _20813_ (.A1(_12740_),
    .A2(_05090_),
    .B1(_12722_),
    .B2(_05091_),
    .X(_02169_));
 sky130_fd_sc_hd__a22o_1 _20814_ (.A1(_12737_),
    .A2(_05090_),
    .B1(_12720_),
    .B2(_05091_),
    .X(_02170_));
 sky130_fd_sc_hd__buf_1 _20815_ (.A(\mem_wordsize[1] ),
    .X(_05092_));
 sky130_fd_sc_hd__buf_1 _20816_ (.A(_04560_),
    .X(_05093_));
 sky130_fd_sc_hd__a22o_1 _20817_ (.A1(_12734_),
    .A2(_05092_),
    .B1(_12717_),
    .B2(_05093_),
    .X(_02171_));
 sky130_fd_sc_hd__a22o_1 _20818_ (.A1(_12732_),
    .A2(_05092_),
    .B1(_12716_),
    .B2(_05093_),
    .X(_02172_));
 sky130_fd_sc_hd__a22o_1 _20819_ (.A1(_12731_),
    .A2(_05092_),
    .B1(_12714_),
    .B2(_05093_),
    .X(_02173_));
 sky130_fd_sc_hd__a22o_1 _20820_ (.A1(_12727_),
    .A2(_05092_),
    .B1(_12711_),
    .B2(_05093_),
    .X(_02174_));
 sky130_fd_sc_hd__nor2_1 _20821_ (.A(_04949_),
    .B(net421),
    .Y(_02175_));
 sky130_fd_sc_hd__clkbuf_2 _20822_ (.A(_13966_),
    .X(_02318_));
 sky130_fd_sc_hd__nor2_1 _20823_ (.A(_02318_),
    .B(net420),
    .Y(_02176_));
 sky130_fd_sc_hd__nor2_1 _20824_ (.A(_02321_),
    .B(net420),
    .Y(_02177_));
 sky130_fd_sc_hd__buf_1 _20825_ (.A(_04412_),
    .X(_05094_));
 sky130_fd_sc_hd__nor2_1 _20826_ (.A(_02324_),
    .B(_05094_),
    .Y(_02178_));
 sky130_fd_sc_hd__nor2_1 _20827_ (.A(_02327_),
    .B(_05094_),
    .Y(_02179_));
 sky130_fd_sc_hd__nor2_1 _20828_ (.A(_02330_),
    .B(_05094_),
    .Y(_02180_));
 sky130_fd_sc_hd__nor2_1 _20829_ (.A(_02333_),
    .B(_05094_),
    .Y(_02181_));
 sky130_fd_sc_hd__nor2_1 _20830_ (.A(_02336_),
    .B(_04412_),
    .Y(_02182_));
 sky130_fd_sc_hd__or2_4 _20831_ (.A(_12558_),
    .B(_12559_),
    .X(_02183_));
 sky130_fd_sc_hd__or2_1 _20832_ (.A(\irq_pending[3] ),
    .B(net26),
    .X(_02214_));
 sky130_fd_sc_hd__and2_1 _20833_ (.A(_11873_),
    .B(_02214_),
    .X(_02215_));
 sky130_fd_sc_hd__or2_1 _20834_ (.A(\irq_pending[4] ),
    .B(net27),
    .X(_02218_));
 sky130_fd_sc_hd__and2_1 _20835_ (.A(_11872_),
    .B(_02218_),
    .X(_02219_));
 sky130_fd_sc_hd__or2_1 _20836_ (.A(_12346_),
    .B(net28),
    .X(_02221_));
 sky130_fd_sc_hd__and2_1 _20837_ (.A(\irq_mask[5] ),
    .B(_02221_),
    .X(_02222_));
 sky130_fd_sc_hd__or2_1 _20838_ (.A(\irq_pending[6] ),
    .B(net29),
    .X(_02224_));
 sky130_fd_sc_hd__and2_1 _20839_ (.A(_11870_),
    .B(_02224_),
    .X(_02225_));
 sky130_fd_sc_hd__or2_1 _20840_ (.A(_12342_),
    .B(net30),
    .X(_02227_));
 sky130_fd_sc_hd__and2_1 _20841_ (.A(\irq_mask[7] ),
    .B(_02227_),
    .X(_02228_));
 sky130_fd_sc_hd__or2_1 _20842_ (.A(\irq_pending[8] ),
    .B(net31),
    .X(_02230_));
 sky130_fd_sc_hd__and2_1 _20843_ (.A(_11866_),
    .B(_02230_),
    .X(_02231_));
 sky130_fd_sc_hd__or2_1 _20844_ (.A(_12336_),
    .B(net32),
    .X(_02233_));
 sky130_fd_sc_hd__and2_1 _20845_ (.A(\irq_mask[9] ),
    .B(_02233_),
    .X(_02234_));
 sky130_fd_sc_hd__or2_1 _20846_ (.A(\irq_pending[10] ),
    .B(net2),
    .X(_02236_));
 sky130_fd_sc_hd__and2_1 _20847_ (.A(_11864_),
    .B(_02236_),
    .X(_02237_));
 sky130_fd_sc_hd__or2_1 _20848_ (.A(_12332_),
    .B(net3),
    .X(_02239_));
 sky130_fd_sc_hd__and2_1 _20849_ (.A(\irq_mask[11] ),
    .B(_02239_),
    .X(_02240_));
 sky130_fd_sc_hd__or2_1 _20850_ (.A(\irq_pending[12] ),
    .B(net4),
    .X(_02242_));
 sky130_fd_sc_hd__and2_1 _20851_ (.A(_11861_),
    .B(_02242_),
    .X(_02243_));
 sky130_fd_sc_hd__or2_1 _20852_ (.A(_12326_),
    .B(net5),
    .X(_02245_));
 sky130_fd_sc_hd__and2_1 _20853_ (.A(\irq_mask[13] ),
    .B(_02245_),
    .X(_02246_));
 sky130_fd_sc_hd__or2_1 _20854_ (.A(\irq_pending[14] ),
    .B(net6),
    .X(_02248_));
 sky130_fd_sc_hd__and2_1 _20855_ (.A(_11858_),
    .B(_02248_),
    .X(_02249_));
 sky130_fd_sc_hd__or2_1 _20856_ (.A(_12322_),
    .B(net7),
    .X(_02251_));
 sky130_fd_sc_hd__and2_1 _20857_ (.A(\irq_mask[15] ),
    .B(_02251_),
    .X(_02252_));
 sky130_fd_sc_hd__or2_1 _20858_ (.A(\irq_pending[16] ),
    .B(net8),
    .X(_02254_));
 sky130_fd_sc_hd__and2_1 _20859_ (.A(_11853_),
    .B(_02254_),
    .X(_02255_));
 sky130_fd_sc_hd__or2_1 _20860_ (.A(\irq_pending[17] ),
    .B(net9),
    .X(_02257_));
 sky130_fd_sc_hd__and2_1 _20861_ (.A(_11852_),
    .B(_02257_),
    .X(_02258_));
 sky130_fd_sc_hd__or2_1 _20862_ (.A(_12313_),
    .B(net10),
    .X(_02260_));
 sky130_fd_sc_hd__and2_1 _20863_ (.A(\irq_mask[18] ),
    .B(_02260_),
    .X(_02261_));
 sky130_fd_sc_hd__or2_1 _20864_ (.A(\irq_pending[19] ),
    .B(net11),
    .X(_02263_));
 sky130_fd_sc_hd__and2_1 _20865_ (.A(_11846_),
    .B(_02263_),
    .X(_02264_));
 sky130_fd_sc_hd__or2_1 _20866_ (.A(_12306_),
    .B(net467),
    .X(_02266_));
 sky130_fd_sc_hd__and2_1 _20867_ (.A(\irq_mask[20] ),
    .B(_02266_),
    .X(_02267_));
 sky130_fd_sc_hd__or2_1 _20868_ (.A(\irq_pending[21] ),
    .B(net14),
    .X(_02269_));
 sky130_fd_sc_hd__and2_1 _20869_ (.A(_11845_),
    .B(_02269_),
    .X(_02270_));
 sky130_fd_sc_hd__or2_1 _20870_ (.A(_12301_),
    .B(net15),
    .X(_02272_));
 sky130_fd_sc_hd__and2_1 _20871_ (.A(\irq_mask[22] ),
    .B(_02272_),
    .X(_02273_));
 sky130_fd_sc_hd__or2_1 _20872_ (.A(\irq_pending[23] ),
    .B(net16),
    .X(_02275_));
 sky130_fd_sc_hd__and2_1 _20873_ (.A(_11839_),
    .B(_02275_),
    .X(_02276_));
 sky130_fd_sc_hd__or2_1 _20874_ (.A(_12293_),
    .B(net17),
    .X(_02278_));
 sky130_fd_sc_hd__and2_1 _20875_ (.A(\irq_mask[24] ),
    .B(_02278_),
    .X(_02279_));
 sky130_fd_sc_hd__or2_1 _20876_ (.A(\irq_pending[25] ),
    .B(net18),
    .X(_02281_));
 sky130_fd_sc_hd__and2_1 _20877_ (.A(_11838_),
    .B(_02281_),
    .X(_02282_));
 sky130_fd_sc_hd__or2_1 _20878_ (.A(_12290_),
    .B(net19),
    .X(_02284_));
 sky130_fd_sc_hd__and2_1 _20879_ (.A(\irq_mask[26] ),
    .B(_02284_),
    .X(_02285_));
 sky130_fd_sc_hd__or2_1 _20880_ (.A(\irq_pending[27] ),
    .B(net466),
    .X(_02287_));
 sky130_fd_sc_hd__and2_1 _20881_ (.A(_11834_),
    .B(_02287_),
    .X(_02288_));
 sky130_fd_sc_hd__or2_1 _20882_ (.A(_12284_),
    .B(net465),
    .X(_02290_));
 sky130_fd_sc_hd__and2_1 _20883_ (.A(\irq_mask[28] ),
    .B(_02290_),
    .X(_02291_));
 sky130_fd_sc_hd__or2_1 _20884_ (.A(\irq_pending[29] ),
    .B(net22),
    .X(_02293_));
 sky130_fd_sc_hd__and2_1 _20885_ (.A(_11833_),
    .B(_02293_),
    .X(_02294_));
 sky130_fd_sc_hd__or2_1 _20886_ (.A(_12279_),
    .B(net24),
    .X(_02296_));
 sky130_fd_sc_hd__and2_1 _20887_ (.A(\irq_mask[30] ),
    .B(_02296_),
    .X(_02297_));
 sky130_fd_sc_hd__or2_1 _20888_ (.A(\irq_pending[31] ),
    .B(net25),
    .X(_02299_));
 sky130_fd_sc_hd__and2_1 _20889_ (.A(_11814_),
    .B(_02299_),
    .X(_02300_));
 sky130_fd_sc_hd__or4_4 _20890_ (.A(\timer[3] ),
    .B(\timer[2] ),
    .C(\timer[7] ),
    .D(\timer[6] ),
    .X(_05095_));
 sky130_fd_sc_hd__or4_4 _20891_ (.A(\timer[19] ),
    .B(\timer[18] ),
    .C(\timer[15] ),
    .D(\timer[14] ),
    .X(_05096_));
 sky130_fd_sc_hd__or4_4 _20892_ (.A(\timer[21] ),
    .B(\timer[20] ),
    .C(\timer[23] ),
    .D(\timer[22] ),
    .X(_05097_));
 sky130_fd_sc_hd__or4_4 _20893_ (.A(\timer[31] ),
    .B(\timer[30] ),
    .C(\timer[27] ),
    .D(\timer[26] ),
    .X(_05098_));
 sky130_fd_sc_hd__or4_4 _20894_ (.A(_05095_),
    .B(_05096_),
    .C(_05097_),
    .D(_05098_),
    .X(_05099_));
 sky130_fd_sc_hd__or4_4 _20895_ (.A(\timer[9] ),
    .B(\timer[8] ),
    .C(\timer[11] ),
    .D(\timer[10] ),
    .X(_05100_));
 sky130_fd_sc_hd__or4_4 _20896_ (.A(\timer[5] ),
    .B(_14202_),
    .C(\timer[29] ),
    .D(\timer[28] ),
    .X(_05101_));
 sky130_fd_sc_hd__or4_4 _20897_ (.A(\timer[25] ),
    .B(\timer[24] ),
    .C(\timer[1] ),
    .D(_14201_),
    .X(_05102_));
 sky130_fd_sc_hd__or4_4 _20898_ (.A(\timer[13] ),
    .B(\timer[12] ),
    .C(\timer[17] ),
    .D(\timer[16] ),
    .X(_05103_));
 sky130_fd_sc_hd__or4_4 _20899_ (.A(_05100_),
    .B(_05101_),
    .C(_05102_),
    .D(_05103_),
    .X(_05104_));
 sky130_fd_sc_hd__o21ai_1 _20900_ (.A1(_05099_),
    .A2(_05104_),
    .B1(_11621_),
    .Y(_02302_));
 sky130_fd_sc_hd__or2_1 _20901_ (.A(_02303_),
    .B(net1),
    .X(_02304_));
 sky130_fd_sc_hd__and2_1 _20902_ (.A(\irq_mask[0] ),
    .B(_02304_),
    .X(_02305_));
 sky130_fd_sc_hd__nor2_2 _20903_ (.A(_12355_),
    .B(net23),
    .Y(_02307_));
 sky130_fd_sc_hd__or2_1 _20904_ (.A(_12354_),
    .B(_02307_),
    .X(_02308_));
 sky130_fd_sc_hd__nor2_1 _20905_ (.A(_11827_),
    .B(_02310_),
    .Y(_02311_));
 sky130_fd_sc_hd__or2_1 _20906_ (.A(_14021_),
    .B(_02311_),
    .X(_02312_));
 sky130_fd_sc_hd__or2_1 _20907_ (.A(_02313_),
    .B(_14021_),
    .X(_02314_));
 sky130_fd_sc_hd__or2_1 _20908_ (.A(_02316_),
    .B(_14021_),
    .X(_02317_));
 sky130_fd_sc_hd__o32a_1 _20909_ (.A1(_02387_),
    .A2(net322),
    .A3(_14103_),
    .B1(_02390_),
    .B2(_04201_),
    .X(_05105_));
 sky130_fd_sc_hd__o22a_1 _20910_ (.A1(_02393_),
    .A2(_13410_),
    .B1(_14101_),
    .B2(_05105_),
    .X(_05106_));
 sky130_fd_sc_hd__o22a_1 _20911_ (.A1(_02396_),
    .A2(_04213_),
    .B1(_14099_),
    .B2(_05106_),
    .X(_05107_));
 sky130_fd_sc_hd__o22a_1 _20912_ (.A1(_02399_),
    .A2(_13403_),
    .B1(_14092_),
    .B2(_05107_),
    .X(_05108_));
 sky130_fd_sc_hd__o22a_1 _20913_ (.A1(_02402_),
    .A2(_13400_),
    .B1(_14090_),
    .B2(_05108_),
    .X(_05109_));
 sky130_fd_sc_hd__or2_1 _20914_ (.A(_14097_),
    .B(_05109_),
    .X(_05110_));
 sky130_fd_sc_hd__o32a_1 _20915_ (.A1(_02363_),
    .A2(_13437_),
    .A3(_14085_),
    .B1(_02366_),
    .B2(_13435_),
    .X(_05111_));
 sky130_fd_sc_hd__o22a_1 _20916_ (.A1(_02369_),
    .A2(_13433_),
    .B1(_14083_),
    .B2(_05111_),
    .X(_05112_));
 sky130_fd_sc_hd__o22a_1 _20917_ (.A1(_02372_),
    .A2(_13430_),
    .B1(_14087_),
    .B2(_05112_),
    .X(_05113_));
 sky130_fd_sc_hd__o22a_1 _20918_ (.A1(_02375_),
    .A2(_13427_),
    .B1(_14078_),
    .B2(_05113_),
    .X(_05114_));
 sky130_fd_sc_hd__o22a_1 _20919_ (.A1(_02378_),
    .A2(_13425_),
    .B1(_14074_),
    .B2(_05114_),
    .X(_05115_));
 sky130_fd_sc_hd__o22a_1 _20920_ (.A1(_02381_),
    .A2(_13423_),
    .B1(_14076_),
    .B2(_05115_),
    .X(_05116_));
 sky130_fd_sc_hd__o32a_1 _20921_ (.A1(_02351_),
    .A2(_13450_),
    .A3(_14129_),
    .B1(_02354_),
    .B2(_13448_),
    .X(_05117_));
 sky130_fd_sc_hd__o22a_1 _20922_ (.A1(_02357_),
    .A2(_13446_),
    .B1(_14131_),
    .B2(_05117_),
    .X(_05118_));
 sky130_fd_sc_hd__o21a_1 _20923_ (.A1(_13966_),
    .A2(_00048_),
    .B1(_13484_),
    .X(_05119_));
 sky130_fd_sc_hd__o32a_1 _20924_ (.A1(_00049_),
    .A2(_14122_),
    .A3(_05119_),
    .B1(_13962_),
    .B2(_13482_),
    .X(_05120_));
 sky130_fd_sc_hd__o22a_1 _20925_ (.A1(_13957_),
    .A2(_13478_),
    .B1(_14115_),
    .B2(_05120_),
    .X(_05121_));
 sky130_fd_sc_hd__o22a_1 _20926_ (.A1(_13952_),
    .A2(_13474_),
    .B1(_14118_),
    .B2(_05121_),
    .X(_05122_));
 sky130_fd_sc_hd__o22a_1 _20927_ (.A1(_02330_),
    .A2(_13471_),
    .B1(_14109_),
    .B2(_05122_),
    .X(_05123_));
 sky130_fd_sc_hd__o22a_1 _20928_ (.A1(_04980_),
    .A2(_13468_),
    .B1(_14120_),
    .B2(_05123_),
    .X(_05124_));
 sky130_fd_sc_hd__o22a_1 _20929_ (.A1(_02336_),
    .A2(_13465_),
    .B1(_14111_),
    .B2(_05124_),
    .X(_05125_));
 sky130_fd_sc_hd__o32a_1 _20930_ (.A1(_02339_),
    .A2(_13460_),
    .A3(_14138_),
    .B1(_02342_),
    .B2(_13458_),
    .X(_05126_));
 sky130_fd_sc_hd__o22a_1 _20931_ (.A1(_02345_),
    .A2(_13456_),
    .B1(_14140_),
    .B2(_05126_),
    .X(_05127_));
 sky130_fd_sc_hd__or2_1 _20932_ (.A(_14134_),
    .B(_05127_),
    .X(_05128_));
 sky130_fd_sc_hd__o221a_1 _20933_ (.A1(_02348_),
    .A2(_13453_),
    .B1(_14141_),
    .B2(_05125_),
    .C1(_05128_),
    .X(_05129_));
 sky130_fd_sc_hd__or2_2 _20934_ (.A(_14132_),
    .B(_05129_),
    .X(_05130_));
 sky130_fd_sc_hd__o221ai_2 _20935_ (.A1(_02360_),
    .A2(_13442_),
    .B1(_14125_),
    .B2(_05118_),
    .C1(_05130_),
    .Y(_05131_));
 sky130_fd_sc_hd__or3b_4 _20936_ (.A(_14079_),
    .B(_14088_),
    .C_N(_05131_),
    .X(_05132_));
 sky130_fd_sc_hd__o221a_1 _20937_ (.A1(_02384_),
    .A2(_13420_),
    .B1(_14072_),
    .B2(_05116_),
    .C1(_05132_),
    .X(_05133_));
 sky130_fd_sc_hd__or2_1 _20938_ (.A(_14107_),
    .B(_05133_),
    .X(_05134_));
 sky130_fd_sc_hd__o311a_1 _20939_ (.A1(_05084_),
    .A2(_13398_),
    .A3(_14094_),
    .B1(_05110_),
    .C1(_05134_),
    .X(_05135_));
 sky130_fd_sc_hd__o21a_1 _20940_ (.A1(_11682_),
    .A2(_11714_),
    .B1(_05135_),
    .X(_05136_));
 sky130_fd_sc_hd__nor2_1 _20941_ (.A(_00000_),
    .B(_05136_),
    .Y(_00002_));
 sky130_vsdinv _20942_ (.A(_05135_),
    .Y(_05137_));
 sky130_fd_sc_hd__o221a_2 _20943_ (.A1(_14094_),
    .A2(_05137_),
    .B1(_13394_),
    .B2(_11714_),
    .C1(_14143_),
    .X(_00001_));
 sky130_vsdinv _20944_ (.A(\pcpi_mul.rs2[0] ),
    .Y(_05138_));
 sky130_fd_sc_hd__buf_1 _20945_ (.A(_05138_),
    .X(_05139_));
 sky130_fd_sc_hd__buf_1 _20946_ (.A(_05139_),
    .X(_05140_));
 sky130_fd_sc_hd__buf_2 _20947_ (.A(_05140_),
    .X(_05141_));
 sky130_fd_sc_hd__buf_1 _20948_ (.A(_05141_),
    .X(_05142_));
 sky130_fd_sc_hd__clkbuf_4 _20949_ (.A(_05142_),
    .X(_05143_));
 sky130_fd_sc_hd__clkbuf_4 _20950_ (.A(_05143_),
    .X(_05144_));
 sky130_vsdinv _20951_ (.A(\pcpi_mul.rs1[0] ),
    .Y(_05145_));
 sky130_fd_sc_hd__buf_1 _20952_ (.A(_05145_),
    .X(_05146_));
 sky130_fd_sc_hd__clkbuf_2 _20953_ (.A(_05146_),
    .X(_05147_));
 sky130_fd_sc_hd__clkbuf_2 _20954_ (.A(_05147_),
    .X(_05148_));
 sky130_fd_sc_hd__buf_2 _20955_ (.A(_05148_),
    .X(_05149_));
 sky130_fd_sc_hd__clkbuf_2 _20956_ (.A(_05149_),
    .X(_05150_));
 sky130_fd_sc_hd__buf_1 _20957_ (.A(_05150_),
    .X(_05151_));
 sky130_fd_sc_hd__clkbuf_2 _20958_ (.A(_05151_),
    .X(_05152_));
 sky130_fd_sc_hd__buf_1 _20959_ (.A(_05152_),
    .X(_05153_));
 sky130_fd_sc_hd__buf_1 _20960_ (.A(_05153_),
    .X(_05154_));
 sky130_fd_sc_hd__nor2_1 _20961_ (.A(_05144_),
    .B(_05154_),
    .Y(_02623_));
 sky130_fd_sc_hd__or2_1 _20962_ (.A(net211),
    .B(net200),
    .X(_05155_));
 sky130_fd_sc_hd__o21ai_1 _20963_ (.A1(_02318_),
    .A2(_04949_),
    .B1(_05155_),
    .Y(_02319_));
 sky130_vsdinv _20964_ (.A(_02320_),
    .Y(_05156_));
 sky130_fd_sc_hd__o22a_1 _20965_ (.A1(_14256_),
    .A2(_05156_),
    .B1(_13484_),
    .B2(_02320_),
    .X(_05157_));
 sky130_vsdinv _20966_ (.A(_05157_),
    .Y(_05158_));
 sky130_fd_sc_hd__o32a_1 _20967_ (.A1(_04949_),
    .A2(_13488_),
    .A3(_05157_),
    .B1(_14070_),
    .B2(_05158_),
    .X(_02602_));
 sky130_fd_sc_hd__or2_1 _20968_ (.A(net222),
    .B(_05155_),
    .X(_05159_));
 sky130_fd_sc_hd__a21bo_1 _20969_ (.A1(_12741_),
    .A2(_05155_),
    .B1_N(_05159_),
    .X(_02322_));
 sky130_fd_sc_hd__o22a_1 _20970_ (.A1(_04413_),
    .A2(_05156_),
    .B1(_14070_),
    .B2(_05158_),
    .X(_05160_));
 sky130_fd_sc_hd__nor2_1 _20971_ (.A(_13481_),
    .B(_02323_),
    .Y(_05161_));
 sky130_fd_sc_hd__a21o_1 _20972_ (.A1(_13483_),
    .A2(_02323_),
    .B1(_05161_),
    .X(_05162_));
 sky130_fd_sc_hd__o2bb2a_1 _20973_ (.A1_N(_05160_),
    .A2_N(_05162_),
    .B1(_05160_),
    .B2(_05162_),
    .X(_02613_));
 sky130_fd_sc_hd__or2_1 _20974_ (.A(net225),
    .B(_05159_),
    .X(_05163_));
 sky130_vsdinv _20975_ (.A(_05163_),
    .Y(_05164_));
 sky130_fd_sc_hd__a21o_1 _20976_ (.A1(_12738_),
    .A2(_05159_),
    .B1(_05164_),
    .X(_02325_));
 sky130_fd_sc_hd__o2bb2a_1 _20977_ (.A1_N(_13481_),
    .A2_N(_02323_),
    .B1(_05160_),
    .B2(_05161_),
    .X(_05165_));
 sky130_fd_sc_hd__nor2_1 _20978_ (.A(_13477_),
    .B(_02326_),
    .Y(_05166_));
 sky130_fd_sc_hd__a21o_1 _20979_ (.A1(_13479_),
    .A2(_02326_),
    .B1(_05166_),
    .X(_05167_));
 sky130_fd_sc_hd__o2bb2a_1 _20980_ (.A1_N(_05165_),
    .A2_N(_05167_),
    .B1(_05165_),
    .B2(_05167_),
    .X(_02616_));
 sky130_fd_sc_hd__or2_1 _20981_ (.A(net226),
    .B(_05163_),
    .X(_05168_));
 sky130_fd_sc_hd__o21ai_1 _20982_ (.A1(_02327_),
    .A2(_05164_),
    .B1(_05168_),
    .Y(_02328_));
 sky130_fd_sc_hd__o2bb2a_1 _20983_ (.A1_N(_13477_),
    .A2_N(_02326_),
    .B1(_05165_),
    .B2(_05166_),
    .X(_05169_));
 sky130_fd_sc_hd__nor2_1 _20984_ (.A(_13473_),
    .B(_02329_),
    .Y(_05170_));
 sky130_fd_sc_hd__a21o_1 _20985_ (.A1(_13475_),
    .A2(_02329_),
    .B1(_05170_),
    .X(_05171_));
 sky130_fd_sc_hd__o2bb2a_1 _20986_ (.A1_N(_05169_),
    .A2_N(_05171_),
    .B1(_05169_),
    .B2(_05171_),
    .X(_02617_));
 sky130_fd_sc_hd__or2_1 _20987_ (.A(net227),
    .B(_05168_),
    .X(_05172_));
 sky130_vsdinv _20988_ (.A(_05172_),
    .Y(_05173_));
 sky130_fd_sc_hd__a21o_1 _20989_ (.A1(_12733_),
    .A2(_05168_),
    .B1(_05173_),
    .X(_02331_));
 sky130_fd_sc_hd__o2bb2a_1 _20990_ (.A1_N(_13473_),
    .A2_N(_02329_),
    .B1(_05169_),
    .B2(_05170_),
    .X(_05174_));
 sky130_fd_sc_hd__nor2_1 _20991_ (.A(_13470_),
    .B(_02332_),
    .Y(_05175_));
 sky130_fd_sc_hd__a21o_1 _20992_ (.A1(_13472_),
    .A2(_02332_),
    .B1(_05175_),
    .X(_05176_));
 sky130_fd_sc_hd__o2bb2a_1 _20993_ (.A1_N(_05174_),
    .A2_N(_05176_),
    .B1(_05174_),
    .B2(_05176_),
    .X(_02618_));
 sky130_fd_sc_hd__or2_1 _20994_ (.A(net228),
    .B(_05172_),
    .X(_05177_));
 sky130_fd_sc_hd__o21ai_1 _20995_ (.A1(_02333_),
    .A2(_05173_),
    .B1(_05177_),
    .Y(_02334_));
 sky130_fd_sc_hd__o2bb2ai_2 _20996_ (.A1_N(_13470_),
    .A2_N(_02332_),
    .B1(_05174_),
    .B2(_05175_),
    .Y(_05178_));
 sky130_fd_sc_hd__o2bb2a_1 _20997_ (.A1_N(_13467_),
    .A2_N(_02335_),
    .B1(_13467_),
    .B2(_02335_),
    .X(_05179_));
 sky130_fd_sc_hd__o2bb2a_1 _20998_ (.A1_N(_05178_),
    .A2_N(_05179_),
    .B1(_05178_),
    .B2(_05179_),
    .X(_02619_));
 sky130_fd_sc_hd__or2_1 _20999_ (.A(net229),
    .B(_05177_),
    .X(_05180_));
 sky130_vsdinv _21000_ (.A(_05180_),
    .Y(_05181_));
 sky130_fd_sc_hd__a21o_1 _21001_ (.A1(_12728_),
    .A2(_05177_),
    .B1(_05181_),
    .X(_02337_));
 sky130_fd_sc_hd__o2bb2a_1 _21002_ (.A1_N(_13464_),
    .A2_N(_02338_),
    .B1(_13463_),
    .B2(_02338_),
    .X(_05182_));
 sky130_fd_sc_hd__a22o_1 _21003_ (.A1(_13469_),
    .A2(_02335_),
    .B1(_05178_),
    .B2(_05179_),
    .X(_05183_));
 sky130_fd_sc_hd__a2bb2oi_1 _21004_ (.A1_N(_05182_),
    .A2_N(_05183_),
    .B1(_05182_),
    .B2(_05183_),
    .Y(_02620_));
 sky130_fd_sc_hd__or2_1 _21005_ (.A(net368),
    .B(_05180_),
    .X(_05184_));
 sky130_fd_sc_hd__o21ai_1 _21006_ (.A1(_02339_),
    .A2(_05181_),
    .B1(_05184_),
    .Y(_02340_));
 sky130_fd_sc_hd__or2_1 _21007_ (.A(_13463_),
    .B(_02338_),
    .X(_05185_));
 sky130_fd_sc_hd__a32o_1 _21008_ (.A1(_13467_),
    .A2(_02335_),
    .A3(_05185_),
    .B1(_13464_),
    .B2(_02338_),
    .X(_05186_));
 sky130_fd_sc_hd__a31o_1 _21009_ (.A1(_05179_),
    .A2(_05182_),
    .A3(_05178_),
    .B1(_05186_),
    .X(_05187_));
 sky130_fd_sc_hd__o2bb2a_2 _21010_ (.A1_N(_13459_),
    .A2_N(_02341_),
    .B1(_13459_),
    .B2(_02341_),
    .X(_05188_));
 sky130_fd_sc_hd__o2bb2a_1 _21011_ (.A1_N(_05187_),
    .A2_N(_05188_),
    .B1(_05187_),
    .B2(_05188_),
    .X(_02621_));
 sky130_fd_sc_hd__or2_1 _21012_ (.A(net369),
    .B(_05184_),
    .X(_05189_));
 sky130_vsdinv _21013_ (.A(_05189_),
    .Y(_05190_));
 sky130_fd_sc_hd__a21o_1 _21014_ (.A1(_12724_),
    .A2(_05184_),
    .B1(_05190_),
    .X(_02343_));
 sky130_fd_sc_hd__o2bb2a_2 _21015_ (.A1_N(_13457_),
    .A2_N(_02344_),
    .B1(_04097_),
    .B2(_02344_),
    .X(_05191_));
 sky130_fd_sc_hd__a22o_1 _21016_ (.A1(_13461_),
    .A2(_02341_),
    .B1(_05187_),
    .B2(_05188_),
    .X(_05192_));
 sky130_fd_sc_hd__a2bb2oi_1 _21017_ (.A1_N(_05191_),
    .A2_N(_05192_),
    .B1(_05191_),
    .B2(_05192_),
    .Y(_02622_));
 sky130_fd_sc_hd__or2_1 _21018_ (.A(net339),
    .B(_05189_),
    .X(_05193_));
 sky130_fd_sc_hd__o21ai_1 _21019_ (.A1(_02345_),
    .A2(_05190_),
    .B1(_05193_),
    .Y(_02346_));
 sky130_vsdinv _21020_ (.A(_02347_),
    .Y(_05194_));
 sky130_fd_sc_hd__a22o_1 _21021_ (.A1(_13455_),
    .A2(_02347_),
    .B1(_04112_),
    .B2(_05194_),
    .X(_05195_));
 sky130_fd_sc_hd__or2_1 _21022_ (.A(net337),
    .B(_02344_),
    .X(_05196_));
 sky130_fd_sc_hd__a32o_1 _21023_ (.A1(_13460_),
    .A2(_02341_),
    .A3(_05196_),
    .B1(_13457_),
    .B2(_02344_),
    .X(_05197_));
 sky130_fd_sc_hd__a31oi_4 _21024_ (.A1(_05188_),
    .A2(_05191_),
    .A3(_05187_),
    .B1(_05197_),
    .Y(_05198_));
 sky130_fd_sc_hd__a2bb2oi_1 _21025_ (.A1_N(_05195_),
    .A2_N(_05198_),
    .B1(_05195_),
    .B2(_05198_),
    .Y(_02592_));
 sky130_fd_sc_hd__or2_1 _21026_ (.A(net340),
    .B(_05193_),
    .X(_05199_));
 sky130_vsdinv _21027_ (.A(_05199_),
    .Y(_05200_));
 sky130_fd_sc_hd__a21o_1 _21028_ (.A1(_12720_),
    .A2(_05193_),
    .B1(_05200_),
    .X(_02349_));
 sky130_vsdinv _21029_ (.A(_02350_),
    .Y(_05201_));
 sky130_fd_sc_hd__a22o_1 _21030_ (.A1(_13452_),
    .A2(_02350_),
    .B1(_04117_),
    .B2(_05201_),
    .X(_05202_));
 sky130_fd_sc_hd__o22a_1 _21031_ (.A1(_04112_),
    .A2(_05194_),
    .B1(_05195_),
    .B2(_05198_),
    .X(_05203_));
 sky130_fd_sc_hd__a2bb2oi_1 _21032_ (.A1_N(_05202_),
    .A2_N(_05203_),
    .B1(_05202_),
    .B2(_05203_),
    .Y(_02593_));
 sky130_fd_sc_hd__or2_1 _21033_ (.A(net341),
    .B(_05199_),
    .X(_05204_));
 sky130_fd_sc_hd__o21ai_1 _21034_ (.A1(_02351_),
    .A2(_05200_),
    .B1(_05204_),
    .Y(_02352_));
 sky130_vsdinv _21035_ (.A(_02353_),
    .Y(_05205_));
 sky130_fd_sc_hd__a22o_1 _21036_ (.A1(_13449_),
    .A2(_02353_),
    .B1(_04125_),
    .B2(_05205_),
    .X(_05206_));
 sky130_fd_sc_hd__o22a_1 _21037_ (.A1(_04117_),
    .A2(_05201_),
    .B1(_05202_),
    .B2(_05203_),
    .X(_05207_));
 sky130_fd_sc_hd__a2bb2oi_1 _21038_ (.A1_N(_05206_),
    .A2_N(_05207_),
    .B1(_05206_),
    .B2(_05207_),
    .Y(_02594_));
 sky130_fd_sc_hd__or2_1 _21039_ (.A(net342),
    .B(_05204_),
    .X(_05208_));
 sky130_vsdinv _21040_ (.A(_05208_),
    .Y(_05209_));
 sky130_fd_sc_hd__a21o_1 _21041_ (.A1(_12716_),
    .A2(_05204_),
    .B1(_05209_),
    .X(_02355_));
 sky130_vsdinv _21042_ (.A(_02356_),
    .Y(_05210_));
 sky130_fd_sc_hd__a22o_1 _21043_ (.A1(_13447_),
    .A2(_02356_),
    .B1(_04130_),
    .B2(_05210_),
    .X(_05211_));
 sky130_fd_sc_hd__o22a_1 _21044_ (.A1(_04125_),
    .A2(_05205_),
    .B1(_05206_),
    .B2(_05207_),
    .X(_05212_));
 sky130_fd_sc_hd__a2bb2oi_1 _21045_ (.A1_N(_05211_),
    .A2_N(_05212_),
    .B1(_05211_),
    .B2(_05212_),
    .Y(_02595_));
 sky130_fd_sc_hd__or2_1 _21046_ (.A(net343),
    .B(_05208_),
    .X(_05213_));
 sky130_fd_sc_hd__o21ai_1 _21047_ (.A1(_02357_),
    .A2(_05209_),
    .B1(_05213_),
    .Y(_02358_));
 sky130_vsdinv _21048_ (.A(_02359_),
    .Y(_05214_));
 sky130_fd_sc_hd__a22o_1 _21049_ (.A1(_13445_),
    .A2(_02359_),
    .B1(_04136_),
    .B2(_05214_),
    .X(_05215_));
 sky130_fd_sc_hd__o22a_1 _21050_ (.A1(_04130_),
    .A2(_05210_),
    .B1(_05211_),
    .B2(_05212_),
    .X(_05216_));
 sky130_fd_sc_hd__a2bb2oi_1 _21051_ (.A1_N(_05215_),
    .A2_N(_05216_),
    .B1(_05215_),
    .B2(_05216_),
    .Y(_02596_));
 sky130_fd_sc_hd__or2_1 _21052_ (.A(net344),
    .B(_05213_),
    .X(_05217_));
 sky130_vsdinv _21053_ (.A(_05217_),
    .Y(_05218_));
 sky130_fd_sc_hd__a21o_1 _21054_ (.A1(_12711_),
    .A2(_05213_),
    .B1(_05218_),
    .X(_02361_));
 sky130_vsdinv _21055_ (.A(_02362_),
    .Y(_05219_));
 sky130_fd_sc_hd__a22o_1 _21056_ (.A1(_13441_),
    .A2(_02362_),
    .B1(_04140_),
    .B2(_05219_),
    .X(_05220_));
 sky130_fd_sc_hd__o22a_2 _21057_ (.A1(_04136_),
    .A2(_05214_),
    .B1(_05215_),
    .B2(_05216_),
    .X(_05221_));
 sky130_fd_sc_hd__a2bb2oi_1 _21058_ (.A1_N(_05220_),
    .A2_N(_05221_),
    .B1(_05220_),
    .B2(_05221_),
    .Y(_02597_));
 sky130_fd_sc_hd__or2_1 _21059_ (.A(net345),
    .B(_05217_),
    .X(_05222_));
 sky130_fd_sc_hd__o21ai_1 _21060_ (.A1(_02363_),
    .A2(_05218_),
    .B1(_05222_),
    .Y(_02364_));
 sky130_fd_sc_hd__o22ai_4 _21061_ (.A1(_04140_),
    .A2(_05219_),
    .B1(_05220_),
    .B2(_05221_),
    .Y(_05223_));
 sky130_fd_sc_hd__o2bb2a_2 _21062_ (.A1_N(_13436_),
    .A2_N(_02365_),
    .B1(_13436_),
    .B2(_02365_),
    .X(_05224_));
 sky130_fd_sc_hd__o2bb2a_1 _21063_ (.A1_N(_05223_),
    .A2_N(_05224_),
    .B1(_05223_),
    .B2(_05224_),
    .X(_02598_));
 sky130_fd_sc_hd__or2_1 _21064_ (.A(net346),
    .B(_05222_),
    .X(_05225_));
 sky130_vsdinv _21065_ (.A(_05225_),
    .Y(_05226_));
 sky130_fd_sc_hd__a21o_1 _21066_ (.A1(_12706_),
    .A2(_05222_),
    .B1(_05226_),
    .X(_02367_));
 sky130_fd_sc_hd__o2bb2a_2 _21067_ (.A1_N(_04149_),
    .A2_N(_02368_),
    .B1(_04149_),
    .B2(_02368_),
    .X(_05227_));
 sky130_fd_sc_hd__a22o_1 _21068_ (.A1(_13438_),
    .A2(_02365_),
    .B1(_05223_),
    .B2(_05224_),
    .X(_05228_));
 sky130_fd_sc_hd__a2bb2oi_1 _21069_ (.A1_N(_05227_),
    .A2_N(_05228_),
    .B1(_05227_),
    .B2(_05228_),
    .Y(_02599_));
 sky130_fd_sc_hd__or2_1 _21070_ (.A(net347),
    .B(_05225_),
    .X(_05229_));
 sky130_fd_sc_hd__o21ai_1 _21071_ (.A1(_02369_),
    .A2(_05226_),
    .B1(_05229_),
    .Y(_02370_));
 sky130_vsdinv _21072_ (.A(_02371_),
    .Y(_05230_));
 sky130_fd_sc_hd__a22o_1 _21073_ (.A1(_13432_),
    .A2(_02371_),
    .B1(_04154_),
    .B2(_05230_),
    .X(_05231_));
 sky130_fd_sc_hd__or2_1 _21074_ (.A(net314),
    .B(_02368_),
    .X(_05232_));
 sky130_fd_sc_hd__a32o_1 _21075_ (.A1(_13437_),
    .A2(_02365_),
    .A3(_05232_),
    .B1(_13434_),
    .B2(_02368_),
    .X(_05233_));
 sky130_fd_sc_hd__a31oi_4 _21076_ (.A1(_05224_),
    .A2(_05227_),
    .A3(_05223_),
    .B1(_05233_),
    .Y(_05234_));
 sky130_fd_sc_hd__a2bb2oi_1 _21077_ (.A1_N(_05231_),
    .A2_N(_05234_),
    .B1(_05231_),
    .B2(_05234_),
    .Y(_02600_));
 sky130_fd_sc_hd__or2_1 _21078_ (.A(net348),
    .B(_05229_),
    .X(_05235_));
 sky130_vsdinv _21079_ (.A(_05235_),
    .Y(_05236_));
 sky130_fd_sc_hd__a21o_1 _21080_ (.A1(_12703_),
    .A2(_05229_),
    .B1(_05236_),
    .X(_02373_));
 sky130_vsdinv _21081_ (.A(_02374_),
    .Y(_05237_));
 sky130_fd_sc_hd__a22o_1 _21082_ (.A1(_13429_),
    .A2(_02374_),
    .B1(_04162_),
    .B2(_05237_),
    .X(_05238_));
 sky130_fd_sc_hd__o22a_1 _21083_ (.A1(_04155_),
    .A2(_05230_),
    .B1(_05231_),
    .B2(_05234_),
    .X(_05239_));
 sky130_fd_sc_hd__a2bb2oi_1 _21084_ (.A1_N(_05238_),
    .A2_N(_05239_),
    .B1(_05238_),
    .B2(_05239_),
    .Y(_02601_));
 sky130_fd_sc_hd__or2_1 _21085_ (.A(net350),
    .B(_05235_),
    .X(_05240_));
 sky130_fd_sc_hd__o21ai_1 _21086_ (.A1(_02375_),
    .A2(_05236_),
    .B1(_05240_),
    .Y(_02376_));
 sky130_vsdinv _21087_ (.A(_02377_),
    .Y(_05241_));
 sky130_fd_sc_hd__a22o_1 _21088_ (.A1(_13426_),
    .A2(_02377_),
    .B1(_04167_),
    .B2(_05241_),
    .X(_05242_));
 sky130_fd_sc_hd__o22a_1 _21089_ (.A1(_04163_),
    .A2(_05237_),
    .B1(_05238_),
    .B2(_05239_),
    .X(_05243_));
 sky130_fd_sc_hd__a2bb2oi_1 _21090_ (.A1_N(_05242_),
    .A2_N(_05243_),
    .B1(_05242_),
    .B2(_05243_),
    .Y(_02603_));
 sky130_fd_sc_hd__or2_1 _21091_ (.A(net351),
    .B(_05240_),
    .X(_05244_));
 sky130_vsdinv _21092_ (.A(_05244_),
    .Y(_05245_));
 sky130_fd_sc_hd__a21o_1 _21093_ (.A1(_12700_),
    .A2(_05240_),
    .B1(_05245_),
    .X(_02379_));
 sky130_vsdinv _21094_ (.A(_02380_),
    .Y(_05246_));
 sky130_fd_sc_hd__a22o_1 _21095_ (.A1(_13424_),
    .A2(_02380_),
    .B1(_04174_),
    .B2(_05246_),
    .X(_05247_));
 sky130_fd_sc_hd__o22a_1 _21096_ (.A1(_04168_),
    .A2(_05241_),
    .B1(_05242_),
    .B2(_05243_),
    .X(_05248_));
 sky130_fd_sc_hd__a2bb2oi_1 _21097_ (.A1_N(_05247_),
    .A2_N(_05248_),
    .B1(_05247_),
    .B2(_05248_),
    .Y(_02604_));
 sky130_fd_sc_hd__or2_1 _21098_ (.A(net352),
    .B(_05244_),
    .X(_05249_));
 sky130_fd_sc_hd__o21ai_1 _21099_ (.A1(_02381_),
    .A2(_05245_),
    .B1(_05249_),
    .Y(_02382_));
 sky130_vsdinv _21100_ (.A(_02383_),
    .Y(_05250_));
 sky130_fd_sc_hd__a22o_1 _21101_ (.A1(_13422_),
    .A2(_02383_),
    .B1(_04179_),
    .B2(_05250_),
    .X(_05251_));
 sky130_fd_sc_hd__o22a_1 _21102_ (.A1(_04175_),
    .A2(_05246_),
    .B1(_05247_),
    .B2(_05248_),
    .X(_05252_));
 sky130_fd_sc_hd__a2bb2oi_1 _21103_ (.A1_N(_05251_),
    .A2_N(_05252_),
    .B1(_05251_),
    .B2(_05252_),
    .Y(_02605_));
 sky130_fd_sc_hd__or2_1 _21104_ (.A(net353),
    .B(_05249_),
    .X(_05253_));
 sky130_vsdinv _21105_ (.A(_05253_),
    .Y(_05254_));
 sky130_fd_sc_hd__a21o_1 _21106_ (.A1(_12697_),
    .A2(_05249_),
    .B1(_05254_),
    .X(_02385_));
 sky130_vsdinv _21107_ (.A(_02386_),
    .Y(_05255_));
 sky130_fd_sc_hd__a22o_1 _21108_ (.A1(_13419_),
    .A2(_02386_),
    .B1(_04185_),
    .B2(_05255_),
    .X(_05256_));
 sky130_fd_sc_hd__o22a_2 _21109_ (.A1(_04180_),
    .A2(_05250_),
    .B1(_05251_),
    .B2(_05252_),
    .X(_05257_));
 sky130_fd_sc_hd__a2bb2oi_1 _21110_ (.A1_N(_05256_),
    .A2_N(_05257_),
    .B1(_05256_),
    .B2(_05257_),
    .Y(_02606_));
 sky130_fd_sc_hd__or2_1 _21111_ (.A(net354),
    .B(_05253_),
    .X(_05258_));
 sky130_fd_sc_hd__o21ai_1 _21112_ (.A1(_02387_),
    .A2(_05254_),
    .B1(_05258_),
    .Y(_02388_));
 sky130_fd_sc_hd__o22ai_4 _21113_ (.A1(_04186_),
    .A2(_05255_),
    .B1(_05256_),
    .B2(_05257_),
    .Y(_05259_));
 sky130_fd_sc_hd__o2bb2a_1 _21114_ (.A1_N(_13415_),
    .A2_N(_02389_),
    .B1(_13415_),
    .B2(_02389_),
    .X(_05260_));
 sky130_fd_sc_hd__o2bb2a_1 _21115_ (.A1_N(_05259_),
    .A2_N(_05260_),
    .B1(_05259_),
    .B2(_05260_),
    .X(_02607_));
 sky130_fd_sc_hd__or2_1 _21116_ (.A(_12694_),
    .B(_05258_),
    .X(_05261_));
 sky130_vsdinv _21117_ (.A(_05261_),
    .Y(_05262_));
 sky130_fd_sc_hd__a21o_1 _21118_ (.A1(_12694_),
    .A2(_05258_),
    .B1(_05262_),
    .X(_02391_));
 sky130_fd_sc_hd__o2bb2a_1 _21119_ (.A1_N(_04201_),
    .A2_N(_02392_),
    .B1(_04201_),
    .B2(_02392_),
    .X(_05263_));
 sky130_fd_sc_hd__a22o_1 _21120_ (.A1(_13417_),
    .A2(_02389_),
    .B1(_05259_),
    .B2(_05260_),
    .X(_05264_));
 sky130_fd_sc_hd__a2bb2oi_1 _21121_ (.A1_N(_05263_),
    .A2_N(_05264_),
    .B1(_05263_),
    .B2(_05264_),
    .Y(_02608_));
 sky130_fd_sc_hd__or2_1 _21122_ (.A(_12693_),
    .B(_05261_),
    .X(_05265_));
 sky130_fd_sc_hd__o21ai_1 _21123_ (.A1(_02393_),
    .A2(_05262_),
    .B1(_05265_),
    .Y(_02394_));
 sky130_fd_sc_hd__or2_1 _21124_ (.A(_13413_),
    .B(_02392_),
    .X(_05266_));
 sky130_fd_sc_hd__a32o_1 _21125_ (.A1(_13416_),
    .A2(_02389_),
    .A3(_05266_),
    .B1(_13414_),
    .B2(_02392_),
    .X(_05267_));
 sky130_fd_sc_hd__a31o_1 _21126_ (.A1(_05260_),
    .A2(_05263_),
    .A3(_05259_),
    .B1(_05267_),
    .X(_05268_));
 sky130_fd_sc_hd__o2bb2a_1 _21127_ (.A1_N(_13411_),
    .A2_N(_02395_),
    .B1(_13410_),
    .B2(_02395_),
    .X(_05269_));
 sky130_fd_sc_hd__o2bb2a_1 _21128_ (.A1_N(_05268_),
    .A2_N(_05269_),
    .B1(_05268_),
    .B2(_05269_),
    .X(_02609_));
 sky130_fd_sc_hd__or2_1 _21129_ (.A(_12691_),
    .B(_05265_),
    .X(_05270_));
 sky130_vsdinv _21130_ (.A(_05270_),
    .Y(_05271_));
 sky130_fd_sc_hd__a21o_1 _21131_ (.A1(_12691_),
    .A2(_05265_),
    .B1(_05271_),
    .X(_02397_));
 sky130_fd_sc_hd__o2bb2a_1 _21132_ (.A1_N(_04213_),
    .A2_N(_02398_),
    .B1(_04213_),
    .B2(_02398_),
    .X(_05272_));
 sky130_fd_sc_hd__a22o_1 _21133_ (.A1(_13412_),
    .A2(_02395_),
    .B1(_05268_),
    .B2(_05269_),
    .X(_05273_));
 sky130_fd_sc_hd__a2bb2oi_1 _21134_ (.A1_N(_05272_),
    .A2_N(_05273_),
    .B1(_05272_),
    .B2(_05273_),
    .Y(_02610_));
 sky130_fd_sc_hd__or2_1 _21135_ (.A(_12688_),
    .B(_05270_),
    .X(_05274_));
 sky130_fd_sc_hd__o21ai_1 _21136_ (.A1(_02399_),
    .A2(_05271_),
    .B1(_05274_),
    .Y(_02400_));
 sky130_fd_sc_hd__or2_1 _21137_ (.A(_13407_),
    .B(_02398_),
    .X(_05275_));
 sky130_fd_sc_hd__a32o_1 _21138_ (.A1(_13411_),
    .A2(_02395_),
    .A3(_05275_),
    .B1(_13408_),
    .B2(_02398_),
    .X(_05276_));
 sky130_fd_sc_hd__a31o_1 _21139_ (.A1(_05269_),
    .A2(_05272_),
    .A3(_05268_),
    .B1(_05276_),
    .X(_05277_));
 sky130_fd_sc_hd__nor2_1 _21140_ (.A(_13403_),
    .B(_02401_),
    .Y(_05278_));
 sky130_fd_sc_hd__a21oi_1 _21141_ (.A1(_13405_),
    .A2(_02401_),
    .B1(_05278_),
    .Y(_05279_));
 sky130_vsdinv _21142_ (.A(_05277_),
    .Y(_05280_));
 sky130_vsdinv _21143_ (.A(_05279_),
    .Y(_05281_));
 sky130_fd_sc_hd__o22a_1 _21144_ (.A1(_05277_),
    .A2(_05279_),
    .B1(_05280_),
    .B2(_05281_),
    .X(_02611_));
 sky130_fd_sc_hd__or2_1 _21145_ (.A(_12687_),
    .B(_05274_),
    .X(_05282_));
 sky130_vsdinv _21146_ (.A(_05282_),
    .Y(_05283_));
 sky130_fd_sc_hd__a21o_1 _21147_ (.A1(_12687_),
    .A2(_05274_),
    .B1(_05283_),
    .X(_02403_));
 sky130_fd_sc_hd__o2bb2a_1 _21148_ (.A1_N(_13404_),
    .A2_N(_02401_),
    .B1(_05280_),
    .B2(_05278_),
    .X(_05284_));
 sky130_fd_sc_hd__nor2_1 _21149_ (.A(_13401_),
    .B(_02404_),
    .Y(_05285_));
 sky130_fd_sc_hd__a21o_1 _21150_ (.A1(_13402_),
    .A2(_02404_),
    .B1(_05285_),
    .X(_05286_));
 sky130_fd_sc_hd__o2bb2a_1 _21151_ (.A1_N(_05284_),
    .A2_N(_05286_),
    .B1(_05284_),
    .B2(_05286_),
    .X(_02612_));
 sky130_fd_sc_hd__or2_1 _21152_ (.A(_12686_),
    .B(_05282_),
    .X(_05287_));
 sky130_fd_sc_hd__o21ai_1 _21153_ (.A1(_02405_),
    .A2(_05283_),
    .B1(_05287_),
    .Y(_02406_));
 sky130_vsdinv _21154_ (.A(_02407_),
    .Y(_05288_));
 sky130_fd_sc_hd__a22o_1 _21155_ (.A1(_13399_),
    .A2(_02407_),
    .B1(_04233_),
    .B2(_05288_),
    .X(_05289_));
 sky130_fd_sc_hd__o2bb2a_1 _21156_ (.A1_N(_13401_),
    .A2_N(_02404_),
    .B1(_05284_),
    .B2(_05285_),
    .X(_05290_));
 sky130_fd_sc_hd__a2bb2oi_1 _21157_ (.A1_N(_05289_),
    .A2_N(_05290_),
    .B1(_05289_),
    .B2(_05290_),
    .Y(_02614_));
 sky130_fd_sc_hd__a32o_1 _21158_ (.A1(_02405_),
    .A2(_05283_),
    .A3(_11712_),
    .B1(_11714_),
    .B2(_05287_),
    .X(_02408_));
 sky130_fd_sc_hd__o22ai_1 _21159_ (.A1(_04233_),
    .A2(_05288_),
    .B1(_05289_),
    .B2(_05290_),
    .Y(_05291_));
 sky130_fd_sc_hd__a2bb2o_1 _21160_ (.A1_N(_11684_),
    .A2_N(_02409_),
    .B1(_11684_),
    .B2(_02409_),
    .X(_05292_));
 sky130_fd_sc_hd__a2bb2o_1 _21161_ (.A1_N(_05291_),
    .A2_N(_05292_),
    .B1(_05291_),
    .B2(_05292_),
    .X(_02615_));
 sky130_vsdinv _21162_ (.A(\pcpi_mul.rs1[1] ),
    .Y(_05293_));
 sky130_fd_sc_hd__buf_1 _21163_ (.A(_05293_),
    .X(_05294_));
 sky130_fd_sc_hd__buf_1 _21164_ (.A(_05294_),
    .X(_05295_));
 sky130_fd_sc_hd__clkbuf_2 _21165_ (.A(_05295_),
    .X(_05296_));
 sky130_fd_sc_hd__clkbuf_2 _21166_ (.A(_05296_),
    .X(_05297_));
 sky130_fd_sc_hd__clkbuf_2 _21167_ (.A(_05297_),
    .X(_05298_));
 sky130_fd_sc_hd__buf_2 _21168_ (.A(_05298_),
    .X(_05299_));
 sky130_fd_sc_hd__buf_1 _21169_ (.A(_05299_),
    .X(_05300_));
 sky130_vsdinv _21170_ (.A(\pcpi_mul.rs2[1] ),
    .Y(_05301_));
 sky130_fd_sc_hd__buf_1 _21171_ (.A(_05301_),
    .X(_05302_));
 sky130_fd_sc_hd__buf_1 _21172_ (.A(_05302_),
    .X(_05303_));
 sky130_fd_sc_hd__clkbuf_2 _21173_ (.A(_05303_),
    .X(_05304_));
 sky130_fd_sc_hd__buf_2 _21174_ (.A(_05304_),
    .X(_05305_));
 sky130_fd_sc_hd__clkbuf_2 _21175_ (.A(_05305_),
    .X(_05306_));
 sky130_fd_sc_hd__buf_2 _21176_ (.A(_05306_),
    .X(_05307_));
 sky130_fd_sc_hd__buf_2 _21177_ (.A(_05307_),
    .X(_05308_));
 sky130_fd_sc_hd__o22a_1 _21178_ (.A1(_05144_),
    .A2(_05300_),
    .B1(_05308_),
    .B2(_05154_),
    .X(_05309_));
 sky130_fd_sc_hd__or4_4 _21179_ (.A(_05144_),
    .B(_05299_),
    .C(_05308_),
    .D(_05153_),
    .X(_05310_));
 sky130_fd_sc_hd__nor2b_1 _21180_ (.A(_05309_),
    .B_N(_05310_),
    .Y(_02624_));
 sky130_fd_sc_hd__buf_2 _21181_ (.A(_05142_),
    .X(_05311_));
 sky130_vsdinv _21182_ (.A(\pcpi_mul.rs1[2] ),
    .Y(_05312_));
 sky130_fd_sc_hd__buf_1 _21183_ (.A(_05312_),
    .X(_05313_));
 sky130_fd_sc_hd__clkbuf_2 _21184_ (.A(_05313_),
    .X(_05314_));
 sky130_fd_sc_hd__clkbuf_2 _21185_ (.A(_05314_),
    .X(_05315_));
 sky130_fd_sc_hd__clkbuf_2 _21186_ (.A(_05315_),
    .X(_05316_));
 sky130_fd_sc_hd__clkbuf_2 _21187_ (.A(_05295_),
    .X(_05317_));
 sky130_fd_sc_hd__clkbuf_2 _21188_ (.A(_05317_),
    .X(_05318_));
 sky130_fd_sc_hd__clkbuf_2 _21189_ (.A(_05318_),
    .X(_05319_));
 sky130_vsdinv _21190_ (.A(\pcpi_mul.rs2[2] ),
    .Y(_05320_));
 sky130_fd_sc_hd__buf_1 _21191_ (.A(_05320_),
    .X(_05321_));
 sky130_fd_sc_hd__clkbuf_4 _21192_ (.A(_05321_),
    .X(_05322_));
 sky130_fd_sc_hd__buf_1 _21193_ (.A(_05322_),
    .X(_05323_));
 sky130_fd_sc_hd__clkbuf_2 _21194_ (.A(_05147_),
    .X(_05324_));
 sky130_fd_sc_hd__clkbuf_2 _21195_ (.A(_05324_),
    .X(_05325_));
 sky130_fd_sc_hd__o22a_1 _21196_ (.A1(_05305_),
    .A2(_05319_),
    .B1(_05323_),
    .B2(_05325_),
    .X(_05326_));
 sky130_fd_sc_hd__or4_4 _21197_ (.A(_05304_),
    .B(_05318_),
    .C(_05322_),
    .D(_05148_),
    .X(_05327_));
 sky130_vsdinv _21198_ (.A(_05327_),
    .Y(_05328_));
 sky130_fd_sc_hd__or2_1 _21199_ (.A(_05326_),
    .B(_05328_),
    .X(_05329_));
 sky130_fd_sc_hd__or3_4 _21200_ (.A(_05311_),
    .B(_05316_),
    .C(_05329_),
    .X(_05330_));
 sky130_vsdinv _21201_ (.A(_05330_),
    .Y(_05331_));
 sky130_fd_sc_hd__o21a_1 _21202_ (.A1(_05143_),
    .A2(_05316_),
    .B1(_05329_),
    .X(_05332_));
 sky130_fd_sc_hd__or2_1 _21203_ (.A(_05331_),
    .B(_05332_),
    .X(_05333_));
 sky130_fd_sc_hd__or2_1 _21204_ (.A(_05310_),
    .B(_05333_),
    .X(_05334_));
 sky130_fd_sc_hd__a21boi_1 _21205_ (.A1(_05310_),
    .A2(_05333_),
    .B1_N(_05334_),
    .Y(_02625_));
 sky130_vsdinv _21206_ (.A(\pcpi_mul.rs1[3] ),
    .Y(_05335_));
 sky130_fd_sc_hd__buf_1 _21207_ (.A(_05335_),
    .X(_05336_));
 sky130_fd_sc_hd__buf_1 _21208_ (.A(_05336_),
    .X(_05337_));
 sky130_fd_sc_hd__clkbuf_2 _21209_ (.A(_05337_),
    .X(_05338_));
 sky130_fd_sc_hd__clkbuf_2 _21210_ (.A(_05338_),
    .X(_05339_));
 sky130_fd_sc_hd__buf_2 _21211_ (.A(_05339_),
    .X(_05340_));
 sky130_fd_sc_hd__or2_1 _21212_ (.A(_05141_),
    .B(_05340_),
    .X(_05341_));
 sky130_fd_sc_hd__buf_1 _21213_ (.A(_05313_),
    .X(_05342_));
 sky130_fd_sc_hd__clkbuf_2 _21214_ (.A(_05342_),
    .X(_05343_));
 sky130_fd_sc_hd__o22a_1 _21215_ (.A1(_05321_),
    .A2(_05317_),
    .B1(_05304_),
    .B2(_05343_),
    .X(_05344_));
 sky130_fd_sc_hd__buf_1 _21216_ (.A(_13618_),
    .X(_05345_));
 sky130_fd_sc_hd__buf_1 _21217_ (.A(_05345_),
    .X(_05346_));
 sky130_fd_sc_hd__and4_1 _21218_ (.A(_13172_),
    .B(_13623_),
    .C(_13177_),
    .D(_05346_),
    .X(_05347_));
 sky130_fd_sc_hd__nor2_1 _21219_ (.A(_05344_),
    .B(_05347_),
    .Y(_05348_));
 sky130_vsdinv _21220_ (.A(\pcpi_mul.rs2[3] ),
    .Y(_05349_));
 sky130_fd_sc_hd__buf_1 _21221_ (.A(_05349_),
    .X(_05350_));
 sky130_fd_sc_hd__buf_1 _21222_ (.A(_05350_),
    .X(_05351_));
 sky130_fd_sc_hd__nor2_1 _21223_ (.A(_05351_),
    .B(_05149_),
    .Y(_05352_));
 sky130_fd_sc_hd__a2bb2o_1 _21224_ (.A1_N(_05348_),
    .A2_N(_05352_),
    .B1(_05348_),
    .B2(_05352_),
    .X(_05353_));
 sky130_fd_sc_hd__or2_2 _21225_ (.A(_05341_),
    .B(_05353_),
    .X(_05354_));
 sky130_fd_sc_hd__a21bo_1 _21226_ (.A1(_05341_),
    .A2(_05353_),
    .B1_N(_05354_),
    .X(_05355_));
 sky130_vsdinv _21227_ (.A(_05355_),
    .Y(_05356_));
 sky130_fd_sc_hd__o22a_1 _21228_ (.A1(_05331_),
    .A2(_05356_),
    .B1(_05330_),
    .B2(_05355_),
    .X(_05357_));
 sky130_fd_sc_hd__a2bb2o_1 _21229_ (.A1_N(_05328_),
    .A2_N(_05357_),
    .B1(_05328_),
    .B2(_05356_),
    .X(_05358_));
 sky130_fd_sc_hd__or2_1 _21230_ (.A(_05334_),
    .B(_05358_),
    .X(_05359_));
 sky130_fd_sc_hd__a21boi_1 _21231_ (.A1(_05334_),
    .A2(_05358_),
    .B1_N(_05359_),
    .Y(_02626_));
 sky130_vsdinv _21232_ (.A(\pcpi_mul.rs2[4] ),
    .Y(_05360_));
 sky130_fd_sc_hd__buf_1 _21233_ (.A(_05360_),
    .X(_05361_));
 sky130_fd_sc_hd__clkbuf_2 _21234_ (.A(_05361_),
    .X(_05362_));
 sky130_fd_sc_hd__clkbuf_2 _21235_ (.A(_05146_),
    .X(_05363_));
 sky130_vsdinv _21236_ (.A(\pcpi_mul.rs1[4] ),
    .Y(_05364_));
 sky130_fd_sc_hd__buf_1 _21237_ (.A(_05364_),
    .X(_05365_));
 sky130_fd_sc_hd__buf_1 _21238_ (.A(_05365_),
    .X(_05366_));
 sky130_fd_sc_hd__o22a_1 _21239_ (.A1(_05362_),
    .A2(_05363_),
    .B1(_05140_),
    .B2(_05366_),
    .X(_05367_));
 sky130_fd_sc_hd__buf_1 _21240_ (.A(_05138_),
    .X(_05368_));
 sky130_fd_sc_hd__buf_1 _21241_ (.A(_05365_),
    .X(_05369_));
 sky130_fd_sc_hd__or4_4 _21242_ (.A(_05361_),
    .B(_05147_),
    .C(_05368_),
    .D(_05369_),
    .X(_05370_));
 sky130_fd_sc_hd__or2b_1 _21243_ (.A(_05367_),
    .B_N(_05370_),
    .X(_05371_));
 sky130_fd_sc_hd__buf_1 _21244_ (.A(_05320_),
    .X(_05372_));
 sky130_fd_sc_hd__o22a_1 _21245_ (.A1(_05372_),
    .A2(_05342_),
    .B1(_05303_),
    .B2(_05337_),
    .X(_05373_));
 sky130_fd_sc_hd__buf_1 _21246_ (.A(_13171_),
    .X(_05374_));
 sky130_fd_sc_hd__buf_1 _21247_ (.A(_13176_),
    .X(_05375_));
 sky130_fd_sc_hd__buf_1 _21248_ (.A(_13614_),
    .X(_05376_));
 sky130_fd_sc_hd__and4_1 _21249_ (.A(_05374_),
    .B(_05345_),
    .C(_05375_),
    .D(_05376_),
    .X(_05377_));
 sky130_fd_sc_hd__nor2_2 _21250_ (.A(_05373_),
    .B(_05377_),
    .Y(_05378_));
 sky130_fd_sc_hd__buf_1 _21251_ (.A(_05295_),
    .X(_05379_));
 sky130_fd_sc_hd__buf_2 _21252_ (.A(_05379_),
    .X(_05380_));
 sky130_fd_sc_hd__nor2_2 _21253_ (.A(_05350_),
    .B(_05380_),
    .Y(_05381_));
 sky130_fd_sc_hd__a2bb2o_1 _21254_ (.A1_N(_05378_),
    .A2_N(_05381_),
    .B1(_05378_),
    .B2(_05381_),
    .X(_05382_));
 sky130_fd_sc_hd__or2_1 _21255_ (.A(_05371_),
    .B(_05382_),
    .X(_05383_));
 sky130_fd_sc_hd__a21bo_1 _21256_ (.A1(_05371_),
    .A2(_05382_),
    .B1_N(_05383_),
    .X(_05384_));
 sky130_fd_sc_hd__o2bb2a_1 _21257_ (.A1_N(_05354_),
    .A2_N(_05384_),
    .B1(_05354_),
    .B2(_05384_),
    .X(_05385_));
 sky130_vsdinv _21258_ (.A(_05385_),
    .Y(_05386_));
 sky130_fd_sc_hd__a31o_1 _21259_ (.A1(\pcpi_mul.rs2[3] ),
    .A2(_13626_),
    .A3(_05348_),
    .B1(_05347_),
    .X(_05387_));
 sky130_vsdinv _21260_ (.A(_05387_),
    .Y(_05388_));
 sky130_fd_sc_hd__a22o_1 _21261_ (.A1(_05386_),
    .A2(_05388_),
    .B1(_05385_),
    .B2(_05387_),
    .X(_05389_));
 sky130_fd_sc_hd__o22a_1 _21262_ (.A1(_05330_),
    .A2(_05355_),
    .B1(_05327_),
    .B2(_05355_),
    .X(_05390_));
 sky130_fd_sc_hd__or2_1 _21263_ (.A(_05389_),
    .B(_05390_),
    .X(_05391_));
 sky130_vsdinv _21264_ (.A(_05391_),
    .Y(_05392_));
 sky130_fd_sc_hd__a21o_1 _21265_ (.A1(_05389_),
    .A2(_05390_),
    .B1(_05392_),
    .X(_05393_));
 sky130_fd_sc_hd__or2_1 _21266_ (.A(_05359_),
    .B(_05393_),
    .X(_05394_));
 sky130_vsdinv _21267_ (.A(_05394_),
    .Y(_05395_));
 sky130_fd_sc_hd__a21oi_1 _21268_ (.A1(_05359_),
    .A2(_05393_),
    .B1(_05395_),
    .Y(_02627_));
 sky130_fd_sc_hd__o22a_1 _21269_ (.A1(_05354_),
    .A2(_05384_),
    .B1(_05386_),
    .B2(_05388_),
    .X(_05396_));
 sky130_fd_sc_hd__a21oi_2 _21270_ (.A1(_05378_),
    .A2(_05381_),
    .B1(_05377_),
    .Y(_05397_));
 sky130_vsdinv _21271_ (.A(\pcpi_mul.rs1[5] ),
    .Y(_05398_));
 sky130_fd_sc_hd__buf_1 _21272_ (.A(_05398_),
    .X(_05399_));
 sky130_fd_sc_hd__or2_1 _21273_ (.A(_05139_),
    .B(_05399_),
    .X(_05400_));
 sky130_fd_sc_hd__and4_1 _21274_ (.A(_13163_),
    .B(_13622_),
    .C(_13157_),
    .D(\pcpi_mul.rs1[0] ),
    .X(_05401_));
 sky130_fd_sc_hd__buf_1 _21275_ (.A(_05360_),
    .X(_05402_));
 sky130_vsdinv _21276_ (.A(\pcpi_mul.rs2[5] ),
    .Y(_05403_));
 sky130_fd_sc_hd__buf_1 _21277_ (.A(_05403_),
    .X(_05404_));
 sky130_fd_sc_hd__o22a_1 _21278_ (.A1(_05402_),
    .A2(_05294_),
    .B1(_05404_),
    .B2(_05145_),
    .X(_05405_));
 sky130_fd_sc_hd__or2_1 _21279_ (.A(_05401_),
    .B(_05405_),
    .X(_05406_));
 sky130_fd_sc_hd__a2bb2o_1 _21280_ (.A1_N(_05400_),
    .A2_N(_05406_),
    .B1(_05400_),
    .B2(_05406_),
    .X(_05407_));
 sky130_fd_sc_hd__a2bb2o_1 _21281_ (.A1_N(_05370_),
    .A2_N(_05407_),
    .B1(_05370_),
    .B2(_05407_),
    .X(_05408_));
 sky130_fd_sc_hd__or2_1 _21282_ (.A(_05351_),
    .B(_05343_),
    .X(_05409_));
 sky130_fd_sc_hd__and4_1 _21283_ (.A(_13172_),
    .B(_05376_),
    .C(_13177_),
    .D(_13611_),
    .X(_05410_));
 sky130_fd_sc_hd__o22a_1 _21284_ (.A1(_05321_),
    .A2(_05337_),
    .B1(_05303_),
    .B2(_05369_),
    .X(_05411_));
 sky130_fd_sc_hd__or2_1 _21285_ (.A(_05410_),
    .B(_05411_),
    .X(_05412_));
 sky130_fd_sc_hd__a2bb2o_1 _21286_ (.A1_N(_05409_),
    .A2_N(_05412_),
    .B1(_05409_),
    .B2(_05412_),
    .X(_05413_));
 sky130_fd_sc_hd__a2bb2o_1 _21287_ (.A1_N(_05408_),
    .A2_N(_05413_),
    .B1(_05408_),
    .B2(_05413_),
    .X(_05414_));
 sky130_fd_sc_hd__a2bb2o_1 _21288_ (.A1_N(_05383_),
    .A2_N(_05414_),
    .B1(_05383_),
    .B2(_05414_),
    .X(_05415_));
 sky130_fd_sc_hd__a2bb2o_1 _21289_ (.A1_N(_05397_),
    .A2_N(_05415_),
    .B1(_05397_),
    .B2(_05415_),
    .X(_05416_));
 sky130_fd_sc_hd__or2_1 _21290_ (.A(_05396_),
    .B(_05416_),
    .X(_05417_));
 sky130_fd_sc_hd__a21bo_1 _21291_ (.A1(_05396_),
    .A2(_05416_),
    .B1_N(_05417_),
    .X(_05418_));
 sky130_fd_sc_hd__or2_1 _21292_ (.A(_05394_),
    .B(_05418_),
    .X(_05419_));
 sky130_vsdinv _21293_ (.A(\pcpi_mul.rs2[6] ),
    .Y(_05420_));
 sky130_fd_sc_hd__buf_4 _21294_ (.A(_05420_),
    .X(_05421_));
 sky130_fd_sc_hd__buf_1 _21295_ (.A(_05421_),
    .X(_05422_));
 sky130_fd_sc_hd__buf_2 _21296_ (.A(_05422_),
    .X(_05423_));
 sky130_fd_sc_hd__buf_1 _21297_ (.A(_05423_),
    .X(_05424_));
 sky130_fd_sc_hd__clkbuf_4 _21298_ (.A(_05424_),
    .X(_05425_));
 sky130_fd_sc_hd__or2_2 _21299_ (.A(_05425_),
    .B(_05151_),
    .X(_05426_));
 sky130_fd_sc_hd__o21ba_1 _21300_ (.A1(_05409_),
    .A2(_05412_),
    .B1_N(_05410_),
    .X(_05427_));
 sky130_fd_sc_hd__and4_1 _21301_ (.A(_13171_),
    .B(_13610_),
    .C(_13176_),
    .D(_13606_),
    .X(_05428_));
 sky130_fd_sc_hd__o22a_1 _21302_ (.A1(_05320_),
    .A2(_05364_),
    .B1(_05302_),
    .B2(_05399_),
    .X(_05429_));
 sky130_fd_sc_hd__or2_1 _21303_ (.A(_05428_),
    .B(_05429_),
    .X(_05430_));
 sky130_fd_sc_hd__or2_1 _21304_ (.A(_05349_),
    .B(_05337_),
    .X(_05431_));
 sky130_fd_sc_hd__a2bb2o_1 _21305_ (.A1_N(_05430_),
    .A2_N(_05431_),
    .B1(_05430_),
    .B2(_05431_),
    .X(_05432_));
 sky130_fd_sc_hd__and4_1 _21306_ (.A(_13157_),
    .B(_13621_),
    .C(_13163_),
    .D(_13618_),
    .X(_05433_));
 sky130_fd_sc_hd__o22a_1 _21307_ (.A1(_05403_),
    .A2(_05294_),
    .B1(_05402_),
    .B2(_05313_),
    .X(_05434_));
 sky130_fd_sc_hd__or2_1 _21308_ (.A(_05433_),
    .B(_05434_),
    .X(_05435_));
 sky130_vsdinv _21309_ (.A(\pcpi_mul.rs1[6] ),
    .Y(_05436_));
 sky130_fd_sc_hd__or2_1 _21310_ (.A(_05139_),
    .B(_05436_),
    .X(_05437_));
 sky130_fd_sc_hd__a2bb2o_1 _21311_ (.A1_N(_05435_),
    .A2_N(_05437_),
    .B1(_05435_),
    .B2(_05437_),
    .X(_05438_));
 sky130_fd_sc_hd__o21ba_1 _21312_ (.A1(_05400_),
    .A2(_05406_),
    .B1_N(_05401_),
    .X(_05439_));
 sky130_fd_sc_hd__a2bb2o_1 _21313_ (.A1_N(_05438_),
    .A2_N(_05439_),
    .B1(_05438_),
    .B2(_05439_),
    .X(_05440_));
 sky130_fd_sc_hd__a2bb2o_1 _21314_ (.A1_N(_05432_),
    .A2_N(_05440_),
    .B1(_05432_),
    .B2(_05440_),
    .X(_05441_));
 sky130_fd_sc_hd__o22a_1 _21315_ (.A1(_05370_),
    .A2(_05407_),
    .B1(_05408_),
    .B2(_05413_),
    .X(_05442_));
 sky130_fd_sc_hd__a2bb2o_1 _21316_ (.A1_N(_05441_),
    .A2_N(_05442_),
    .B1(_05441_),
    .B2(_05442_),
    .X(_05443_));
 sky130_fd_sc_hd__a2bb2o_1 _21317_ (.A1_N(_05427_),
    .A2_N(_05443_),
    .B1(_05427_),
    .B2(_05443_),
    .X(_05444_));
 sky130_fd_sc_hd__or2_1 _21318_ (.A(_05426_),
    .B(_05444_),
    .X(_05445_));
 sky130_fd_sc_hd__a21bo_1 _21319_ (.A1(_05426_),
    .A2(_05444_),
    .B1_N(_05445_),
    .X(_05446_));
 sky130_fd_sc_hd__o22a_1 _21320_ (.A1(_05383_),
    .A2(_05414_),
    .B1(_05397_),
    .B2(_05415_),
    .X(_05447_));
 sky130_fd_sc_hd__or2_2 _21321_ (.A(_05446_),
    .B(_05447_),
    .X(_05448_));
 sky130_fd_sc_hd__a21bo_1 _21322_ (.A1(_05446_),
    .A2(_05447_),
    .B1_N(_05448_),
    .X(_05449_));
 sky130_fd_sc_hd__or2_1 _21323_ (.A(_05391_),
    .B(_05418_),
    .X(_05450_));
 sky130_fd_sc_hd__nand2_1 _21324_ (.A(_05417_),
    .B(_05450_),
    .Y(_05451_));
 sky130_fd_sc_hd__a2bb2oi_2 _21325_ (.A1_N(_05449_),
    .A2_N(_05451_),
    .B1(_05449_),
    .B2(_05451_),
    .Y(_05452_));
 sky130_fd_sc_hd__a2bb2oi_1 _21326_ (.A1_N(_05419_),
    .A2_N(_05452_),
    .B1(_05419_),
    .B2(_05452_),
    .Y(_02683_));
 sky130_fd_sc_hd__o22a_1 _21327_ (.A1(_05419_),
    .A2(_05452_),
    .B1(_05449_),
    .B2(_05450_),
    .X(_05453_));
 sky130_vsdinv _21328_ (.A(\pcpi_mul.rs2[7] ),
    .Y(_05454_));
 sky130_fd_sc_hd__buf_1 _21329_ (.A(_05454_),
    .X(_05455_));
 sky130_fd_sc_hd__clkbuf_2 _21330_ (.A(_05455_),
    .X(_05456_));
 sky130_fd_sc_hd__buf_2 _21331_ (.A(_05456_),
    .X(_05457_));
 sky130_fd_sc_hd__buf_2 _21332_ (.A(_05457_),
    .X(_05458_));
 sky130_fd_sc_hd__buf_1 _21333_ (.A(_05324_),
    .X(_05459_));
 sky130_fd_sc_hd__clkbuf_4 _21334_ (.A(_05422_),
    .X(_05460_));
 sky130_fd_sc_hd__o22a_2 _21335_ (.A1(_05458_),
    .A2(_05459_),
    .B1(_05460_),
    .B2(_05298_),
    .X(_05461_));
 sky130_fd_sc_hd__or4_4 _21336_ (.A(_05455_),
    .B(_05146_),
    .C(_05420_),
    .D(_05379_),
    .X(_05462_));
 sky130_fd_sc_hd__or2b_1 _21337_ (.A(_05461_),
    .B_N(_05462_),
    .X(_05463_));
 sky130_fd_sc_hd__o21ba_1 _21338_ (.A1(_05430_),
    .A2(_05431_),
    .B1_N(_05428_),
    .X(_05464_));
 sky130_fd_sc_hd__and4_1 _21339_ (.A(_13171_),
    .B(_13606_),
    .C(_13176_),
    .D(\pcpi_mul.rs1[6] ),
    .X(_05465_));
 sky130_fd_sc_hd__o22a_1 _21340_ (.A1(_05320_),
    .A2(_05399_),
    .B1(_05301_),
    .B2(_05436_),
    .X(_05466_));
 sky130_fd_sc_hd__or2_1 _21341_ (.A(_05465_),
    .B(_05466_),
    .X(_05467_));
 sky130_fd_sc_hd__or2_1 _21342_ (.A(_05349_),
    .B(_05365_),
    .X(_05468_));
 sky130_fd_sc_hd__a2bb2o_1 _21343_ (.A1_N(_05467_),
    .A2_N(_05468_),
    .B1(_05467_),
    .B2(_05468_),
    .X(_05469_));
 sky130_fd_sc_hd__and4_1 _21344_ (.A(_13157_),
    .B(_13618_),
    .C(_13163_),
    .D(\pcpi_mul.rs1[3] ),
    .X(_05470_));
 sky130_fd_sc_hd__o22a_1 _21345_ (.A1(_05403_),
    .A2(_05312_),
    .B1(_05402_),
    .B2(_05335_),
    .X(_05471_));
 sky130_fd_sc_hd__or2_1 _21346_ (.A(_05470_),
    .B(_05471_),
    .X(_05472_));
 sky130_vsdinv _21347_ (.A(\pcpi_mul.rs1[7] ),
    .Y(_05473_));
 sky130_fd_sc_hd__or2_1 _21348_ (.A(_05139_),
    .B(_05473_),
    .X(_05474_));
 sky130_fd_sc_hd__a2bb2o_1 _21349_ (.A1_N(_05472_),
    .A2_N(_05474_),
    .B1(_05472_),
    .B2(_05474_),
    .X(_05475_));
 sky130_fd_sc_hd__o21ba_1 _21350_ (.A1(_05435_),
    .A2(_05437_),
    .B1_N(_05433_),
    .X(_05476_));
 sky130_fd_sc_hd__a2bb2o_1 _21351_ (.A1_N(_05475_),
    .A2_N(_05476_),
    .B1(_05475_),
    .B2(_05476_),
    .X(_05477_));
 sky130_fd_sc_hd__a2bb2o_1 _21352_ (.A1_N(_05469_),
    .A2_N(_05477_),
    .B1(_05469_),
    .B2(_05477_),
    .X(_05478_));
 sky130_fd_sc_hd__o22a_1 _21353_ (.A1(_05438_),
    .A2(_05439_),
    .B1(_05432_),
    .B2(_05440_),
    .X(_05479_));
 sky130_fd_sc_hd__a2bb2o_1 _21354_ (.A1_N(_05478_),
    .A2_N(_05479_),
    .B1(_05478_),
    .B2(_05479_),
    .X(_05480_));
 sky130_fd_sc_hd__a2bb2o_1 _21355_ (.A1_N(_05464_),
    .A2_N(_05480_),
    .B1(_05464_),
    .B2(_05480_),
    .X(_05481_));
 sky130_fd_sc_hd__or2_1 _21356_ (.A(_05463_),
    .B(_05481_),
    .X(_05482_));
 sky130_fd_sc_hd__a21bo_1 _21357_ (.A1(_05463_),
    .A2(_05481_),
    .B1_N(_05482_),
    .X(_05483_));
 sky130_fd_sc_hd__or2_1 _21358_ (.A(_05445_),
    .B(_05483_),
    .X(_05484_));
 sky130_fd_sc_hd__a21bo_1 _21359_ (.A1(_05445_),
    .A2(_05483_),
    .B1_N(_05484_),
    .X(_05485_));
 sky130_fd_sc_hd__o22a_1 _21360_ (.A1(_05441_),
    .A2(_05442_),
    .B1(_05427_),
    .B2(_05443_),
    .X(_05486_));
 sky130_fd_sc_hd__or2_1 _21361_ (.A(_05485_),
    .B(_05486_),
    .X(_05487_));
 sky130_fd_sc_hd__a21bo_1 _21362_ (.A1(_05485_),
    .A2(_05486_),
    .B1_N(_05487_),
    .X(_05488_));
 sky130_fd_sc_hd__clkbuf_2 _21363_ (.A(_05488_),
    .X(_05489_));
 sky130_fd_sc_hd__or2_1 _21364_ (.A(_05417_),
    .B(_05449_),
    .X(_05490_));
 sky130_fd_sc_hd__nand2_1 _21365_ (.A(_05448_),
    .B(_05490_),
    .Y(_05491_));
 sky130_fd_sc_hd__a2bb2oi_2 _21366_ (.A1_N(_05489_),
    .A2_N(_05491_),
    .B1(_05488_),
    .B2(_05491_),
    .Y(_05492_));
 sky130_fd_sc_hd__a2bb2oi_1 _21367_ (.A1_N(_05453_),
    .A2_N(_05492_),
    .B1(_05453_),
    .B2(_05492_),
    .Y(_02684_));
 sky130_fd_sc_hd__o22a_1 _21368_ (.A1(_05453_),
    .A2(_05492_),
    .B1(_05489_),
    .B2(_05490_),
    .X(_05493_));
 sky130_fd_sc_hd__and4_1 _21369_ (.A(_13151_),
    .B(_13621_),
    .C(\pcpi_mul.rs2[8] ),
    .D(\pcpi_mul.rs1[0] ),
    .X(_05494_));
 sky130_vsdinv _21370_ (.A(\pcpi_mul.rs2[8] ),
    .Y(_05495_));
 sky130_fd_sc_hd__o22a_1 _21371_ (.A1(_05454_),
    .A2(_05293_),
    .B1(_05495_),
    .B2(_05145_),
    .X(_05496_));
 sky130_fd_sc_hd__or2_1 _21372_ (.A(_05494_),
    .B(_05496_),
    .X(_05497_));
 sky130_fd_sc_hd__or2_1 _21373_ (.A(_05420_),
    .B(_05312_),
    .X(_05498_));
 sky130_fd_sc_hd__a2bb2o_1 _21374_ (.A1_N(_05497_),
    .A2_N(_05498_),
    .B1(_05497_),
    .B2(_05498_),
    .X(_05499_));
 sky130_fd_sc_hd__or2_1 _21375_ (.A(_05462_),
    .B(_05499_),
    .X(_05500_));
 sky130_fd_sc_hd__a21bo_1 _21376_ (.A1(_05462_),
    .A2(_05499_),
    .B1_N(_05500_),
    .X(_05501_));
 sky130_fd_sc_hd__o21ba_1 _21377_ (.A1(_05467_),
    .A2(_05468_),
    .B1_N(_05465_),
    .X(_05502_));
 sky130_fd_sc_hd__and4_1 _21378_ (.A(_05374_),
    .B(_13601_),
    .C(_05375_),
    .D(_13596_),
    .X(_05503_));
 sky130_fd_sc_hd__buf_1 _21379_ (.A(_05436_),
    .X(_05504_));
 sky130_fd_sc_hd__buf_1 _21380_ (.A(_05473_),
    .X(_05505_));
 sky130_fd_sc_hd__o22a_1 _21381_ (.A1(_05372_),
    .A2(_05504_),
    .B1(_05302_),
    .B2(_05505_),
    .X(_05506_));
 sky130_fd_sc_hd__or2_1 _21382_ (.A(_05503_),
    .B(_05506_),
    .X(_05507_));
 sky130_fd_sc_hd__buf_1 _21383_ (.A(_05398_),
    .X(_05508_));
 sky130_fd_sc_hd__clkbuf_2 _21384_ (.A(_05508_),
    .X(_05509_));
 sky130_fd_sc_hd__or2_1 _21385_ (.A(_05350_),
    .B(_05509_),
    .X(_05510_));
 sky130_fd_sc_hd__a2bb2o_1 _21386_ (.A1_N(_05507_),
    .A2_N(_05510_),
    .B1(_05507_),
    .B2(_05510_),
    .X(_05511_));
 sky130_vsdinv _21387_ (.A(\pcpi_mul.rs1[8] ),
    .Y(_05512_));
 sky130_fd_sc_hd__or2_1 _21388_ (.A(_05368_),
    .B(_05512_),
    .X(_05513_));
 sky130_fd_sc_hd__and4_1 _21389_ (.A(_13164_),
    .B(_13610_),
    .C(_13158_),
    .D(_13614_),
    .X(_05514_));
 sky130_fd_sc_hd__o22a_1 _21390_ (.A1(_05361_),
    .A2(_05364_),
    .B1(_05404_),
    .B2(_05336_),
    .X(_05515_));
 sky130_fd_sc_hd__or2_1 _21391_ (.A(_05514_),
    .B(_05515_),
    .X(_05516_));
 sky130_fd_sc_hd__a2bb2o_1 _21392_ (.A1_N(_05513_),
    .A2_N(_05516_),
    .B1(_05513_),
    .B2(_05516_),
    .X(_05517_));
 sky130_fd_sc_hd__o21ba_1 _21393_ (.A1(_05472_),
    .A2(_05474_),
    .B1_N(_05470_),
    .X(_05518_));
 sky130_fd_sc_hd__a2bb2o_1 _21394_ (.A1_N(_05517_),
    .A2_N(_05518_),
    .B1(_05517_),
    .B2(_05518_),
    .X(_05519_));
 sky130_fd_sc_hd__a2bb2o_1 _21395_ (.A1_N(_05511_),
    .A2_N(_05519_),
    .B1(_05511_),
    .B2(_05519_),
    .X(_05520_));
 sky130_fd_sc_hd__o22a_1 _21396_ (.A1(_05475_),
    .A2(_05476_),
    .B1(_05469_),
    .B2(_05477_),
    .X(_05521_));
 sky130_fd_sc_hd__a2bb2o_1 _21397_ (.A1_N(_05520_),
    .A2_N(_05521_),
    .B1(_05520_),
    .B2(_05521_),
    .X(_05522_));
 sky130_fd_sc_hd__a2bb2o_1 _21398_ (.A1_N(_05502_),
    .A2_N(_05522_),
    .B1(_05502_),
    .B2(_05522_),
    .X(_05523_));
 sky130_fd_sc_hd__nor2_2 _21399_ (.A(_05501_),
    .B(_05523_),
    .Y(_05524_));
 sky130_fd_sc_hd__a21o_1 _21400_ (.A1(_05501_),
    .A2(_05523_),
    .B1(_05524_),
    .X(_05525_));
 sky130_fd_sc_hd__or2_1 _21401_ (.A(_05482_),
    .B(_05525_),
    .X(_05526_));
 sky130_fd_sc_hd__a21bo_1 _21402_ (.A1(_05482_),
    .A2(_05525_),
    .B1_N(_05526_),
    .X(_05527_));
 sky130_fd_sc_hd__o22a_1 _21403_ (.A1(_05478_),
    .A2(_05479_),
    .B1(_05464_),
    .B2(_05480_),
    .X(_05528_));
 sky130_fd_sc_hd__a2bb2o_1 _21404_ (.A1_N(_05484_),
    .A2_N(_05528_),
    .B1(_05484_),
    .B2(_05528_),
    .X(_05529_));
 sky130_fd_sc_hd__a2bb2o_2 _21405_ (.A1_N(_05527_),
    .A2_N(_05529_),
    .B1(_05527_),
    .B2(_05529_),
    .X(_05530_));
 sky130_fd_sc_hd__o21ai_2 _21406_ (.A1(_05448_),
    .A2(_05489_),
    .B1(_05487_),
    .Y(_05531_));
 sky130_fd_sc_hd__a2bb2oi_2 _21407_ (.A1_N(_05530_),
    .A2_N(_05531_),
    .B1(_05530_),
    .B2(_05531_),
    .Y(_05532_));
 sky130_fd_sc_hd__a2bb2oi_1 _21408_ (.A1_N(_05493_),
    .A2_N(_05532_),
    .B1(_05493_),
    .B2(_05532_),
    .Y(_02685_));
 sky130_fd_sc_hd__or2_1 _21409_ (.A(_05487_),
    .B(_05530_),
    .X(_05533_));
 sky130_vsdinv _21410_ (.A(\pcpi_mul.rs2[9] ),
    .Y(_05534_));
 sky130_fd_sc_hd__buf_1 _21411_ (.A(_05534_),
    .X(_05535_));
 sky130_fd_sc_hd__buf_2 _21412_ (.A(_05535_),
    .X(_05536_));
 sky130_fd_sc_hd__buf_1 _21413_ (.A(_05536_),
    .X(_05537_));
 sky130_fd_sc_hd__buf_4 _21414_ (.A(_05537_),
    .X(_05538_));
 sky130_fd_sc_hd__or2_4 _21415_ (.A(_05538_),
    .B(_05154_),
    .X(_05539_));
 sky130_fd_sc_hd__and4_1 _21416_ (.A(\pcpi_mul.rs2[8] ),
    .B(_13621_),
    .C(\pcpi_mul.rs2[7] ),
    .D(\pcpi_mul.rs1[2] ),
    .X(_05540_));
 sky130_fd_sc_hd__o22a_1 _21417_ (.A1(_05495_),
    .A2(_05294_),
    .B1(_05454_),
    .B2(_05312_),
    .X(_05541_));
 sky130_fd_sc_hd__or2_1 _21418_ (.A(_05540_),
    .B(_05541_),
    .X(_05542_));
 sky130_fd_sc_hd__or2_1 _21419_ (.A(_05420_),
    .B(_05335_),
    .X(_05543_));
 sky130_fd_sc_hd__a2bb2o_1 _21420_ (.A1_N(_05542_),
    .A2_N(_05543_),
    .B1(_05542_),
    .B2(_05543_),
    .X(_05544_));
 sky130_fd_sc_hd__o21ba_1 _21421_ (.A1(_05497_),
    .A2(_05498_),
    .B1_N(_05494_),
    .X(_05545_));
 sky130_fd_sc_hd__or2_1 _21422_ (.A(_05544_),
    .B(_05545_),
    .X(_05546_));
 sky130_vsdinv _21423_ (.A(_05546_),
    .Y(_05547_));
 sky130_fd_sc_hd__a21o_1 _21424_ (.A1(_05544_),
    .A2(_05545_),
    .B1(_05547_),
    .X(_05548_));
 sky130_fd_sc_hd__or2_1 _21425_ (.A(_05500_),
    .B(_05548_),
    .X(_05549_));
 sky130_vsdinv _21426_ (.A(_05549_),
    .Y(_05550_));
 sky130_fd_sc_hd__a21o_1 _21427_ (.A1(_05500_),
    .A2(_05548_),
    .B1(_05550_),
    .X(_05551_));
 sky130_fd_sc_hd__o21ba_1 _21428_ (.A1(_05507_),
    .A2(_05510_),
    .B1_N(_05503_),
    .X(_05552_));
 sky130_fd_sc_hd__and4_1 _21429_ (.A(_05374_),
    .B(\pcpi_mul.rs1[7] ),
    .C(_05375_),
    .D(\pcpi_mul.rs1[8] ),
    .X(_05553_));
 sky130_fd_sc_hd__o22a_1 _21430_ (.A1(_05372_),
    .A2(_05505_),
    .B1(_05302_),
    .B2(_05512_),
    .X(_05554_));
 sky130_fd_sc_hd__or2_1 _21431_ (.A(_05553_),
    .B(_05554_),
    .X(_05555_));
 sky130_fd_sc_hd__clkbuf_2 _21432_ (.A(_05504_),
    .X(_05556_));
 sky130_fd_sc_hd__or2_1 _21433_ (.A(_05350_),
    .B(_05556_),
    .X(_05557_));
 sky130_fd_sc_hd__a2bb2o_1 _21434_ (.A1_N(_05555_),
    .A2_N(_05557_),
    .B1(_05555_),
    .B2(_05557_),
    .X(_05558_));
 sky130_fd_sc_hd__and4_1 _21435_ (.A(_13158_),
    .B(\pcpi_mul.rs1[4] ),
    .C(_13164_),
    .D(\pcpi_mul.rs1[5] ),
    .X(_05559_));
 sky130_fd_sc_hd__o22a_1 _21436_ (.A1(_05404_),
    .A2(_05364_),
    .B1(_05402_),
    .B2(_05398_),
    .X(_05560_));
 sky130_fd_sc_hd__or2_1 _21437_ (.A(_05559_),
    .B(_05560_),
    .X(_05561_));
 sky130_vsdinv _21438_ (.A(\pcpi_mul.rs1[9] ),
    .Y(_05562_));
 sky130_fd_sc_hd__or2_1 _21439_ (.A(_05368_),
    .B(_05562_),
    .X(_05563_));
 sky130_fd_sc_hd__a2bb2o_1 _21440_ (.A1_N(_05561_),
    .A2_N(_05563_),
    .B1(_05561_),
    .B2(_05563_),
    .X(_05564_));
 sky130_fd_sc_hd__o21ba_1 _21441_ (.A1(_05513_),
    .A2(_05516_),
    .B1_N(_05514_),
    .X(_05565_));
 sky130_fd_sc_hd__a2bb2o_1 _21442_ (.A1_N(_05564_),
    .A2_N(_05565_),
    .B1(_05564_),
    .B2(_05565_),
    .X(_05566_));
 sky130_fd_sc_hd__a2bb2o_1 _21443_ (.A1_N(_05558_),
    .A2_N(_05566_),
    .B1(_05558_),
    .B2(_05566_),
    .X(_05567_));
 sky130_fd_sc_hd__o22a_1 _21444_ (.A1(_05517_),
    .A2(_05518_),
    .B1(_05511_),
    .B2(_05519_),
    .X(_05568_));
 sky130_fd_sc_hd__a2bb2o_1 _21445_ (.A1_N(_05567_),
    .A2_N(_05568_),
    .B1(_05567_),
    .B2(_05568_),
    .X(_05569_));
 sky130_fd_sc_hd__a2bb2o_1 _21446_ (.A1_N(_05552_),
    .A2_N(_05569_),
    .B1(_05552_),
    .B2(_05569_),
    .X(_05570_));
 sky130_fd_sc_hd__or2_1 _21447_ (.A(_05551_),
    .B(_05570_),
    .X(_05571_));
 sky130_fd_sc_hd__a21boi_1 _21448_ (.A1(_05551_),
    .A2(_05570_),
    .B1_N(_05571_),
    .Y(_05572_));
 sky130_fd_sc_hd__nand2_1 _21449_ (.A(_05524_),
    .B(_05572_),
    .Y(_05573_));
 sky130_fd_sc_hd__o21ai_1 _21450_ (.A1(_05524_),
    .A2(_05572_),
    .B1(_05573_),
    .Y(_05574_));
 sky130_fd_sc_hd__or2_1 _21451_ (.A(_05539_),
    .B(_05574_),
    .X(_05575_));
 sky130_fd_sc_hd__a21bo_1 _21452_ (.A1(_05539_),
    .A2(_05574_),
    .B1_N(_05575_),
    .X(_05576_));
 sky130_fd_sc_hd__o22a_1 _21453_ (.A1(_05520_),
    .A2(_05521_),
    .B1(_05502_),
    .B2(_05522_),
    .X(_05577_));
 sky130_fd_sc_hd__a2bb2o_1 _21454_ (.A1_N(_05526_),
    .A2_N(_05577_),
    .B1(_05526_),
    .B2(_05577_),
    .X(_05578_));
 sky130_fd_sc_hd__a2bb2o_1 _21455_ (.A1_N(_05576_),
    .A2_N(_05578_),
    .B1(_05576_),
    .B2(_05578_),
    .X(_05579_));
 sky130_fd_sc_hd__o22a_1 _21456_ (.A1(_05484_),
    .A2(_05528_),
    .B1(_05527_),
    .B2(_05529_),
    .X(_05580_));
 sky130_fd_sc_hd__or2_1 _21457_ (.A(_05579_),
    .B(_05580_),
    .X(_05581_));
 sky130_fd_sc_hd__a21bo_1 _21458_ (.A1(_05579_),
    .A2(_05580_),
    .B1_N(_05581_),
    .X(_05582_));
 sky130_fd_sc_hd__a2bb2o_1 _21459_ (.A1_N(_05533_),
    .A2_N(_05582_),
    .B1(_05533_),
    .B2(_05582_),
    .X(_05583_));
 sky130_fd_sc_hd__o32a_1 _21460_ (.A1(_05448_),
    .A2(_05489_),
    .A3(_05530_),
    .B1(_05493_),
    .B2(_05532_),
    .X(_05584_));
 sky130_fd_sc_hd__a2bb2oi_1 _21461_ (.A1_N(_05583_),
    .A2_N(_05584_),
    .B1(_05583_),
    .B2(_05584_),
    .Y(_02686_));
 sky130_vsdinv _21462_ (.A(\pcpi_mul.rs2[10] ),
    .Y(_05585_));
 sky130_fd_sc_hd__buf_1 _21463_ (.A(_05585_),
    .X(_05586_));
 sky130_fd_sc_hd__clkbuf_2 _21464_ (.A(_05586_),
    .X(_05587_));
 sky130_fd_sc_hd__buf_2 _21465_ (.A(_05587_),
    .X(_05588_));
 sky130_fd_sc_hd__clkbuf_4 _21466_ (.A(_05588_),
    .X(_05589_));
 sky130_fd_sc_hd__buf_1 _21467_ (.A(_05153_),
    .X(_05590_));
 sky130_fd_sc_hd__o22a_2 _21468_ (.A1(_05589_),
    .A2(_05590_),
    .B1(_05538_),
    .B2(_05300_),
    .X(_05591_));
 sky130_fd_sc_hd__buf_2 _21469_ (.A(_05586_),
    .X(_05592_));
 sky130_fd_sc_hd__or4_4 _21470_ (.A(_05592_),
    .B(_05324_),
    .C(_05535_),
    .D(_05297_),
    .X(_05593_));
 sky130_fd_sc_hd__or2b_1 _21471_ (.A(_05591_),
    .B_N(_05593_),
    .X(_05594_));
 sky130_fd_sc_hd__o21ba_1 _21472_ (.A1(_05555_),
    .A2(_05557_),
    .B1_N(_05553_),
    .X(_05595_));
 sky130_fd_sc_hd__and4_1 _21473_ (.A(_05374_),
    .B(_13593_),
    .C(_05375_),
    .D(\pcpi_mul.rs1[9] ),
    .X(_05596_));
 sky130_fd_sc_hd__clkbuf_2 _21474_ (.A(_05512_),
    .X(_05597_));
 sky130_fd_sc_hd__o22a_1 _21475_ (.A1(_05372_),
    .A2(_05597_),
    .B1(_05303_),
    .B2(_05562_),
    .X(_05598_));
 sky130_fd_sc_hd__or2_1 _21476_ (.A(_05596_),
    .B(_05598_),
    .X(_05599_));
 sky130_fd_sc_hd__clkbuf_2 _21477_ (.A(_05473_),
    .X(_05600_));
 sky130_fd_sc_hd__or2_1 _21478_ (.A(_05351_),
    .B(_05600_),
    .X(_05601_));
 sky130_fd_sc_hd__a2bb2o_1 _21479_ (.A1_N(_05599_),
    .A2_N(_05601_),
    .B1(_05599_),
    .B2(_05601_),
    .X(_05602_));
 sky130_vsdinv _21480_ (.A(\pcpi_mul.rs1[10] ),
    .Y(_05603_));
 sky130_fd_sc_hd__or2_1 _21481_ (.A(_05368_),
    .B(_05603_),
    .X(_05604_));
 sky130_fd_sc_hd__and4_1 _21482_ (.A(_13158_),
    .B(_13606_),
    .C(_13164_),
    .D(_13601_),
    .X(_05605_));
 sky130_fd_sc_hd__clkbuf_2 _21483_ (.A(_05404_),
    .X(_05606_));
 sky130_fd_sc_hd__o22a_1 _21484_ (.A1(_05606_),
    .A2(_05399_),
    .B1(_05361_),
    .B2(_05504_),
    .X(_05607_));
 sky130_fd_sc_hd__or2_1 _21485_ (.A(_05605_),
    .B(_05607_),
    .X(_05608_));
 sky130_fd_sc_hd__a2bb2o_1 _21486_ (.A1_N(_05604_),
    .A2_N(_05608_),
    .B1(_05604_),
    .B2(_05608_),
    .X(_05609_));
 sky130_fd_sc_hd__o21ba_1 _21487_ (.A1(_05561_),
    .A2(_05563_),
    .B1_N(_05559_),
    .X(_05610_));
 sky130_fd_sc_hd__a2bb2o_1 _21488_ (.A1_N(_05609_),
    .A2_N(_05610_),
    .B1(_05609_),
    .B2(_05610_),
    .X(_05611_));
 sky130_fd_sc_hd__a2bb2o_1 _21489_ (.A1_N(_05602_),
    .A2_N(_05611_),
    .B1(_05602_),
    .B2(_05611_),
    .X(_05612_));
 sky130_fd_sc_hd__o22a_1 _21490_ (.A1(_05564_),
    .A2(_05565_),
    .B1(_05558_),
    .B2(_05566_),
    .X(_05613_));
 sky130_fd_sc_hd__a2bb2o_1 _21491_ (.A1_N(_05612_),
    .A2_N(_05613_),
    .B1(_05612_),
    .B2(_05613_),
    .X(_05614_));
 sky130_fd_sc_hd__a2bb2o_1 _21492_ (.A1_N(_05595_),
    .A2_N(_05614_),
    .B1(_05595_),
    .B2(_05614_),
    .X(_05615_));
 sky130_fd_sc_hd__or2_1 _21493_ (.A(_05421_),
    .B(_05369_),
    .X(_05616_));
 sky130_fd_sc_hd__o22a_1 _21494_ (.A1(_05495_),
    .A2(_05313_),
    .B1(_05455_),
    .B2(_05336_),
    .X(_05617_));
 sky130_fd_sc_hd__and4_1 _21495_ (.A(_13145_),
    .B(_05345_),
    .C(_13151_),
    .D(_13614_),
    .X(_05618_));
 sky130_fd_sc_hd__or2_1 _21496_ (.A(_05617_),
    .B(_05618_),
    .X(_05619_));
 sky130_fd_sc_hd__a2bb2o_1 _21497_ (.A1_N(_05616_),
    .A2_N(_05619_),
    .B1(_05616_),
    .B2(_05619_),
    .X(_05620_));
 sky130_fd_sc_hd__o21ba_1 _21498_ (.A1(_05542_),
    .A2(_05543_),
    .B1_N(_05540_),
    .X(_05621_));
 sky130_fd_sc_hd__or2_1 _21499_ (.A(_05620_),
    .B(_05621_),
    .X(_05622_));
 sky130_fd_sc_hd__a21bo_1 _21500_ (.A1(_05620_),
    .A2(_05621_),
    .B1_N(_05622_),
    .X(_05623_));
 sky130_fd_sc_hd__buf_1 _21501_ (.A(_05623_),
    .X(_05624_));
 sky130_fd_sc_hd__or2_2 _21502_ (.A(_05547_),
    .B(_05550_),
    .X(_05625_));
 sky130_fd_sc_hd__a2bb2oi_2 _21503_ (.A1_N(_05624_),
    .A2_N(_05625_),
    .B1(_05623_),
    .B2(_05625_),
    .Y(_05626_));
 sky130_fd_sc_hd__a2bb2o_1 _21504_ (.A1_N(_05615_),
    .A2_N(_05626_),
    .B1(_05615_),
    .B2(_05626_),
    .X(_05627_));
 sky130_fd_sc_hd__or2_1 _21505_ (.A(_05571_),
    .B(_05627_),
    .X(_05628_));
 sky130_fd_sc_hd__a21bo_1 _21506_ (.A1(_05571_),
    .A2(_05627_),
    .B1_N(_05628_),
    .X(_05629_));
 sky130_fd_sc_hd__or2_1 _21507_ (.A(_05594_),
    .B(_05629_),
    .X(_05630_));
 sky130_fd_sc_hd__a21bo_1 _21508_ (.A1(_05594_),
    .A2(_05629_),
    .B1_N(_05630_),
    .X(_05631_));
 sky130_fd_sc_hd__a2bb2o_1 _21509_ (.A1_N(_05575_),
    .A2_N(_05631_),
    .B1(_05575_),
    .B2(_05631_),
    .X(_05632_));
 sky130_fd_sc_hd__o22a_1 _21510_ (.A1(_05567_),
    .A2(_05568_),
    .B1(_05552_),
    .B2(_05569_),
    .X(_05633_));
 sky130_fd_sc_hd__or2_1 _21511_ (.A(_05573_),
    .B(_05633_),
    .X(_05634_));
 sky130_fd_sc_hd__a21bo_1 _21512_ (.A1(_05573_),
    .A2(_05633_),
    .B1_N(_05634_),
    .X(_05635_));
 sky130_fd_sc_hd__a2bb2o_1 _21513_ (.A1_N(_05632_),
    .A2_N(_05635_),
    .B1(_05632_),
    .B2(_05635_),
    .X(_05636_));
 sky130_fd_sc_hd__o22a_1 _21514_ (.A1(_05526_),
    .A2(_05577_),
    .B1(_05576_),
    .B2(_05578_),
    .X(_05637_));
 sky130_fd_sc_hd__or2_1 _21515_ (.A(_05636_),
    .B(_05637_),
    .X(_05638_));
 sky130_fd_sc_hd__a21bo_1 _21516_ (.A1(_05636_),
    .A2(_05637_),
    .B1_N(_05638_),
    .X(_05639_));
 sky130_fd_sc_hd__a2bb2o_1 _21517_ (.A1_N(_05581_),
    .A2_N(_05639_),
    .B1(_05581_),
    .B2(_05639_),
    .X(_05640_));
 sky130_fd_sc_hd__o22a_1 _21518_ (.A1(_05533_),
    .A2(_05582_),
    .B1(_05583_),
    .B2(_05584_),
    .X(_05641_));
 sky130_fd_sc_hd__a2bb2oi_1 _21519_ (.A1_N(_05640_),
    .A2_N(_05641_),
    .B1(_05640_),
    .B2(_05641_),
    .Y(_02629_));
 sky130_fd_sc_hd__o22a_1 _21520_ (.A1(_05612_),
    .A2(_05613_),
    .B1(_05595_),
    .B2(_05614_),
    .X(_05642_));
 sky130_fd_sc_hd__or2_1 _21521_ (.A(_05628_),
    .B(_05642_),
    .X(_05643_));
 sky130_fd_sc_hd__a21bo_1 _21522_ (.A1(_05628_),
    .A2(_05642_),
    .B1_N(_05643_),
    .X(_05644_));
 sky130_fd_sc_hd__buf_1 _21523_ (.A(_05314_),
    .X(_05645_));
 sky130_fd_sc_hd__or2_2 _21524_ (.A(_05534_),
    .B(_05645_),
    .X(_05646_));
 sky130_fd_sc_hd__buf_1 _21525_ (.A(_13622_),
    .X(_05647_));
 sky130_fd_sc_hd__and4_1 _21526_ (.A(_13141_),
    .B(_05647_),
    .C(\pcpi_mul.rs2[11] ),
    .D(_13625_),
    .X(_05648_));
 sky130_vsdinv _21527_ (.A(\pcpi_mul.rs2[11] ),
    .Y(_05649_));
 sky130_fd_sc_hd__o22a_1 _21528_ (.A1(_05585_),
    .A2(_05379_),
    .B1(_05649_),
    .B2(_05147_),
    .X(_05650_));
 sky130_fd_sc_hd__or2_1 _21529_ (.A(_05648_),
    .B(_05650_),
    .X(_05651_));
 sky130_fd_sc_hd__a2bb2o_1 _21530_ (.A1_N(_05646_),
    .A2_N(_05651_),
    .B1(_05646_),
    .B2(_05651_),
    .X(_05652_));
 sky130_fd_sc_hd__o21ba_1 _21531_ (.A1(_05599_),
    .A2(_05601_),
    .B1_N(_05596_),
    .X(_05653_));
 sky130_fd_sc_hd__clkbuf_2 _21532_ (.A(_13590_),
    .X(_05654_));
 sky130_fd_sc_hd__clkbuf_2 _21533_ (.A(\pcpi_mul.rs1[10] ),
    .X(_05655_));
 sky130_fd_sc_hd__and4_1 _21534_ (.A(_13172_),
    .B(_05654_),
    .C(_13177_),
    .D(_05655_),
    .X(_05656_));
 sky130_fd_sc_hd__buf_2 _21535_ (.A(_05562_),
    .X(_05657_));
 sky130_fd_sc_hd__clkbuf_2 _21536_ (.A(_05603_),
    .X(_05658_));
 sky130_fd_sc_hd__o22a_1 _21537_ (.A1(_05321_),
    .A2(_05657_),
    .B1(_05304_),
    .B2(_05658_),
    .X(_05659_));
 sky130_fd_sc_hd__or2_1 _21538_ (.A(_05656_),
    .B(_05659_),
    .X(_05660_));
 sky130_fd_sc_hd__buf_2 _21539_ (.A(_05351_),
    .X(_05661_));
 sky130_fd_sc_hd__buf_1 _21540_ (.A(_05597_),
    .X(_05662_));
 sky130_fd_sc_hd__clkbuf_4 _21541_ (.A(_05662_),
    .X(_05663_));
 sky130_fd_sc_hd__or2_1 _21542_ (.A(_05661_),
    .B(_05663_),
    .X(_05664_));
 sky130_fd_sc_hd__a2bb2o_1 _21543_ (.A1_N(_05660_),
    .A2_N(_05664_),
    .B1(_05660_),
    .B2(_05664_),
    .X(_05665_));
 sky130_vsdinv _21544_ (.A(\pcpi_mul.rs1[11] ),
    .Y(_05666_));
 sky130_fd_sc_hd__clkbuf_2 _21545_ (.A(_05666_),
    .X(_05667_));
 sky130_fd_sc_hd__or2_2 _21546_ (.A(_05140_),
    .B(_05667_),
    .X(_05668_));
 sky130_fd_sc_hd__and4_1 _21547_ (.A(_13159_),
    .B(_13602_),
    .C(_13165_),
    .D(_13596_),
    .X(_05669_));
 sky130_fd_sc_hd__o22a_1 _21548_ (.A1(_05606_),
    .A2(_05556_),
    .B1(_05362_),
    .B2(_05505_),
    .X(_05670_));
 sky130_fd_sc_hd__or2_1 _21549_ (.A(_05669_),
    .B(_05670_),
    .X(_05671_));
 sky130_fd_sc_hd__a2bb2o_1 _21550_ (.A1_N(_05668_),
    .A2_N(_05671_),
    .B1(_05668_),
    .B2(_05671_),
    .X(_05672_));
 sky130_fd_sc_hd__o21ba_1 _21551_ (.A1(_05604_),
    .A2(_05608_),
    .B1_N(_05605_),
    .X(_05673_));
 sky130_fd_sc_hd__a2bb2o_1 _21552_ (.A1_N(_05672_),
    .A2_N(_05673_),
    .B1(_05672_),
    .B2(_05673_),
    .X(_05674_));
 sky130_fd_sc_hd__a2bb2o_1 _21553_ (.A1_N(_05665_),
    .A2_N(_05674_),
    .B1(_05665_),
    .B2(_05674_),
    .X(_05675_));
 sky130_fd_sc_hd__o22a_1 _21554_ (.A1(_05609_),
    .A2(_05610_),
    .B1(_05602_),
    .B2(_05611_),
    .X(_05676_));
 sky130_fd_sc_hd__a2bb2o_1 _21555_ (.A1_N(_05675_),
    .A2_N(_05676_),
    .B1(_05675_),
    .B2(_05676_),
    .X(_05677_));
 sky130_fd_sc_hd__a2bb2o_1 _21556_ (.A1_N(_05653_),
    .A2_N(_05677_),
    .B1(_05653_),
    .B2(_05677_),
    .X(_05678_));
 sky130_fd_sc_hd__o21ba_1 _21557_ (.A1(_05616_),
    .A2(_05619_),
    .B1_N(_05618_),
    .X(_05679_));
 sky130_fd_sc_hd__clkbuf_2 _21558_ (.A(_05508_),
    .X(_05680_));
 sky130_fd_sc_hd__or2_1 _21559_ (.A(_05421_),
    .B(_05680_),
    .X(_05681_));
 sky130_fd_sc_hd__clkbuf_4 _21560_ (.A(_05495_),
    .X(_05682_));
 sky130_fd_sc_hd__clkbuf_2 _21561_ (.A(_05336_),
    .X(_05683_));
 sky130_fd_sc_hd__clkbuf_2 _21562_ (.A(_05365_),
    .X(_05684_));
 sky130_fd_sc_hd__o22a_1 _21563_ (.A1(_05682_),
    .A2(_05683_),
    .B1(_05455_),
    .B2(_05684_),
    .X(_05685_));
 sky130_fd_sc_hd__and4_1 _21564_ (.A(_13145_),
    .B(_13615_),
    .C(_13151_),
    .D(_13611_),
    .X(_05686_));
 sky130_fd_sc_hd__or2_1 _21565_ (.A(_05685_),
    .B(_05686_),
    .X(_05687_));
 sky130_fd_sc_hd__a2bb2o_1 _21566_ (.A1_N(_05681_),
    .A2_N(_05687_),
    .B1(_05681_),
    .B2(_05687_),
    .X(_05688_));
 sky130_fd_sc_hd__a2bb2o_1 _21567_ (.A1_N(_05593_),
    .A2_N(_05688_),
    .B1(_05593_),
    .B2(_05688_),
    .X(_05689_));
 sky130_fd_sc_hd__a2bb2o_2 _21568_ (.A1_N(_05679_),
    .A2_N(_05689_),
    .B1(_05679_),
    .B2(_05689_),
    .X(_05690_));
 sky130_fd_sc_hd__o21ai_1 _21569_ (.A1(_05546_),
    .A2(_05624_),
    .B1(_05622_),
    .Y(_05691_));
 sky130_fd_sc_hd__a2bb2oi_1 _21570_ (.A1_N(_05690_),
    .A2_N(_05691_),
    .B1(_05690_),
    .B2(_05691_),
    .Y(_05692_));
 sky130_fd_sc_hd__a2bb2o_1 _21571_ (.A1_N(_05678_),
    .A2_N(_05692_),
    .B1(_05678_),
    .B2(_05692_),
    .X(_05693_));
 sky130_fd_sc_hd__o22a_1 _21572_ (.A1(_05615_),
    .A2(_05626_),
    .B1(_05549_),
    .B2(_05624_),
    .X(_05694_));
 sky130_fd_sc_hd__or2_1 _21573_ (.A(_05693_),
    .B(_05694_),
    .X(_05695_));
 sky130_fd_sc_hd__a21bo_1 _21574_ (.A1(_05693_),
    .A2(_05694_),
    .B1_N(_05695_),
    .X(_05696_));
 sky130_fd_sc_hd__or2_1 _21575_ (.A(_05652_),
    .B(_05696_),
    .X(_05697_));
 sky130_fd_sc_hd__a21bo_1 _21576_ (.A1(_05652_),
    .A2(_05696_),
    .B1_N(_05697_),
    .X(_05698_));
 sky130_fd_sc_hd__a2bb2o_1 _21577_ (.A1_N(_05630_),
    .A2_N(_05698_),
    .B1(_05630_),
    .B2(_05698_),
    .X(_05699_));
 sky130_fd_sc_hd__a2bb2o_1 _21578_ (.A1_N(_05644_),
    .A2_N(_05699_),
    .B1(_05644_),
    .B2(_05699_),
    .X(_05700_));
 sky130_fd_sc_hd__o22a_1 _21579_ (.A1(_05575_),
    .A2(_05631_),
    .B1(_05632_),
    .B2(_05635_),
    .X(_05701_));
 sky130_fd_sc_hd__a2bb2o_1 _21580_ (.A1_N(_05700_),
    .A2_N(_05701_),
    .B1(_05700_),
    .B2(_05701_),
    .X(_05702_));
 sky130_fd_sc_hd__a2bb2o_1 _21581_ (.A1_N(_05634_),
    .A2_N(_05702_),
    .B1(_05634_),
    .B2(_05702_),
    .X(_05703_));
 sky130_fd_sc_hd__a2bb2o_1 _21582_ (.A1_N(_05638_),
    .A2_N(_05703_),
    .B1(_05638_),
    .B2(_05703_),
    .X(_05704_));
 sky130_fd_sc_hd__o22a_1 _21583_ (.A1(_05581_),
    .A2(_05639_),
    .B1(_05640_),
    .B2(_05641_),
    .X(_05705_));
 sky130_fd_sc_hd__a2bb2oi_1 _21584_ (.A1_N(_05704_),
    .A2_N(_05705_),
    .B1(_05704_),
    .B2(_05705_),
    .Y(_02630_));
 sky130_vsdinv _21585_ (.A(\pcpi_mul.rs2[12] ),
    .Y(_05706_));
 sky130_fd_sc_hd__buf_1 _21586_ (.A(_05706_),
    .X(_05707_));
 sky130_fd_sc_hd__clkbuf_4 _21587_ (.A(_05707_),
    .X(_05708_));
 sky130_fd_sc_hd__clkbuf_4 _21588_ (.A(_05708_),
    .X(_05709_));
 sky130_fd_sc_hd__or2_2 _21589_ (.A(_05709_),
    .B(_05151_),
    .X(_05710_));
 sky130_fd_sc_hd__clkbuf_2 _21590_ (.A(_05535_),
    .X(_05711_));
 sky130_fd_sc_hd__or2_1 _21591_ (.A(_05711_),
    .B(_05340_),
    .X(_05712_));
 sky130_fd_sc_hd__buf_1 _21592_ (.A(_05649_),
    .X(_05713_));
 sky130_fd_sc_hd__buf_2 _21593_ (.A(_05713_),
    .X(_05714_));
 sky130_fd_sc_hd__o22a_1 _21594_ (.A1(_05714_),
    .A2(_05318_),
    .B1(_05587_),
    .B2(_05315_),
    .X(_05715_));
 sky130_fd_sc_hd__and4_1 _21595_ (.A(_13136_),
    .B(_13624_),
    .C(_13142_),
    .D(_13620_),
    .X(_05716_));
 sky130_fd_sc_hd__or2_1 _21596_ (.A(_05715_),
    .B(_05716_),
    .X(_05717_));
 sky130_fd_sc_hd__a2bb2o_1 _21597_ (.A1_N(_05712_),
    .A2_N(_05717_),
    .B1(_05712_),
    .B2(_05717_),
    .X(_05718_));
 sky130_fd_sc_hd__or2_1 _21598_ (.A(_05710_),
    .B(_05718_),
    .X(_05719_));
 sky130_fd_sc_hd__a21bo_1 _21599_ (.A1(_05710_),
    .A2(_05718_),
    .B1_N(_05719_),
    .X(_05720_));
 sky130_fd_sc_hd__o21ba_1 _21600_ (.A1(_05660_),
    .A2(_05664_),
    .B1_N(_05656_),
    .X(_05721_));
 sky130_fd_sc_hd__buf_1 _21601_ (.A(_05658_),
    .X(_05722_));
 sky130_fd_sc_hd__clkbuf_2 _21602_ (.A(_05722_),
    .X(_05723_));
 sky130_fd_sc_hd__clkbuf_2 _21603_ (.A(_05666_),
    .X(_05724_));
 sky130_fd_sc_hd__clkbuf_2 _21604_ (.A(_05724_),
    .X(_05725_));
 sky130_fd_sc_hd__o22a_2 _21605_ (.A1(_05323_),
    .A2(_05723_),
    .B1(_05306_),
    .B2(_05725_),
    .X(_05726_));
 sky130_fd_sc_hd__and4_2 _21606_ (.A(_13173_),
    .B(_13588_),
    .C(_13178_),
    .D(_13585_),
    .X(_05727_));
 sky130_fd_sc_hd__nor2_2 _21607_ (.A(_05726_),
    .B(_05727_),
    .Y(_05728_));
 sky130_fd_sc_hd__buf_1 _21608_ (.A(_05657_),
    .X(_05729_));
 sky130_fd_sc_hd__buf_1 _21609_ (.A(_05729_),
    .X(_05730_));
 sky130_fd_sc_hd__buf_2 _21610_ (.A(_05730_),
    .X(_05731_));
 sky130_fd_sc_hd__nor2_2 _21611_ (.A(_05661_),
    .B(_05731_),
    .Y(_05732_));
 sky130_fd_sc_hd__a2bb2o_1 _21612_ (.A1_N(_05728_),
    .A2_N(_05732_),
    .B1(_05728_),
    .B2(_05732_),
    .X(_05733_));
 sky130_vsdinv _21613_ (.A(\pcpi_mul.rs1[12] ),
    .Y(_05734_));
 sky130_fd_sc_hd__clkbuf_2 _21614_ (.A(_05734_),
    .X(_05735_));
 sky130_fd_sc_hd__or2_1 _21615_ (.A(_05141_),
    .B(_05735_),
    .X(_05736_));
 sky130_fd_sc_hd__clkbuf_4 _21616_ (.A(_05606_),
    .X(_05737_));
 sky130_fd_sc_hd__clkbuf_2 _21617_ (.A(_05505_),
    .X(_05738_));
 sky130_fd_sc_hd__clkbuf_4 _21618_ (.A(_05362_),
    .X(_05739_));
 sky130_fd_sc_hd__o22a_1 _21619_ (.A1(_05737_),
    .A2(_05738_),
    .B1(_05739_),
    .B2(_05662_),
    .X(_05740_));
 sky130_fd_sc_hd__buf_1 _21620_ (.A(_13596_),
    .X(_05741_));
 sky130_fd_sc_hd__buf_1 _21621_ (.A(_13593_),
    .X(_05742_));
 sky130_fd_sc_hd__and4_1 _21622_ (.A(_13159_),
    .B(_05741_),
    .C(_13165_),
    .D(_05742_),
    .X(_05743_));
 sky130_fd_sc_hd__or2_1 _21623_ (.A(_05740_),
    .B(_05743_),
    .X(_05744_));
 sky130_fd_sc_hd__a2bb2o_2 _21624_ (.A1_N(_05736_),
    .A2_N(_05744_),
    .B1(_05736_),
    .B2(_05744_),
    .X(_05745_));
 sky130_fd_sc_hd__o21ba_1 _21625_ (.A1(_05668_),
    .A2(_05671_),
    .B1_N(_05669_),
    .X(_05746_));
 sky130_fd_sc_hd__a2bb2o_1 _21626_ (.A1_N(_05745_),
    .A2_N(_05746_),
    .B1(_05745_),
    .B2(_05746_),
    .X(_05747_));
 sky130_fd_sc_hd__a2bb2o_1 _21627_ (.A1_N(_05733_),
    .A2_N(_05747_),
    .B1(_05733_),
    .B2(_05747_),
    .X(_05748_));
 sky130_fd_sc_hd__o22a_1 _21628_ (.A1(_05672_),
    .A2(_05673_),
    .B1(_05665_),
    .B2(_05674_),
    .X(_05749_));
 sky130_fd_sc_hd__a2bb2o_1 _21629_ (.A1_N(_05748_),
    .A2_N(_05749_),
    .B1(_05748_),
    .B2(_05749_),
    .X(_05750_));
 sky130_fd_sc_hd__a2bb2o_1 _21630_ (.A1_N(_05721_),
    .A2_N(_05750_),
    .B1(_05721_),
    .B2(_05750_),
    .X(_05751_));
 sky130_fd_sc_hd__or2_1 _21631_ (.A(_05622_),
    .B(_05690_),
    .X(_05752_));
 sky130_fd_sc_hd__o21ba_1 _21632_ (.A1(_05681_),
    .A2(_05687_),
    .B1_N(_05686_),
    .X(_05753_));
 sky130_fd_sc_hd__o21ba_1 _21633_ (.A1(_05646_),
    .A2(_05651_),
    .B1_N(_05648_),
    .X(_05754_));
 sky130_fd_sc_hd__buf_1 _21634_ (.A(_05556_),
    .X(_05755_));
 sky130_fd_sc_hd__or2_2 _21635_ (.A(_05422_),
    .B(_05755_),
    .X(_05756_));
 sky130_fd_sc_hd__o22a_1 _21636_ (.A1(_05682_),
    .A2(_05684_),
    .B1(_05456_),
    .B2(_05508_),
    .X(_05757_));
 sky130_fd_sc_hd__buf_1 _21637_ (.A(_13610_),
    .X(_05758_));
 sky130_fd_sc_hd__and4_1 _21638_ (.A(_13145_),
    .B(_05758_),
    .C(_13152_),
    .D(_13607_),
    .X(_05759_));
 sky130_fd_sc_hd__or2_1 _21639_ (.A(_05757_),
    .B(_05759_),
    .X(_05760_));
 sky130_fd_sc_hd__a2bb2o_1 _21640_ (.A1_N(_05756_),
    .A2_N(_05760_),
    .B1(_05756_),
    .B2(_05760_),
    .X(_05761_));
 sky130_fd_sc_hd__a2bb2o_1 _21641_ (.A1_N(_05754_),
    .A2_N(_05761_),
    .B1(_05754_),
    .B2(_05761_),
    .X(_05762_));
 sky130_fd_sc_hd__a2bb2o_1 _21642_ (.A1_N(_05753_),
    .A2_N(_05762_),
    .B1(_05753_),
    .B2(_05762_),
    .X(_05763_));
 sky130_fd_sc_hd__o22a_1 _21643_ (.A1(_05593_),
    .A2(_05688_),
    .B1(_05679_),
    .B2(_05689_),
    .X(_05764_));
 sky130_fd_sc_hd__or2_1 _21644_ (.A(_05763_),
    .B(_05764_),
    .X(_05765_));
 sky130_fd_sc_hd__a21bo_1 _21645_ (.A1(_05763_),
    .A2(_05764_),
    .B1_N(_05765_),
    .X(_05766_));
 sky130_fd_sc_hd__a2bb2o_1 _21646_ (.A1_N(_05752_),
    .A2_N(_05766_),
    .B1(_05752_),
    .B2(_05766_),
    .X(_05767_));
 sky130_fd_sc_hd__a2bb2o_1 _21647_ (.A1_N(_05751_),
    .A2_N(_05767_),
    .B1(_05751_),
    .B2(_05767_),
    .X(_05768_));
 sky130_fd_sc_hd__o32a_1 _21648_ (.A1(_05546_),
    .A2(_05624_),
    .A3(_05690_),
    .B1(_05678_),
    .B2(_05692_),
    .X(_05769_));
 sky130_fd_sc_hd__or2_1 _21649_ (.A(_05768_),
    .B(_05769_),
    .X(_05770_));
 sky130_fd_sc_hd__a21bo_1 _21650_ (.A1(_05768_),
    .A2(_05769_),
    .B1_N(_05770_),
    .X(_05771_));
 sky130_fd_sc_hd__or2_1 _21651_ (.A(_05720_),
    .B(_05771_),
    .X(_05772_));
 sky130_fd_sc_hd__a21bo_1 _21652_ (.A1(_05720_),
    .A2(_05771_),
    .B1_N(_05772_),
    .X(_05773_));
 sky130_fd_sc_hd__a2bb2o_1 _21653_ (.A1_N(_05697_),
    .A2_N(_05773_),
    .B1(_05697_),
    .B2(_05773_),
    .X(_05774_));
 sky130_fd_sc_hd__o22a_1 _21654_ (.A1(_05675_),
    .A2(_05676_),
    .B1(_05653_),
    .B2(_05677_),
    .X(_05775_));
 sky130_fd_sc_hd__or2_1 _21655_ (.A(_05695_),
    .B(_05775_),
    .X(_05776_));
 sky130_fd_sc_hd__a21bo_1 _21656_ (.A1(_05695_),
    .A2(_05775_),
    .B1_N(_05776_),
    .X(_05777_));
 sky130_fd_sc_hd__a2bb2o_1 _21657_ (.A1_N(_05774_),
    .A2_N(_05777_),
    .B1(_05774_),
    .B2(_05777_),
    .X(_05778_));
 sky130_fd_sc_hd__o22a_1 _21658_ (.A1(_05630_),
    .A2(_05698_),
    .B1(_05644_),
    .B2(_05699_),
    .X(_05779_));
 sky130_fd_sc_hd__a2bb2o_1 _21659_ (.A1_N(_05778_),
    .A2_N(_05779_),
    .B1(_05778_),
    .B2(_05779_),
    .X(_05780_));
 sky130_fd_sc_hd__a2bb2o_1 _21660_ (.A1_N(_05643_),
    .A2_N(_05780_),
    .B1(_05643_),
    .B2(_05780_),
    .X(_05781_));
 sky130_fd_sc_hd__o22a_1 _21661_ (.A1(_05700_),
    .A2(_05701_),
    .B1(_05634_),
    .B2(_05702_),
    .X(_05782_));
 sky130_fd_sc_hd__a2bb2o_1 _21662_ (.A1_N(_05781_),
    .A2_N(_05782_),
    .B1(_05781_),
    .B2(_05782_),
    .X(_05783_));
 sky130_fd_sc_hd__o22a_1 _21663_ (.A1(_05638_),
    .A2(_05703_),
    .B1(_05704_),
    .B2(_05705_),
    .X(_05784_));
 sky130_fd_sc_hd__a2bb2oi_1 _21664_ (.A1_N(_05783_),
    .A2_N(_05784_),
    .B1(_05783_),
    .B2(_05784_),
    .Y(_02631_));
 sky130_fd_sc_hd__o22a_2 _21665_ (.A1(_05781_),
    .A2(_05782_),
    .B1(_05783_),
    .B2(_05784_),
    .X(_05785_));
 sky130_vsdinv _21666_ (.A(\pcpi_mul.rs2[13] ),
    .Y(_05786_));
 sky130_fd_sc_hd__clkbuf_2 _21667_ (.A(_05786_),
    .X(_05787_));
 sky130_fd_sc_hd__buf_2 _21668_ (.A(_05787_),
    .X(_05788_));
 sky130_fd_sc_hd__clkbuf_4 _21669_ (.A(_05788_),
    .X(_05789_));
 sky130_fd_sc_hd__clkbuf_2 _21670_ (.A(_05706_),
    .X(_05790_));
 sky130_fd_sc_hd__clkbuf_4 _21671_ (.A(_05790_),
    .X(_05791_));
 sky130_fd_sc_hd__buf_1 _21672_ (.A(_05297_),
    .X(_05792_));
 sky130_fd_sc_hd__o22a_1 _21673_ (.A1(_05789_),
    .A2(_05459_),
    .B1(_05791_),
    .B2(_05792_),
    .X(_05793_));
 sky130_fd_sc_hd__clkbuf_4 _21674_ (.A(_05707_),
    .X(_05794_));
 sky130_fd_sc_hd__or4_4 _21675_ (.A(_05789_),
    .B(_05325_),
    .C(_05794_),
    .D(_05792_),
    .X(_05795_));
 sky130_fd_sc_hd__or2b_1 _21676_ (.A(_05793_),
    .B_N(_05795_),
    .X(_05796_));
 sky130_fd_sc_hd__buf_1 _21677_ (.A(_05534_),
    .X(_05797_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _21678_ (.A(_05684_),
    .X(_05798_));
 sky130_fd_sc_hd__clkbuf_2 _21679_ (.A(_05798_),
    .X(_05799_));
 sky130_fd_sc_hd__or2_1 _21680_ (.A(_05797_),
    .B(_05799_),
    .X(_05800_));
 sky130_fd_sc_hd__buf_1 _21681_ (.A(_05649_),
    .X(_05801_));
 sky130_fd_sc_hd__clkbuf_2 _21682_ (.A(_05585_),
    .X(_05802_));
 sky130_fd_sc_hd__clkbuf_2 _21683_ (.A(_05683_),
    .X(_05803_));
 sky130_fd_sc_hd__o22a_1 _21684_ (.A1(_05801_),
    .A2(_05645_),
    .B1(_05802_),
    .B2(_05803_),
    .X(_05804_));
 sky130_fd_sc_hd__buf_1 _21685_ (.A(\pcpi_mul.rs2[11] ),
    .X(_05805_));
 sky130_fd_sc_hd__buf_1 _21686_ (.A(_13619_),
    .X(_05806_));
 sky130_fd_sc_hd__buf_1 _21687_ (.A(\pcpi_mul.rs2[10] ),
    .X(_05807_));
 sky130_fd_sc_hd__buf_1 _21688_ (.A(_13615_),
    .X(_05808_));
 sky130_fd_sc_hd__and4_1 _21689_ (.A(_05805_),
    .B(_05806_),
    .C(_05807_),
    .D(_05808_),
    .X(_05809_));
 sky130_fd_sc_hd__or2_1 _21690_ (.A(_05804_),
    .B(_05809_),
    .X(_05810_));
 sky130_fd_sc_hd__a2bb2o_1 _21691_ (.A1_N(_05800_),
    .A2_N(_05810_),
    .B1(_05800_),
    .B2(_05810_),
    .X(_05811_));
 sky130_fd_sc_hd__or2_1 _21692_ (.A(_05796_),
    .B(_05811_),
    .X(_05812_));
 sky130_fd_sc_hd__a21bo_1 _21693_ (.A1(_05796_),
    .A2(_05811_),
    .B1_N(_05812_),
    .X(_05813_));
 sky130_fd_sc_hd__o22a_1 _21694_ (.A1(_05752_),
    .A2(_05766_),
    .B1(_05751_),
    .B2(_05767_),
    .X(_05814_));
 sky130_fd_sc_hd__a21oi_2 _21695_ (.A1(_05728_),
    .A2(_05732_),
    .B1(_05727_),
    .Y(_05815_));
 sky130_fd_sc_hd__buf_2 _21696_ (.A(_05323_),
    .X(_05816_));
 sky130_fd_sc_hd__clkbuf_2 _21697_ (.A(_05667_),
    .X(_05817_));
 sky130_fd_sc_hd__buf_2 _21698_ (.A(_05817_),
    .X(_05818_));
 sky130_fd_sc_hd__clkbuf_2 _21699_ (.A(_05734_),
    .X(_05819_));
 sky130_fd_sc_hd__buf_1 _21700_ (.A(_05819_),
    .X(_05820_));
 sky130_fd_sc_hd__buf_2 _21701_ (.A(_05820_),
    .X(_05821_));
 sky130_fd_sc_hd__o22a_1 _21702_ (.A1(_05816_),
    .A2(_05818_),
    .B1(_05307_),
    .B2(_05821_),
    .X(_05822_));
 sky130_fd_sc_hd__clkbuf_2 _21703_ (.A(_13173_),
    .X(_05823_));
 sky130_fd_sc_hd__clkbuf_2 _21704_ (.A(_13178_),
    .X(_05824_));
 sky130_fd_sc_hd__and4_2 _21705_ (.A(_05823_),
    .B(_13585_),
    .C(_05824_),
    .D(_13583_),
    .X(_05825_));
 sky130_fd_sc_hd__nor2_2 _21706_ (.A(_05822_),
    .B(_05825_),
    .Y(_05826_));
 sky130_fd_sc_hd__buf_4 _21707_ (.A(_05661_),
    .X(_05827_));
 sky130_fd_sc_hd__buf_2 _21708_ (.A(_05827_),
    .X(_05828_));
 sky130_fd_sc_hd__buf_2 _21709_ (.A(_05603_),
    .X(_05829_));
 sky130_fd_sc_hd__clkbuf_2 _21710_ (.A(_05829_),
    .X(_05830_));
 sky130_fd_sc_hd__buf_2 _21711_ (.A(_05830_),
    .X(_05831_));
 sky130_fd_sc_hd__nor2_2 _21712_ (.A(_05828_),
    .B(_05831_),
    .Y(_05832_));
 sky130_fd_sc_hd__a2bb2o_1 _21713_ (.A1_N(_05826_),
    .A2_N(_05832_),
    .B1(_05826_),
    .B2(_05832_),
    .X(_05833_));
 sky130_fd_sc_hd__buf_1 _21714_ (.A(_05141_),
    .X(_05834_));
 sky130_vsdinv _21715_ (.A(\pcpi_mul.rs1[13] ),
    .Y(_05835_));
 sky130_fd_sc_hd__clkbuf_2 _21716_ (.A(_05835_),
    .X(_05836_));
 sky130_fd_sc_hd__clkbuf_2 _21717_ (.A(_05836_),
    .X(_05837_));
 sky130_fd_sc_hd__or2_2 _21718_ (.A(_05834_),
    .B(_05837_),
    .X(_05838_));
 sky130_fd_sc_hd__buf_1 _21719_ (.A(_05606_),
    .X(_05839_));
 sky130_fd_sc_hd__buf_1 _21720_ (.A(_05597_),
    .X(_05840_));
 sky130_fd_sc_hd__clkbuf_2 _21721_ (.A(_05840_),
    .X(_05841_));
 sky130_fd_sc_hd__buf_1 _21722_ (.A(_05362_),
    .X(_05842_));
 sky130_fd_sc_hd__clkbuf_2 _21723_ (.A(_05729_),
    .X(_05843_));
 sky130_fd_sc_hd__o22a_1 _21724_ (.A1(_05839_),
    .A2(_05841_),
    .B1(_05842_),
    .B2(_05843_),
    .X(_05844_));
 sky130_fd_sc_hd__buf_1 _21725_ (.A(_13159_),
    .X(_05845_));
 sky130_fd_sc_hd__buf_1 _21726_ (.A(_05742_),
    .X(_05846_));
 sky130_fd_sc_hd__buf_1 _21727_ (.A(_13165_),
    .X(_05847_));
 sky130_fd_sc_hd__buf_1 _21728_ (.A(_13590_),
    .X(_05848_));
 sky130_fd_sc_hd__and4_1 _21729_ (.A(_05845_),
    .B(_05846_),
    .C(_05847_),
    .D(_05848_),
    .X(_05849_));
 sky130_fd_sc_hd__or2_1 _21730_ (.A(_05844_),
    .B(_05849_),
    .X(_05850_));
 sky130_fd_sc_hd__a2bb2o_1 _21731_ (.A1_N(_05838_),
    .A2_N(_05850_),
    .B1(_05838_),
    .B2(_05850_),
    .X(_05851_));
 sky130_fd_sc_hd__o21ba_1 _21732_ (.A1(_05736_),
    .A2(_05744_),
    .B1_N(_05743_),
    .X(_05852_));
 sky130_fd_sc_hd__a2bb2o_1 _21733_ (.A1_N(_05851_),
    .A2_N(_05852_),
    .B1(_05851_),
    .B2(_05852_),
    .X(_05853_));
 sky130_fd_sc_hd__a2bb2o_2 _21734_ (.A1_N(_05833_),
    .A2_N(_05853_),
    .B1(_05833_),
    .B2(_05853_),
    .X(_05854_));
 sky130_fd_sc_hd__o22a_1 _21735_ (.A1(_05745_),
    .A2(_05746_),
    .B1(_05733_),
    .B2(_05747_),
    .X(_05855_));
 sky130_fd_sc_hd__a2bb2o_1 _21736_ (.A1_N(_05854_),
    .A2_N(_05855_),
    .B1(_05854_),
    .B2(_05855_),
    .X(_05856_));
 sky130_fd_sc_hd__a2bb2o_1 _21737_ (.A1_N(_05815_),
    .A2_N(_05856_),
    .B1(_05815_),
    .B2(_05856_),
    .X(_05857_));
 sky130_fd_sc_hd__o22a_1 _21738_ (.A1(_05754_),
    .A2(_05761_),
    .B1(_05753_),
    .B2(_05762_),
    .X(_05858_));
 sky130_fd_sc_hd__o21ba_1 _21739_ (.A1(_05756_),
    .A2(_05760_),
    .B1_N(_05759_),
    .X(_05859_));
 sky130_fd_sc_hd__o21ba_1 _21740_ (.A1(_05712_),
    .A2(_05717_),
    .B1_N(_05716_),
    .X(_05860_));
 sky130_fd_sc_hd__clkbuf_2 _21741_ (.A(_05600_),
    .X(_05861_));
 sky130_fd_sc_hd__clkbuf_2 _21742_ (.A(_05861_),
    .X(_05862_));
 sky130_fd_sc_hd__or2_1 _21743_ (.A(_05460_),
    .B(_05862_),
    .X(_05863_));
 sky130_fd_sc_hd__clkbuf_2 _21744_ (.A(_05682_),
    .X(_05864_));
 sky130_fd_sc_hd__clkbuf_2 _21745_ (.A(_05864_),
    .X(_05865_));
 sky130_fd_sc_hd__buf_2 _21746_ (.A(_05509_),
    .X(_05866_));
 sky130_fd_sc_hd__buf_2 _21747_ (.A(_05504_),
    .X(_05867_));
 sky130_fd_sc_hd__buf_1 _21748_ (.A(_05867_),
    .X(_05868_));
 sky130_fd_sc_hd__o22a_1 _21749_ (.A1(_05865_),
    .A2(_05866_),
    .B1(_05457_),
    .B2(_05868_),
    .X(_05869_));
 sky130_fd_sc_hd__clkbuf_2 _21750_ (.A(_13146_),
    .X(_05870_));
 sky130_fd_sc_hd__clkbuf_2 _21751_ (.A(_13152_),
    .X(_05871_));
 sky130_fd_sc_hd__clkbuf_2 _21752_ (.A(_13602_),
    .X(_05872_));
 sky130_fd_sc_hd__and4_1 _21753_ (.A(_05870_),
    .B(_13608_),
    .C(_05871_),
    .D(_05872_),
    .X(_05873_));
 sky130_fd_sc_hd__or2_1 _21754_ (.A(_05869_),
    .B(_05873_),
    .X(_05874_));
 sky130_fd_sc_hd__a2bb2o_2 _21755_ (.A1_N(_05863_),
    .A2_N(_05874_),
    .B1(_05863_),
    .B2(_05874_),
    .X(_05875_));
 sky130_fd_sc_hd__a2bb2o_1 _21756_ (.A1_N(_05860_),
    .A2_N(_05875_),
    .B1(_05860_),
    .B2(_05875_),
    .X(_05876_));
 sky130_fd_sc_hd__a2bb2o_1 _21757_ (.A1_N(_05859_),
    .A2_N(_05876_),
    .B1(_05859_),
    .B2(_05876_),
    .X(_05877_));
 sky130_fd_sc_hd__a2bb2o_1 _21758_ (.A1_N(_05719_),
    .A2_N(_05877_),
    .B1(_05719_),
    .B2(_05877_),
    .X(_05878_));
 sky130_fd_sc_hd__a2bb2o_1 _21759_ (.A1_N(_05858_),
    .A2_N(_05878_),
    .B1(_05858_),
    .B2(_05878_),
    .X(_05879_));
 sky130_fd_sc_hd__a2bb2o_1 _21760_ (.A1_N(_05765_),
    .A2_N(_05879_),
    .B1(_05765_),
    .B2(_05879_),
    .X(_05880_));
 sky130_fd_sc_hd__a2bb2o_1 _21761_ (.A1_N(_05857_),
    .A2_N(_05880_),
    .B1(_05857_),
    .B2(_05880_),
    .X(_05881_));
 sky130_fd_sc_hd__or2_1 _21762_ (.A(_05814_),
    .B(_05881_),
    .X(_05882_));
 sky130_fd_sc_hd__a21bo_1 _21763_ (.A1(_05814_),
    .A2(_05881_),
    .B1_N(_05882_),
    .X(_05883_));
 sky130_fd_sc_hd__or2_1 _21764_ (.A(_05813_),
    .B(_05883_),
    .X(_05884_));
 sky130_fd_sc_hd__a21bo_1 _21765_ (.A1(_05813_),
    .A2(_05883_),
    .B1_N(_05884_),
    .X(_05885_));
 sky130_fd_sc_hd__a2bb2o_1 _21766_ (.A1_N(_05772_),
    .A2_N(_05885_),
    .B1(_05772_),
    .B2(_05885_),
    .X(_05886_));
 sky130_fd_sc_hd__o22a_1 _21767_ (.A1(_05748_),
    .A2(_05749_),
    .B1(_05721_),
    .B2(_05750_),
    .X(_05887_));
 sky130_fd_sc_hd__or2_1 _21768_ (.A(_05770_),
    .B(_05887_),
    .X(_05888_));
 sky130_fd_sc_hd__a21bo_1 _21769_ (.A1(_05770_),
    .A2(_05887_),
    .B1_N(_05888_),
    .X(_05889_));
 sky130_fd_sc_hd__a2bb2o_1 _21770_ (.A1_N(_05886_),
    .A2_N(_05889_),
    .B1(_05886_),
    .B2(_05889_),
    .X(_05890_));
 sky130_fd_sc_hd__o22a_1 _21771_ (.A1(_05697_),
    .A2(_05773_),
    .B1(_05774_),
    .B2(_05777_),
    .X(_05891_));
 sky130_fd_sc_hd__a2bb2o_1 _21772_ (.A1_N(_05890_),
    .A2_N(_05891_),
    .B1(_05890_),
    .B2(_05891_),
    .X(_05892_));
 sky130_fd_sc_hd__a2bb2o_1 _21773_ (.A1_N(_05776_),
    .A2_N(_05892_),
    .B1(_05776_),
    .B2(_05892_),
    .X(_05893_));
 sky130_fd_sc_hd__o22a_1 _21774_ (.A1(_05778_),
    .A2(_05779_),
    .B1(_05643_),
    .B2(_05780_),
    .X(_05894_));
 sky130_fd_sc_hd__a2bb2o_1 _21775_ (.A1_N(_05893_),
    .A2_N(_05894_),
    .B1(_05893_),
    .B2(_05894_),
    .X(_05895_));
 sky130_fd_sc_hd__a2bb2oi_2 _21776_ (.A1_N(_05785_),
    .A2_N(_05895_),
    .B1(_05785_),
    .B2(_05895_),
    .Y(_02632_));
 sky130_fd_sc_hd__o22a_1 _21777_ (.A1(_05854_),
    .A2(_05855_),
    .B1(_05815_),
    .B2(_05856_),
    .X(_05896_));
 sky130_fd_sc_hd__or2_1 _21778_ (.A(_05882_),
    .B(_05896_),
    .X(_05897_));
 sky130_fd_sc_hd__a21bo_1 _21779_ (.A1(_05882_),
    .A2(_05896_),
    .B1_N(_05897_),
    .X(_05898_));
 sky130_fd_sc_hd__clkbuf_2 _21780_ (.A(_05508_),
    .X(_05899_));
 sky130_fd_sc_hd__buf_2 _21781_ (.A(_05899_),
    .X(_05900_));
 sky130_fd_sc_hd__or2_1 _21782_ (.A(_05535_),
    .B(_05900_),
    .X(_05901_));
 sky130_fd_sc_hd__buf_1 _21783_ (.A(_05683_),
    .X(_05902_));
 sky130_fd_sc_hd__o22a_1 _21784_ (.A1(_05713_),
    .A2(_05902_),
    .B1(_05586_),
    .B2(_05798_),
    .X(_05903_));
 sky130_fd_sc_hd__buf_1 _21785_ (.A(_13611_),
    .X(_05904_));
 sky130_fd_sc_hd__and4_1 _21786_ (.A(_13135_),
    .B(_05808_),
    .C(_13141_),
    .D(_05904_),
    .X(_05905_));
 sky130_fd_sc_hd__or2_1 _21787_ (.A(_05903_),
    .B(_05905_),
    .X(_05906_));
 sky130_fd_sc_hd__a2bb2o_1 _21788_ (.A1_N(_05901_),
    .A2_N(_05906_),
    .B1(_05901_),
    .B2(_05906_),
    .X(_05907_));
 sky130_fd_sc_hd__buf_1 _21789_ (.A(_05343_),
    .X(_05908_));
 sky130_fd_sc_hd__or2_1 _21790_ (.A(_05790_),
    .B(_05908_),
    .X(_05909_));
 sky130_fd_sc_hd__clkbuf_2 _21791_ (.A(_05317_),
    .X(_05910_));
 sky130_vsdinv _21792_ (.A(\pcpi_mul.rs2[14] ),
    .Y(_05911_));
 sky130_fd_sc_hd__clkbuf_2 _21793_ (.A(_05911_),
    .X(_05912_));
 sky130_fd_sc_hd__o22a_1 _21794_ (.A1(_05787_),
    .A2(_05910_),
    .B1(_05912_),
    .B2(_05148_),
    .X(_05913_));
 sky130_fd_sc_hd__clkbuf_2 _21795_ (.A(_13131_),
    .X(_05914_));
 sky130_fd_sc_hd__clkbuf_2 _21796_ (.A(_05647_),
    .X(_05915_));
 sky130_fd_sc_hd__buf_1 _21797_ (.A(_13128_),
    .X(_05916_));
 sky130_fd_sc_hd__buf_1 _21798_ (.A(_13625_),
    .X(_05917_));
 sky130_fd_sc_hd__and4_1 _21799_ (.A(_05914_),
    .B(_05915_),
    .C(_05916_),
    .D(_05917_),
    .X(_05918_));
 sky130_fd_sc_hd__or2_1 _21800_ (.A(_05913_),
    .B(_05918_),
    .X(_05919_));
 sky130_fd_sc_hd__a2bb2o_1 _21801_ (.A1_N(_05909_),
    .A2_N(_05919_),
    .B1(_05909_),
    .B2(_05919_),
    .X(_05920_));
 sky130_fd_sc_hd__a2bb2o_1 _21802_ (.A1_N(_05795_),
    .A2_N(_05920_),
    .B1(_05795_),
    .B2(_05920_),
    .X(_05921_));
 sky130_fd_sc_hd__a2bb2o_1 _21803_ (.A1_N(_05907_),
    .A2_N(_05921_),
    .B1(_05907_),
    .B2(_05921_),
    .X(_05922_));
 sky130_fd_sc_hd__o22a_1 _21804_ (.A1(_05765_),
    .A2(_05879_),
    .B1(_05857_),
    .B2(_05880_),
    .X(_05923_));
 sky130_fd_sc_hd__a21oi_4 _21805_ (.A1(_05826_),
    .A2(_05832_),
    .B1(_05825_),
    .Y(_05924_));
 sky130_fd_sc_hd__clkbuf_2 _21806_ (.A(_05322_),
    .X(_05925_));
 sky130_fd_sc_hd__buf_1 _21807_ (.A(_05734_),
    .X(_05926_));
 sky130_fd_sc_hd__buf_1 _21808_ (.A(_05926_),
    .X(_05927_));
 sky130_fd_sc_hd__buf_2 _21809_ (.A(_05927_),
    .X(_05928_));
 sky130_fd_sc_hd__clkbuf_2 _21810_ (.A(_05305_),
    .X(_05929_));
 sky130_fd_sc_hd__buf_1 _21811_ (.A(_05835_),
    .X(_05930_));
 sky130_fd_sc_hd__buf_1 _21812_ (.A(_05930_),
    .X(_05931_));
 sky130_fd_sc_hd__buf_2 _21813_ (.A(_05931_),
    .X(_05932_));
 sky130_fd_sc_hd__o22a_1 _21814_ (.A1(_05925_),
    .A2(_05928_),
    .B1(_05929_),
    .B2(_05932_),
    .X(_05933_));
 sky130_fd_sc_hd__buf_1 _21815_ (.A(_13173_),
    .X(_05934_));
 sky130_fd_sc_hd__buf_1 _21816_ (.A(_13178_),
    .X(_05935_));
 sky130_fd_sc_hd__and4_2 _21817_ (.A(_05934_),
    .B(_13583_),
    .C(_05935_),
    .D(_13580_),
    .X(_05936_));
 sky130_fd_sc_hd__nor2_2 _21818_ (.A(_05933_),
    .B(_05936_),
    .Y(_05937_));
 sky130_fd_sc_hd__clkbuf_4 _21819_ (.A(_05661_),
    .X(_05938_));
 sky130_fd_sc_hd__nor2_4 _21820_ (.A(_05938_),
    .B(_05818_),
    .Y(_05939_));
 sky130_fd_sc_hd__a2bb2o_2 _21821_ (.A1_N(_05937_),
    .A2_N(_05939_),
    .B1(_05937_),
    .B2(_05939_),
    .X(_05940_));
 sky130_fd_sc_hd__clkbuf_4 _21822_ (.A(_05140_),
    .X(_05941_));
 sky130_vsdinv _21823_ (.A(\pcpi_mul.rs1[14] ),
    .Y(_05942_));
 sky130_fd_sc_hd__buf_1 _21824_ (.A(_05942_),
    .X(_05943_));
 sky130_fd_sc_hd__buf_2 _21825_ (.A(_05943_),
    .X(_05944_));
 sky130_fd_sc_hd__or2_2 _21826_ (.A(_05941_),
    .B(_05944_),
    .X(_05945_));
 sky130_fd_sc_hd__clkbuf_2 _21827_ (.A(_05657_),
    .X(_05946_));
 sky130_fd_sc_hd__clkbuf_2 _21828_ (.A(_05658_),
    .X(_05947_));
 sky130_fd_sc_hd__o22a_1 _21829_ (.A1(_05839_),
    .A2(_05946_),
    .B1(_05842_),
    .B2(_05947_),
    .X(_05948_));
 sky130_fd_sc_hd__buf_1 _21830_ (.A(_05655_),
    .X(_05949_));
 sky130_fd_sc_hd__and4_1 _21831_ (.A(_13160_),
    .B(_05848_),
    .C(_13166_),
    .D(_05949_),
    .X(_05950_));
 sky130_fd_sc_hd__or2_1 _21832_ (.A(_05948_),
    .B(_05950_),
    .X(_05951_));
 sky130_fd_sc_hd__a2bb2o_1 _21833_ (.A1_N(_05945_),
    .A2_N(_05951_),
    .B1(_05945_),
    .B2(_05951_),
    .X(_05952_));
 sky130_fd_sc_hd__o21ba_1 _21834_ (.A1(_05838_),
    .A2(_05850_),
    .B1_N(_05849_),
    .X(_05953_));
 sky130_fd_sc_hd__a2bb2o_1 _21835_ (.A1_N(_05952_),
    .A2_N(_05953_),
    .B1(_05952_),
    .B2(_05953_),
    .X(_05954_));
 sky130_fd_sc_hd__a2bb2o_1 _21836_ (.A1_N(_05940_),
    .A2_N(_05954_),
    .B1(_05940_),
    .B2(_05954_),
    .X(_05955_));
 sky130_fd_sc_hd__o22a_1 _21837_ (.A1(_05851_),
    .A2(_05852_),
    .B1(_05833_),
    .B2(_05853_),
    .X(_05956_));
 sky130_fd_sc_hd__a2bb2o_1 _21838_ (.A1_N(_05955_),
    .A2_N(_05956_),
    .B1(_05955_),
    .B2(_05956_),
    .X(_05957_));
 sky130_fd_sc_hd__a2bb2o_2 _21839_ (.A1_N(_05924_),
    .A2_N(_05957_),
    .B1(_05924_),
    .B2(_05957_),
    .X(_05958_));
 sky130_fd_sc_hd__o22a_1 _21840_ (.A1(_05860_),
    .A2(_05875_),
    .B1(_05859_),
    .B2(_05876_),
    .X(_05959_));
 sky130_fd_sc_hd__o21ba_1 _21841_ (.A1(_05863_),
    .A2(_05874_),
    .B1_N(_05873_),
    .X(_05960_));
 sky130_fd_sc_hd__o21ba_1 _21842_ (.A1(_05800_),
    .A2(_05810_),
    .B1_N(_05809_),
    .X(_05961_));
 sky130_fd_sc_hd__buf_1 _21843_ (.A(_05422_),
    .X(_05962_));
 sky130_fd_sc_hd__clkbuf_2 _21844_ (.A(_05840_),
    .X(_05963_));
 sky130_fd_sc_hd__or2_1 _21845_ (.A(_05962_),
    .B(_05963_),
    .X(_05964_));
 sky130_fd_sc_hd__clkbuf_2 _21846_ (.A(_05864_),
    .X(_05965_));
 sky130_fd_sc_hd__clkbuf_2 _21847_ (.A(_05456_),
    .X(_05966_));
 sky130_fd_sc_hd__buf_1 _21848_ (.A(_05600_),
    .X(_05967_));
 sky130_fd_sc_hd__o22a_1 _21849_ (.A1(_05965_),
    .A2(_05755_),
    .B1(_05966_),
    .B2(_05967_),
    .X(_05968_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _21850_ (.A(_13601_),
    .X(_05969_));
 sky130_fd_sc_hd__and4_1 _21851_ (.A(_13147_),
    .B(_05969_),
    .C(_13153_),
    .D(_13597_),
    .X(_05970_));
 sky130_fd_sc_hd__or2_1 _21852_ (.A(_05968_),
    .B(_05970_),
    .X(_05971_));
 sky130_fd_sc_hd__a2bb2o_1 _21853_ (.A1_N(_05964_),
    .A2_N(_05971_),
    .B1(_05964_),
    .B2(_05971_),
    .X(_05972_));
 sky130_fd_sc_hd__a2bb2o_1 _21854_ (.A1_N(_05961_),
    .A2_N(_05972_),
    .B1(_05961_),
    .B2(_05972_),
    .X(_05973_));
 sky130_fd_sc_hd__a2bb2o_1 _21855_ (.A1_N(_05960_),
    .A2_N(_05973_),
    .B1(_05960_),
    .B2(_05973_),
    .X(_05974_));
 sky130_fd_sc_hd__a2bb2o_1 _21856_ (.A1_N(_05812_),
    .A2_N(_05974_),
    .B1(_05812_),
    .B2(_05974_),
    .X(_05975_));
 sky130_fd_sc_hd__a2bb2o_1 _21857_ (.A1_N(_05959_),
    .A2_N(_05975_),
    .B1(_05959_),
    .B2(_05975_),
    .X(_05976_));
 sky130_fd_sc_hd__o22a_1 _21858_ (.A1(_05719_),
    .A2(_05877_),
    .B1(_05858_),
    .B2(_05878_),
    .X(_05977_));
 sky130_fd_sc_hd__a2bb2o_1 _21859_ (.A1_N(_05976_),
    .A2_N(_05977_),
    .B1(_05976_),
    .B2(_05977_),
    .X(_05978_));
 sky130_fd_sc_hd__a2bb2o_1 _21860_ (.A1_N(_05958_),
    .A2_N(_05978_),
    .B1(_05958_),
    .B2(_05978_),
    .X(_05979_));
 sky130_fd_sc_hd__or2_1 _21861_ (.A(_05923_),
    .B(_05979_),
    .X(_05980_));
 sky130_fd_sc_hd__a21bo_1 _21862_ (.A1(_05923_),
    .A2(_05979_),
    .B1_N(_05980_),
    .X(_05981_));
 sky130_fd_sc_hd__or2_1 _21863_ (.A(_05922_),
    .B(_05981_),
    .X(_05982_));
 sky130_fd_sc_hd__a21bo_1 _21864_ (.A1(_05922_),
    .A2(_05981_),
    .B1_N(_05982_),
    .X(_05983_));
 sky130_fd_sc_hd__a2bb2o_1 _21865_ (.A1_N(_05884_),
    .A2_N(_05983_),
    .B1(_05884_),
    .B2(_05983_),
    .X(_05984_));
 sky130_fd_sc_hd__a2bb2o_1 _21866_ (.A1_N(_05898_),
    .A2_N(_05984_),
    .B1(_05898_),
    .B2(_05984_),
    .X(_05985_));
 sky130_fd_sc_hd__o22a_1 _21867_ (.A1(_05772_),
    .A2(_05885_),
    .B1(_05886_),
    .B2(_05889_),
    .X(_05986_));
 sky130_fd_sc_hd__a2bb2o_1 _21868_ (.A1_N(_05985_),
    .A2_N(_05986_),
    .B1(_05985_),
    .B2(_05986_),
    .X(_05987_));
 sky130_fd_sc_hd__a2bb2o_1 _21869_ (.A1_N(_05888_),
    .A2_N(_05987_),
    .B1(_05888_),
    .B2(_05987_),
    .X(_05988_));
 sky130_fd_sc_hd__o22a_1 _21870_ (.A1(_05890_),
    .A2(_05891_),
    .B1(_05776_),
    .B2(_05892_),
    .X(_05989_));
 sky130_fd_sc_hd__a2bb2o_2 _21871_ (.A1_N(_05988_),
    .A2_N(_05989_),
    .B1(_05988_),
    .B2(_05989_),
    .X(_05990_));
 sky130_fd_sc_hd__o22a_2 _21872_ (.A1(_05893_),
    .A2(_05894_),
    .B1(_05785_),
    .B2(_05895_),
    .X(_05991_));
 sky130_fd_sc_hd__a2bb2oi_4 _21873_ (.A1_N(_05990_),
    .A2_N(_05991_),
    .B1(_05990_),
    .B2(_05991_),
    .Y(_02633_));
 sky130_fd_sc_hd__o22a_2 _21874_ (.A1(_05988_),
    .A2(_05989_),
    .B1(_05990_),
    .B2(_05991_),
    .X(_05992_));
 sky130_fd_sc_hd__o22a_2 _21875_ (.A1(_05955_),
    .A2(_05956_),
    .B1(_05924_),
    .B2(_05957_),
    .X(_05993_));
 sky130_fd_sc_hd__or2_1 _21876_ (.A(_05980_),
    .B(_05993_),
    .X(_05994_));
 sky130_fd_sc_hd__a21bo_1 _21877_ (.A1(_05980_),
    .A2(_05993_),
    .B1_N(_05994_),
    .X(_05995_));
 sky130_vsdinv _21878_ (.A(\pcpi_mul.rs2[15] ),
    .Y(_05996_));
 sky130_fd_sc_hd__buf_1 _21879_ (.A(_05996_),
    .X(_05997_));
 sky130_fd_sc_hd__buf_4 _21880_ (.A(_05997_),
    .X(_05998_));
 sky130_fd_sc_hd__buf_2 _21881_ (.A(_05998_),
    .X(_05999_));
 sky130_fd_sc_hd__buf_2 _21882_ (.A(_05999_),
    .X(_06000_));
 sky130_fd_sc_hd__buf_4 _21883_ (.A(_06000_),
    .X(_06001_));
 sky130_fd_sc_hd__or2_4 _21884_ (.A(_06001_),
    .B(_05590_),
    .X(_06002_));
 sky130_fd_sc_hd__clkbuf_2 _21885_ (.A(_05755_),
    .X(_06003_));
 sky130_fd_sc_hd__or2_1 _21886_ (.A(_05797_),
    .B(_06003_),
    .X(_06004_));
 sky130_fd_sc_hd__clkbuf_2 _21887_ (.A(_05369_),
    .X(_06005_));
 sky130_fd_sc_hd__o22a_1 _21888_ (.A1(_05713_),
    .A2(_06005_),
    .B1(_05586_),
    .B2(_05899_),
    .X(_06006_));
 sky130_fd_sc_hd__buf_1 _21889_ (.A(_13607_),
    .X(_06007_));
 sky130_fd_sc_hd__and4_1 _21890_ (.A(_05805_),
    .B(_05904_),
    .C(_05807_),
    .D(_06007_),
    .X(_06008_));
 sky130_fd_sc_hd__or2_1 _21891_ (.A(_06006_),
    .B(_06008_),
    .X(_06009_));
 sky130_fd_sc_hd__a2bb2o_1 _21892_ (.A1_N(_06004_),
    .A2_N(_06009_),
    .B1(_06004_),
    .B2(_06009_),
    .X(_06010_));
 sky130_fd_sc_hd__clkbuf_2 _21893_ (.A(_05902_),
    .X(_06011_));
 sky130_fd_sc_hd__or2_1 _21894_ (.A(_05790_),
    .B(_06011_),
    .X(_06012_));
 sky130_fd_sc_hd__clkbuf_2 _21895_ (.A(_05911_),
    .X(_06013_));
 sky130_fd_sc_hd__clkbuf_2 _21896_ (.A(_05786_),
    .X(_06014_));
 sky130_fd_sc_hd__clkbuf_2 _21897_ (.A(_05314_),
    .X(_06015_));
 sky130_fd_sc_hd__o22a_1 _21898_ (.A1(_06013_),
    .A2(_05380_),
    .B1(_06014_),
    .B2(_06015_),
    .X(_06016_));
 sky130_fd_sc_hd__buf_1 _21899_ (.A(_13131_),
    .X(_06017_));
 sky130_fd_sc_hd__and4_1 _21900_ (.A(_05916_),
    .B(_05915_),
    .C(_06017_),
    .D(_05806_),
    .X(_06018_));
 sky130_fd_sc_hd__or2_1 _21901_ (.A(_06016_),
    .B(_06018_),
    .X(_06019_));
 sky130_fd_sc_hd__a2bb2o_1 _21902_ (.A1_N(_06012_),
    .A2_N(_06019_),
    .B1(_06012_),
    .B2(_06019_),
    .X(_06020_));
 sky130_fd_sc_hd__o21ba_1 _21903_ (.A1(_05909_),
    .A2(_05919_),
    .B1_N(_05918_),
    .X(_06021_));
 sky130_fd_sc_hd__a2bb2o_1 _21904_ (.A1_N(_06020_),
    .A2_N(_06021_),
    .B1(_06020_),
    .B2(_06021_),
    .X(_06022_));
 sky130_fd_sc_hd__a2bb2o_1 _21905_ (.A1_N(_06010_),
    .A2_N(_06022_),
    .B1(_06010_),
    .B2(_06022_),
    .X(_06023_));
 sky130_fd_sc_hd__nor2_2 _21906_ (.A(_06002_),
    .B(_06023_),
    .Y(_06024_));
 sky130_fd_sc_hd__a21oi_2 _21907_ (.A1(_06002_),
    .A2(_06023_),
    .B1(_06024_),
    .Y(_06025_));
 sky130_fd_sc_hd__o22a_1 _21908_ (.A1(_05976_),
    .A2(_05977_),
    .B1(_05958_),
    .B2(_05978_),
    .X(_06026_));
 sky130_fd_sc_hd__a21oi_4 _21909_ (.A1(_05937_),
    .A2(_05939_),
    .B1(_05936_),
    .Y(_06027_));
 sky130_fd_sc_hd__clkbuf_2 _21910_ (.A(_05930_),
    .X(_06028_));
 sky130_fd_sc_hd__clkbuf_2 _21911_ (.A(_06028_),
    .X(_06029_));
 sky130_fd_sc_hd__buf_1 _21912_ (.A(_05942_),
    .X(_06030_));
 sky130_fd_sc_hd__buf_1 _21913_ (.A(_06030_),
    .X(_06031_));
 sky130_fd_sc_hd__clkbuf_4 _21914_ (.A(_06031_),
    .X(_06032_));
 sky130_fd_sc_hd__o22a_2 _21915_ (.A1(_05925_),
    .A2(_06029_),
    .B1(_05306_),
    .B2(_06032_),
    .X(_06033_));
 sky130_fd_sc_hd__and4_2 _21916_ (.A(_05934_),
    .B(_13580_),
    .C(_05935_),
    .D(_13576_),
    .X(_06034_));
 sky130_fd_sc_hd__nor2_2 _21917_ (.A(_06033_),
    .B(_06034_),
    .Y(_06035_));
 sky130_fd_sc_hd__nor2_4 _21918_ (.A(_05827_),
    .B(_05821_),
    .Y(_06036_));
 sky130_fd_sc_hd__a2bb2o_1 _21919_ (.A1_N(_06035_),
    .A2_N(_06036_),
    .B1(_06035_),
    .B2(_06036_),
    .X(_06037_));
 sky130_vsdinv _21920_ (.A(\pcpi_mul.rs1[15] ),
    .Y(_06038_));
 sky130_fd_sc_hd__buf_1 _21921_ (.A(_06038_),
    .X(_06039_));
 sky130_fd_sc_hd__clkbuf_2 _21922_ (.A(_06039_),
    .X(_06040_));
 sky130_fd_sc_hd__or2_2 _21923_ (.A(_05941_),
    .B(_06040_),
    .X(_06041_));
 sky130_fd_sc_hd__clkbuf_2 _21924_ (.A(_05658_),
    .X(_06042_));
 sky130_fd_sc_hd__clkbuf_2 _21925_ (.A(_05666_),
    .X(_06043_));
 sky130_fd_sc_hd__o22a_1 _21926_ (.A1(_05737_),
    .A2(_06042_),
    .B1(_05739_),
    .B2(_06043_),
    .X(_06044_));
 sky130_fd_sc_hd__and4_1 _21927_ (.A(_13160_),
    .B(_05949_),
    .C(_13166_),
    .D(_13584_),
    .X(_06045_));
 sky130_fd_sc_hd__or2_1 _21928_ (.A(_06044_),
    .B(_06045_),
    .X(_06046_));
 sky130_fd_sc_hd__a2bb2o_1 _21929_ (.A1_N(_06041_),
    .A2_N(_06046_),
    .B1(_06041_),
    .B2(_06046_),
    .X(_06047_));
 sky130_fd_sc_hd__o21ba_1 _21930_ (.A1(_05945_),
    .A2(_05951_),
    .B1_N(_05950_),
    .X(_06048_));
 sky130_fd_sc_hd__a2bb2o_1 _21931_ (.A1_N(_06047_),
    .A2_N(_06048_),
    .B1(_06047_),
    .B2(_06048_),
    .X(_06049_));
 sky130_fd_sc_hd__a2bb2o_1 _21932_ (.A1_N(_06037_),
    .A2_N(_06049_),
    .B1(_06037_),
    .B2(_06049_),
    .X(_06050_));
 sky130_fd_sc_hd__o22a_1 _21933_ (.A1(_05952_),
    .A2(_05953_),
    .B1(_05940_),
    .B2(_05954_),
    .X(_06051_));
 sky130_fd_sc_hd__a2bb2o_1 _21934_ (.A1_N(_06050_),
    .A2_N(_06051_),
    .B1(_06050_),
    .B2(_06051_),
    .X(_06052_));
 sky130_fd_sc_hd__a2bb2o_1 _21935_ (.A1_N(_06027_),
    .A2_N(_06052_),
    .B1(_06027_),
    .B2(_06052_),
    .X(_06053_));
 sky130_fd_sc_hd__o22a_1 _21936_ (.A1(_05961_),
    .A2(_05972_),
    .B1(_05960_),
    .B2(_05973_),
    .X(_06054_));
 sky130_fd_sc_hd__o22a_1 _21937_ (.A1(_05795_),
    .A2(_05920_),
    .B1(_05907_),
    .B2(_05921_),
    .X(_06055_));
 sky130_fd_sc_hd__o21ba_1 _21938_ (.A1(_05964_),
    .A2(_05971_),
    .B1_N(_05970_),
    .X(_06056_));
 sky130_fd_sc_hd__o21ba_1 _21939_ (.A1(_05901_),
    .A2(_05906_),
    .B1_N(_05905_),
    .X(_06057_));
 sky130_fd_sc_hd__or2_2 _21940_ (.A(_05962_),
    .B(_05730_),
    .X(_06058_));
 sky130_fd_sc_hd__o22a_1 _21941_ (.A1(_05864_),
    .A2(_05738_),
    .B1(_05966_),
    .B2(_05662_),
    .X(_06059_));
 sky130_fd_sc_hd__and4_1 _21942_ (.A(_13147_),
    .B(_13597_),
    .C(_13153_),
    .D(_05742_),
    .X(_06060_));
 sky130_fd_sc_hd__or2_1 _21943_ (.A(_06059_),
    .B(_06060_),
    .X(_06061_));
 sky130_fd_sc_hd__a2bb2o_1 _21944_ (.A1_N(_06058_),
    .A2_N(_06061_),
    .B1(_06058_),
    .B2(_06061_),
    .X(_06062_));
 sky130_fd_sc_hd__a2bb2o_1 _21945_ (.A1_N(_06057_),
    .A2_N(_06062_),
    .B1(_06057_),
    .B2(_06062_),
    .X(_06063_));
 sky130_fd_sc_hd__a2bb2o_1 _21946_ (.A1_N(_06056_),
    .A2_N(_06063_),
    .B1(_06056_),
    .B2(_06063_),
    .X(_06064_));
 sky130_fd_sc_hd__a2bb2o_1 _21947_ (.A1_N(_06055_),
    .A2_N(_06064_),
    .B1(_06055_),
    .B2(_06064_),
    .X(_06065_));
 sky130_fd_sc_hd__a2bb2o_1 _21948_ (.A1_N(_06054_),
    .A2_N(_06065_),
    .B1(_06054_),
    .B2(_06065_),
    .X(_06066_));
 sky130_fd_sc_hd__o22a_1 _21949_ (.A1(_05812_),
    .A2(_05974_),
    .B1(_05959_),
    .B2(_05975_),
    .X(_06067_));
 sky130_fd_sc_hd__a2bb2o_1 _21950_ (.A1_N(_06066_),
    .A2_N(_06067_),
    .B1(_06066_),
    .B2(_06067_),
    .X(_06068_));
 sky130_fd_sc_hd__a2bb2o_1 _21951_ (.A1_N(_06053_),
    .A2_N(_06068_),
    .B1(_06053_),
    .B2(_06068_),
    .X(_06069_));
 sky130_fd_sc_hd__or2_1 _21952_ (.A(_06026_),
    .B(_06069_),
    .X(_06070_));
 sky130_fd_sc_hd__a21boi_1 _21953_ (.A1(_06026_),
    .A2(_06069_),
    .B1_N(_06070_),
    .Y(_06071_));
 sky130_fd_sc_hd__nand2_1 _21954_ (.A(_06025_),
    .B(_06071_),
    .Y(_06072_));
 sky130_fd_sc_hd__o21ai_1 _21955_ (.A1(_06025_),
    .A2(_06071_),
    .B1(_06072_),
    .Y(_06073_));
 sky130_fd_sc_hd__a2bb2o_1 _21956_ (.A1_N(_05982_),
    .A2_N(_06073_),
    .B1(_05982_),
    .B2(_06073_),
    .X(_06074_));
 sky130_fd_sc_hd__a2bb2o_1 _21957_ (.A1_N(_05995_),
    .A2_N(_06074_),
    .B1(_05995_),
    .B2(_06074_),
    .X(_06075_));
 sky130_fd_sc_hd__o22a_1 _21958_ (.A1(_05884_),
    .A2(_05983_),
    .B1(_05898_),
    .B2(_05984_),
    .X(_06076_));
 sky130_fd_sc_hd__a2bb2o_1 _21959_ (.A1_N(_06075_),
    .A2_N(_06076_),
    .B1(_06075_),
    .B2(_06076_),
    .X(_06077_));
 sky130_fd_sc_hd__a2bb2o_1 _21960_ (.A1_N(_05897_),
    .A2_N(_06077_),
    .B1(_05897_),
    .B2(_06077_),
    .X(_06078_));
 sky130_fd_sc_hd__o22a_1 _21961_ (.A1(_05985_),
    .A2(_05986_),
    .B1(_05888_),
    .B2(_05987_),
    .X(_06079_));
 sky130_fd_sc_hd__a2bb2o_2 _21962_ (.A1_N(_06078_),
    .A2_N(_06079_),
    .B1(_06078_),
    .B2(_06079_),
    .X(_06080_));
 sky130_fd_sc_hd__a2bb2oi_4 _21963_ (.A1_N(_05992_),
    .A2_N(_06080_),
    .B1(_05992_),
    .B2(_06080_),
    .Y(_02634_));
 sky130_fd_sc_hd__o22a_1 _21964_ (.A1(_06078_),
    .A2(_06079_),
    .B1(_05992_),
    .B2(_06080_),
    .X(_06081_));
 sky130_fd_sc_hd__buf_2 _21965_ (.A(_06081_),
    .X(_06082_));
 sky130_fd_sc_hd__o22a_1 _21966_ (.A1(_06050_),
    .A2(_06051_),
    .B1(_06027_),
    .B2(_06052_),
    .X(_06083_));
 sky130_fd_sc_hd__or2_1 _21967_ (.A(_06070_),
    .B(_06083_),
    .X(_06084_));
 sky130_fd_sc_hd__a21bo_1 _21968_ (.A1(_06070_),
    .A2(_06083_),
    .B1_N(_06084_),
    .X(_06085_));
 sky130_vsdinv _21969_ (.A(\pcpi_mul.rs2[16] ),
    .Y(_06086_));
 sky130_fd_sc_hd__buf_1 _21970_ (.A(_06086_),
    .X(_06087_));
 sky130_fd_sc_hd__buf_2 _21971_ (.A(_06087_),
    .X(_06088_));
 sky130_fd_sc_hd__clkbuf_2 _21972_ (.A(_06088_),
    .X(_06089_));
 sky130_fd_sc_hd__clkbuf_4 _21973_ (.A(_06089_),
    .X(_06090_));
 sky130_fd_sc_hd__o22a_2 _21974_ (.A1(_06090_),
    .A2(_05152_),
    .B1(_06001_),
    .B2(_05299_),
    .X(_06091_));
 sky130_fd_sc_hd__clkbuf_2 _21975_ (.A(_06087_),
    .X(_06092_));
 sky130_fd_sc_hd__clkbuf_4 _21976_ (.A(_06092_),
    .X(_06093_));
 sky130_fd_sc_hd__clkbuf_4 _21977_ (.A(_06093_),
    .X(_06094_));
 sky130_fd_sc_hd__buf_1 _21978_ (.A(_05996_),
    .X(_06095_));
 sky130_fd_sc_hd__buf_2 _21979_ (.A(_06095_),
    .X(_06096_));
 sky130_fd_sc_hd__or4_4 _21980_ (.A(_06094_),
    .B(_05459_),
    .C(_06096_),
    .D(_05792_),
    .X(_06097_));
 sky130_fd_sc_hd__or2b_2 _21981_ (.A(_06091_),
    .B_N(_06097_),
    .X(_06098_));
 sky130_fd_sc_hd__clkbuf_2 _21982_ (.A(_05738_),
    .X(_06099_));
 sky130_fd_sc_hd__or2_1 _21983_ (.A(_05536_),
    .B(_06099_),
    .X(_06100_));
 sky130_fd_sc_hd__buf_2 _21984_ (.A(_05556_),
    .X(_06101_));
 sky130_fd_sc_hd__o22a_1 _21985_ (.A1(_05801_),
    .A2(_05899_),
    .B1(_05587_),
    .B2(_06101_),
    .X(_06102_));
 sky130_fd_sc_hd__clkbuf_2 _21986_ (.A(_13135_),
    .X(_06103_));
 sky130_fd_sc_hd__clkbuf_2 _21987_ (.A(_13141_),
    .X(_06104_));
 sky130_fd_sc_hd__and4_1 _21988_ (.A(_06103_),
    .B(_06007_),
    .C(_06104_),
    .D(_13603_),
    .X(_06105_));
 sky130_fd_sc_hd__or2_1 _21989_ (.A(_06102_),
    .B(_06105_),
    .X(_06106_));
 sky130_fd_sc_hd__a2bb2o_1 _21990_ (.A1_N(_06100_),
    .A2_N(_06106_),
    .B1(_06100_),
    .B2(_06106_),
    .X(_06107_));
 sky130_fd_sc_hd__clkbuf_2 _21991_ (.A(_05707_),
    .X(_06108_));
 sky130_fd_sc_hd__or2_1 _21992_ (.A(_06108_),
    .B(_05799_),
    .X(_06109_));
 sky130_fd_sc_hd__clkbuf_2 _21993_ (.A(_05911_),
    .X(_06110_));
 sky130_fd_sc_hd__clkbuf_2 _21994_ (.A(_05787_),
    .X(_06111_));
 sky130_fd_sc_hd__clkbuf_2 _21995_ (.A(_05338_),
    .X(_06112_));
 sky130_fd_sc_hd__o22a_1 _21996_ (.A1(_06110_),
    .A2(_06015_),
    .B1(_06111_),
    .B2(_06112_),
    .X(_06113_));
 sky130_fd_sc_hd__clkbuf_2 _21997_ (.A(_13128_),
    .X(_06114_));
 sky130_fd_sc_hd__clkbuf_2 _21998_ (.A(_13619_),
    .X(_06115_));
 sky130_fd_sc_hd__clkbuf_2 _21999_ (.A(_13615_),
    .X(_06116_));
 sky130_fd_sc_hd__and4_1 _22000_ (.A(_06114_),
    .B(_06115_),
    .C(_05914_),
    .D(_06116_),
    .X(_06117_));
 sky130_fd_sc_hd__or2_1 _22001_ (.A(_06113_),
    .B(_06117_),
    .X(_06118_));
 sky130_fd_sc_hd__a2bb2o_1 _22002_ (.A1_N(_06109_),
    .A2_N(_06118_),
    .B1(_06109_),
    .B2(_06118_),
    .X(_06119_));
 sky130_fd_sc_hd__o21ba_1 _22003_ (.A1(_06012_),
    .A2(_06019_),
    .B1_N(_06018_),
    .X(_06120_));
 sky130_fd_sc_hd__a2bb2o_1 _22004_ (.A1_N(_06119_),
    .A2_N(_06120_),
    .B1(_06119_),
    .B2(_06120_),
    .X(_06121_));
 sky130_fd_sc_hd__a2bb2o_1 _22005_ (.A1_N(_06107_),
    .A2_N(_06121_),
    .B1(_06107_),
    .B2(_06121_),
    .X(_06122_));
 sky130_fd_sc_hd__nor2_2 _22006_ (.A(_06098_),
    .B(_06122_),
    .Y(_06123_));
 sky130_fd_sc_hd__a21oi_2 _22007_ (.A1(_06098_),
    .A2(_06122_),
    .B1(_06123_),
    .Y(_06124_));
 sky130_fd_sc_hd__nand2_1 _22008_ (.A(_06024_),
    .B(_06124_),
    .Y(_06125_));
 sky130_fd_sc_hd__o21ai_1 _22009_ (.A1(_06024_),
    .A2(_06124_),
    .B1(_06125_),
    .Y(_06126_));
 sky130_fd_sc_hd__o22a_1 _22010_ (.A1(_06066_),
    .A2(_06067_),
    .B1(_06053_),
    .B2(_06068_),
    .X(_06127_));
 sky130_fd_sc_hd__a21oi_2 _22011_ (.A1(_06035_),
    .A2(_06036_),
    .B1(_06034_),
    .Y(_06128_));
 sky130_fd_sc_hd__buf_1 _22012_ (.A(_06030_),
    .X(_06129_));
 sky130_fd_sc_hd__clkbuf_2 _22013_ (.A(_06129_),
    .X(_06130_));
 sky130_fd_sc_hd__clkbuf_2 _22014_ (.A(_06039_),
    .X(_06131_));
 sky130_fd_sc_hd__clkbuf_2 _22015_ (.A(_06131_),
    .X(_06132_));
 sky130_fd_sc_hd__o22a_2 _22016_ (.A1(_05925_),
    .A2(_06130_),
    .B1(_05929_),
    .B2(_06132_),
    .X(_06133_));
 sky130_fd_sc_hd__and4_4 _22017_ (.A(_05934_),
    .B(_13576_),
    .C(_05935_),
    .D(_13571_),
    .X(_06134_));
 sky130_fd_sc_hd__nor2_2 _22018_ (.A(_06133_),
    .B(_06134_),
    .Y(_06135_));
 sky130_fd_sc_hd__nor2_4 _22019_ (.A(_05938_),
    .B(_05932_),
    .Y(_06136_));
 sky130_fd_sc_hd__a2bb2o_1 _22020_ (.A1_N(_06135_),
    .A2_N(_06136_),
    .B1(_06135_),
    .B2(_06136_),
    .X(_06137_));
 sky130_vsdinv _22021_ (.A(\pcpi_mul.rs1[16] ),
    .Y(_06138_));
 sky130_fd_sc_hd__buf_1 _22022_ (.A(_06138_),
    .X(_06139_));
 sky130_fd_sc_hd__buf_2 _22023_ (.A(_06139_),
    .X(_06140_));
 sky130_fd_sc_hd__or2_2 _22024_ (.A(_05941_),
    .B(_06140_),
    .X(_06141_));
 sky130_fd_sc_hd__o22a_1 _22025_ (.A1(_05839_),
    .A2(_06043_),
    .B1(_05842_),
    .B2(_05735_),
    .X(_06142_));
 sky130_fd_sc_hd__buf_1 _22026_ (.A(\pcpi_mul.rs1[11] ),
    .X(_06143_));
 sky130_fd_sc_hd__buf_1 _22027_ (.A(_06143_),
    .X(_06144_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _22028_ (.A(\pcpi_mul.rs1[12] ),
    .X(_06145_));
 sky130_fd_sc_hd__and4_1 _22029_ (.A(_05845_),
    .B(_06144_),
    .C(_05847_),
    .D(_06145_),
    .X(_06146_));
 sky130_fd_sc_hd__or2_1 _22030_ (.A(_06142_),
    .B(_06146_),
    .X(_06147_));
 sky130_fd_sc_hd__a2bb2o_1 _22031_ (.A1_N(_06141_),
    .A2_N(_06147_),
    .B1(_06141_),
    .B2(_06147_),
    .X(_06148_));
 sky130_fd_sc_hd__o21ba_1 _22032_ (.A1(_06041_),
    .A2(_06046_),
    .B1_N(_06045_),
    .X(_06149_));
 sky130_fd_sc_hd__a2bb2o_1 _22033_ (.A1_N(_06148_),
    .A2_N(_06149_),
    .B1(_06148_),
    .B2(_06149_),
    .X(_06150_));
 sky130_fd_sc_hd__a2bb2o_1 _22034_ (.A1_N(_06137_),
    .A2_N(_06150_),
    .B1(_06137_),
    .B2(_06150_),
    .X(_06151_));
 sky130_fd_sc_hd__o22a_1 _22035_ (.A1(_06047_),
    .A2(_06048_),
    .B1(_06037_),
    .B2(_06049_),
    .X(_06152_));
 sky130_fd_sc_hd__a2bb2o_1 _22036_ (.A1_N(_06151_),
    .A2_N(_06152_),
    .B1(_06151_),
    .B2(_06152_),
    .X(_06153_));
 sky130_fd_sc_hd__a2bb2o_1 _22037_ (.A1_N(_06128_),
    .A2_N(_06153_),
    .B1(_06128_),
    .B2(_06153_),
    .X(_06154_));
 sky130_fd_sc_hd__o22a_1 _22038_ (.A1(_06057_),
    .A2(_06062_),
    .B1(_06056_),
    .B2(_06063_),
    .X(_06155_));
 sky130_fd_sc_hd__o22a_1 _22039_ (.A1(_06020_),
    .A2(_06021_),
    .B1(_06010_),
    .B2(_06022_),
    .X(_06156_));
 sky130_fd_sc_hd__o21ba_1 _22040_ (.A1(_06058_),
    .A2(_06061_),
    .B1_N(_06060_),
    .X(_06157_));
 sky130_fd_sc_hd__o21ba_1 _22041_ (.A1(_06004_),
    .A2(_06009_),
    .B1_N(_06008_),
    .X(_06158_));
 sky130_fd_sc_hd__or2_1 _22042_ (.A(_05962_),
    .B(_05947_),
    .X(_06159_));
 sky130_fd_sc_hd__o22a_1 _22043_ (.A1(_05965_),
    .A2(_05840_),
    .B1(_05966_),
    .B2(_05729_),
    .X(_06160_));
 sky130_fd_sc_hd__and4_1 _22044_ (.A(_13147_),
    .B(_05742_),
    .C(_13153_),
    .D(_13590_),
    .X(_06161_));
 sky130_fd_sc_hd__or2_1 _22045_ (.A(_06160_),
    .B(_06161_),
    .X(_06162_));
 sky130_fd_sc_hd__a2bb2o_1 _22046_ (.A1_N(_06159_),
    .A2_N(_06162_),
    .B1(_06159_),
    .B2(_06162_),
    .X(_06163_));
 sky130_fd_sc_hd__a2bb2o_1 _22047_ (.A1_N(_06158_),
    .A2_N(_06163_),
    .B1(_06158_),
    .B2(_06163_),
    .X(_06164_));
 sky130_fd_sc_hd__a2bb2o_1 _22048_ (.A1_N(_06157_),
    .A2_N(_06164_),
    .B1(_06157_),
    .B2(_06164_),
    .X(_06165_));
 sky130_fd_sc_hd__a2bb2o_1 _22049_ (.A1_N(_06156_),
    .A2_N(_06165_),
    .B1(_06156_),
    .B2(_06165_),
    .X(_06166_));
 sky130_fd_sc_hd__a2bb2o_1 _22050_ (.A1_N(_06155_),
    .A2_N(_06166_),
    .B1(_06155_),
    .B2(_06166_),
    .X(_06167_));
 sky130_fd_sc_hd__o22a_1 _22051_ (.A1(_06055_),
    .A2(_06064_),
    .B1(_06054_),
    .B2(_06065_),
    .X(_06168_));
 sky130_fd_sc_hd__a2bb2o_1 _22052_ (.A1_N(_06167_),
    .A2_N(_06168_),
    .B1(_06167_),
    .B2(_06168_),
    .X(_06169_));
 sky130_fd_sc_hd__a2bb2o_1 _22053_ (.A1_N(_06154_),
    .A2_N(_06169_),
    .B1(_06154_),
    .B2(_06169_),
    .X(_06170_));
 sky130_fd_sc_hd__or2_1 _22054_ (.A(_06127_),
    .B(_06170_),
    .X(_06171_));
 sky130_fd_sc_hd__a21bo_1 _22055_ (.A1(_06127_),
    .A2(_06170_),
    .B1_N(_06171_),
    .X(_06172_));
 sky130_fd_sc_hd__or2_1 _22056_ (.A(_06126_),
    .B(_06172_),
    .X(_06173_));
 sky130_fd_sc_hd__a21bo_1 _22057_ (.A1(_06126_),
    .A2(_06172_),
    .B1_N(_06173_),
    .X(_06174_));
 sky130_fd_sc_hd__a2bb2o_1 _22058_ (.A1_N(_06072_),
    .A2_N(_06174_),
    .B1(_06072_),
    .B2(_06174_),
    .X(_06175_));
 sky130_fd_sc_hd__a2bb2o_1 _22059_ (.A1_N(_06085_),
    .A2_N(_06175_),
    .B1(_06085_),
    .B2(_06175_),
    .X(_06176_));
 sky130_fd_sc_hd__o22a_1 _22060_ (.A1(_05982_),
    .A2(_06073_),
    .B1(_05995_),
    .B2(_06074_),
    .X(_06177_));
 sky130_fd_sc_hd__a2bb2o_1 _22061_ (.A1_N(_06176_),
    .A2_N(_06177_),
    .B1(_06176_),
    .B2(_06177_),
    .X(_06178_));
 sky130_fd_sc_hd__a2bb2o_1 _22062_ (.A1_N(_05994_),
    .A2_N(_06178_),
    .B1(_05994_),
    .B2(_06178_),
    .X(_06179_));
 sky130_fd_sc_hd__o22a_1 _22063_ (.A1(_06075_),
    .A2(_06076_),
    .B1(_05897_),
    .B2(_06077_),
    .X(_06180_));
 sky130_fd_sc_hd__or2_1 _22064_ (.A(_06179_),
    .B(_06180_),
    .X(_06181_));
 sky130_fd_sc_hd__a21bo_1 _22065_ (.A1(_06179_),
    .A2(_06180_),
    .B1_N(_06181_),
    .X(_06182_));
 sky130_fd_sc_hd__buf_2 _22066_ (.A(_06182_),
    .X(_06183_));
 sky130_fd_sc_hd__a2bb2oi_4 _22067_ (.A1_N(_06082_),
    .A2_N(_06183_),
    .B1(_06082_),
    .B2(_06183_),
    .Y(_02635_));
 sky130_fd_sc_hd__o22a_1 _22068_ (.A1(_06151_),
    .A2(_06152_),
    .B1(_06128_),
    .B2(_06153_),
    .X(_06184_));
 sky130_fd_sc_hd__or2_1 _22069_ (.A(_06171_),
    .B(_06184_),
    .X(_06185_));
 sky130_fd_sc_hd__a21bo_1 _22070_ (.A1(_06171_),
    .A2(_06184_),
    .B1_N(_06185_),
    .X(_06186_));
 sky130_fd_sc_hd__clkbuf_2 _22071_ (.A(_05314_),
    .X(_06187_));
 sky130_fd_sc_hd__or2_1 _22072_ (.A(_05997_),
    .B(_06187_),
    .X(_06188_));
 sky130_vsdinv _22073_ (.A(\pcpi_mul.rs2[17] ),
    .Y(_06189_));
 sky130_fd_sc_hd__o22a_1 _22074_ (.A1(_06086_),
    .A2(_05379_),
    .B1(_06189_),
    .B2(_05146_),
    .X(_06190_));
 sky130_fd_sc_hd__and4_1 _22075_ (.A(_13120_),
    .B(_05647_),
    .C(\pcpi_mul.rs2[17] ),
    .D(_13625_),
    .X(_06191_));
 sky130_fd_sc_hd__or2_1 _22076_ (.A(_06190_),
    .B(_06191_),
    .X(_06192_));
 sky130_fd_sc_hd__a2bb2o_1 _22077_ (.A1_N(_06188_),
    .A2_N(_06192_),
    .B1(_06188_),
    .B2(_06192_),
    .X(_06193_));
 sky130_fd_sc_hd__or2_2 _22078_ (.A(_06097_),
    .B(_06193_),
    .X(_06194_));
 sky130_fd_sc_hd__a21bo_1 _22079_ (.A1(_06097_),
    .A2(_06193_),
    .B1_N(_06194_),
    .X(_06195_));
 sky130_fd_sc_hd__or2_1 _22080_ (.A(_05797_),
    .B(_05663_),
    .X(_06196_));
 sky130_fd_sc_hd__o22a_1 _22081_ (.A1(_05801_),
    .A2(_05755_),
    .B1(_05802_),
    .B2(_05967_),
    .X(_06197_));
 sky130_fd_sc_hd__and4_1 _22082_ (.A(_05805_),
    .B(_05969_),
    .C(_05807_),
    .D(_05741_),
    .X(_06198_));
 sky130_fd_sc_hd__or2_1 _22083_ (.A(_06197_),
    .B(_06198_),
    .X(_06199_));
 sky130_fd_sc_hd__a2bb2o_1 _22084_ (.A1_N(_06196_),
    .A2_N(_06199_),
    .B1(_06196_),
    .B2(_06199_),
    .X(_06200_));
 sky130_fd_sc_hd__clkbuf_2 _22085_ (.A(_05680_),
    .X(_06201_));
 sky130_fd_sc_hd__or2_1 _22086_ (.A(_06108_),
    .B(_06201_),
    .X(_06202_));
 sky130_fd_sc_hd__o22a_1 _22087_ (.A1(_05912_),
    .A2(_05902_),
    .B1(_06014_),
    .B2(_06005_),
    .X(_06203_));
 sky130_fd_sc_hd__buf_1 _22088_ (.A(_05376_),
    .X(_06204_));
 sky130_fd_sc_hd__and4_1 _22089_ (.A(_05916_),
    .B(_06204_),
    .C(_06017_),
    .D(_05904_),
    .X(_06205_));
 sky130_fd_sc_hd__or2_1 _22090_ (.A(_06203_),
    .B(_06205_),
    .X(_06206_));
 sky130_fd_sc_hd__a2bb2o_1 _22091_ (.A1_N(_06202_),
    .A2_N(_06206_),
    .B1(_06202_),
    .B2(_06206_),
    .X(_06207_));
 sky130_fd_sc_hd__o21ba_1 _22092_ (.A1(_06109_),
    .A2(_06118_),
    .B1_N(_06117_),
    .X(_06208_));
 sky130_fd_sc_hd__a2bb2o_1 _22093_ (.A1_N(_06207_),
    .A2_N(_06208_),
    .B1(_06207_),
    .B2(_06208_),
    .X(_06209_));
 sky130_fd_sc_hd__a2bb2o_1 _22094_ (.A1_N(_06200_),
    .A2_N(_06209_),
    .B1(_06200_),
    .B2(_06209_),
    .X(_06210_));
 sky130_fd_sc_hd__nor2_2 _22095_ (.A(_06195_),
    .B(_06210_),
    .Y(_06211_));
 sky130_fd_sc_hd__a21oi_2 _22096_ (.A1(_06195_),
    .A2(_06210_),
    .B1(_06211_),
    .Y(_06212_));
 sky130_fd_sc_hd__nand2_1 _22097_ (.A(_06123_),
    .B(_06212_),
    .Y(_06213_));
 sky130_fd_sc_hd__o21ai_1 _22098_ (.A1(_06123_),
    .A2(_06212_),
    .B1(_06213_),
    .Y(_06214_));
 sky130_fd_sc_hd__o22a_1 _22099_ (.A1(_06167_),
    .A2(_06168_),
    .B1(_06154_),
    .B2(_06169_),
    .X(_06215_));
 sky130_fd_sc_hd__a21oi_2 _22100_ (.A1(_06135_),
    .A2(_06136_),
    .B1(_06134_),
    .Y(_06216_));
 sky130_fd_sc_hd__buf_2 _22101_ (.A(_05323_),
    .X(_06217_));
 sky130_fd_sc_hd__buf_1 _22102_ (.A(_06139_),
    .X(_06218_));
 sky130_fd_sc_hd__clkbuf_4 _22103_ (.A(_06218_),
    .X(_06219_));
 sky130_fd_sc_hd__o22a_1 _22104_ (.A1(_06217_),
    .A2(_06132_),
    .B1(_05307_),
    .B2(_06219_),
    .X(_06220_));
 sky130_fd_sc_hd__and4_2 _22105_ (.A(_13174_),
    .B(_13571_),
    .C(_13179_),
    .D(_13568_),
    .X(_06221_));
 sky130_fd_sc_hd__nor2_1 _22106_ (.A(_06220_),
    .B(_06221_),
    .Y(_06222_));
 sky130_fd_sc_hd__nor2_4 _22107_ (.A(_05938_),
    .B(_06032_),
    .Y(_06223_));
 sky130_fd_sc_hd__a2bb2o_1 _22108_ (.A1_N(_06222_),
    .A2_N(_06223_),
    .B1(_06222_),
    .B2(_06223_),
    .X(_06224_));
 sky130_vsdinv _22109_ (.A(\pcpi_mul.rs1[17] ),
    .Y(_06225_));
 sky130_fd_sc_hd__buf_1 _22110_ (.A(_06225_),
    .X(_06226_));
 sky130_fd_sc_hd__clkbuf_2 _22111_ (.A(_06226_),
    .X(_06227_));
 sky130_fd_sc_hd__or2_1 _22112_ (.A(_05834_),
    .B(_06227_),
    .X(_06228_));
 sky130_fd_sc_hd__clkbuf_2 _22113_ (.A(_05737_),
    .X(_06229_));
 sky130_fd_sc_hd__clkbuf_2 _22114_ (.A(_05739_),
    .X(_06230_));
 sky130_fd_sc_hd__clkbuf_2 _22115_ (.A(_05930_),
    .X(_06231_));
 sky130_fd_sc_hd__o22a_1 _22116_ (.A1(_06229_),
    .A2(_05735_),
    .B1(_06230_),
    .B2(_06231_),
    .X(_06232_));
 sky130_fd_sc_hd__clkbuf_2 _22117_ (.A(_13160_),
    .X(_06233_));
 sky130_fd_sc_hd__buf_1 _22118_ (.A(_13581_),
    .X(_06234_));
 sky130_fd_sc_hd__clkbuf_2 _22119_ (.A(_13166_),
    .X(_06235_));
 sky130_fd_sc_hd__buf_1 _22120_ (.A(_13578_),
    .X(_06236_));
 sky130_fd_sc_hd__and4_1 _22121_ (.A(_06233_),
    .B(_06234_),
    .C(_06235_),
    .D(_06236_),
    .X(_06237_));
 sky130_fd_sc_hd__or2_1 _22122_ (.A(_06232_),
    .B(_06237_),
    .X(_06238_));
 sky130_fd_sc_hd__a2bb2o_2 _22123_ (.A1_N(_06228_),
    .A2_N(_06238_),
    .B1(_06228_),
    .B2(_06238_),
    .X(_06239_));
 sky130_fd_sc_hd__o21ba_1 _22124_ (.A1(_06141_),
    .A2(_06147_),
    .B1_N(_06146_),
    .X(_06240_));
 sky130_fd_sc_hd__a2bb2o_1 _22125_ (.A1_N(_06239_),
    .A2_N(_06240_),
    .B1(_06239_),
    .B2(_06240_),
    .X(_06241_));
 sky130_fd_sc_hd__a2bb2o_1 _22126_ (.A1_N(_06224_),
    .A2_N(_06241_),
    .B1(_06224_),
    .B2(_06241_),
    .X(_06242_));
 sky130_fd_sc_hd__o22a_1 _22127_ (.A1(_06148_),
    .A2(_06149_),
    .B1(_06137_),
    .B2(_06150_),
    .X(_06243_));
 sky130_fd_sc_hd__a2bb2o_1 _22128_ (.A1_N(_06242_),
    .A2_N(_06243_),
    .B1(_06242_),
    .B2(_06243_),
    .X(_06244_));
 sky130_fd_sc_hd__a2bb2o_1 _22129_ (.A1_N(_06216_),
    .A2_N(_06244_),
    .B1(_06216_),
    .B2(_06244_),
    .X(_06245_));
 sky130_fd_sc_hd__o22a_1 _22130_ (.A1(_06158_),
    .A2(_06163_),
    .B1(_06157_),
    .B2(_06164_),
    .X(_06246_));
 sky130_fd_sc_hd__o22a_1 _22131_ (.A1(_06119_),
    .A2(_06120_),
    .B1(_06107_),
    .B2(_06121_),
    .X(_06247_));
 sky130_fd_sc_hd__o21ba_1 _22132_ (.A1(_06159_),
    .A2(_06162_),
    .B1_N(_06161_),
    .X(_06248_));
 sky130_fd_sc_hd__o21ba_1 _22133_ (.A1(_06100_),
    .A2(_06106_),
    .B1_N(_06105_),
    .X(_06249_));
 sky130_fd_sc_hd__or2_1 _22134_ (.A(_05423_),
    .B(_05817_),
    .X(_06250_));
 sky130_fd_sc_hd__clkbuf_2 _22135_ (.A(_05657_),
    .X(_06251_));
 sky130_fd_sc_hd__clkbuf_2 _22136_ (.A(_05456_),
    .X(_06252_));
 sky130_fd_sc_hd__o22a_1 _22137_ (.A1(_05865_),
    .A2(_06251_),
    .B1(_06252_),
    .B2(_05829_),
    .X(_06253_));
 sky130_fd_sc_hd__buf_1 _22138_ (.A(_13146_),
    .X(_06254_));
 sky130_fd_sc_hd__clkbuf_2 _22139_ (.A(_13152_),
    .X(_06255_));
 sky130_fd_sc_hd__and4_1 _22140_ (.A(_06254_),
    .B(_05654_),
    .C(_06255_),
    .D(_13587_),
    .X(_06256_));
 sky130_fd_sc_hd__or2_1 _22141_ (.A(_06253_),
    .B(_06256_),
    .X(_06257_));
 sky130_fd_sc_hd__a2bb2o_2 _22142_ (.A1_N(_06250_),
    .A2_N(_06257_),
    .B1(_06250_),
    .B2(_06257_),
    .X(_06258_));
 sky130_fd_sc_hd__a2bb2o_1 _22143_ (.A1_N(_06249_),
    .A2_N(_06258_),
    .B1(_06249_),
    .B2(_06258_),
    .X(_06259_));
 sky130_fd_sc_hd__a2bb2o_1 _22144_ (.A1_N(_06248_),
    .A2_N(_06259_),
    .B1(_06248_),
    .B2(_06259_),
    .X(_06260_));
 sky130_fd_sc_hd__a2bb2o_1 _22145_ (.A1_N(_06247_),
    .A2_N(_06260_),
    .B1(_06247_),
    .B2(_06260_),
    .X(_06261_));
 sky130_fd_sc_hd__a2bb2o_1 _22146_ (.A1_N(_06246_),
    .A2_N(_06261_),
    .B1(_06246_),
    .B2(_06261_),
    .X(_06262_));
 sky130_fd_sc_hd__o22a_1 _22147_ (.A1(_06156_),
    .A2(_06165_),
    .B1(_06155_),
    .B2(_06166_),
    .X(_06263_));
 sky130_fd_sc_hd__a2bb2o_1 _22148_ (.A1_N(_06262_),
    .A2_N(_06263_),
    .B1(_06262_),
    .B2(_06263_),
    .X(_06264_));
 sky130_fd_sc_hd__a2bb2o_1 _22149_ (.A1_N(_06245_),
    .A2_N(_06264_),
    .B1(_06245_),
    .B2(_06264_),
    .X(_06265_));
 sky130_fd_sc_hd__a2bb2o_1 _22150_ (.A1_N(_06125_),
    .A2_N(_06265_),
    .B1(_06125_),
    .B2(_06265_),
    .X(_06266_));
 sky130_fd_sc_hd__a2bb2o_1 _22151_ (.A1_N(_06215_),
    .A2_N(_06266_),
    .B1(_06215_),
    .B2(_06266_),
    .X(_06267_));
 sky130_fd_sc_hd__or2_1 _22152_ (.A(_06214_),
    .B(_06267_),
    .X(_06268_));
 sky130_fd_sc_hd__a21bo_1 _22153_ (.A1(_06214_),
    .A2(_06267_),
    .B1_N(_06268_),
    .X(_06269_));
 sky130_fd_sc_hd__a2bb2o_1 _22154_ (.A1_N(_06173_),
    .A2_N(_06269_),
    .B1(_06173_),
    .B2(_06269_),
    .X(_06270_));
 sky130_fd_sc_hd__a2bb2o_1 _22155_ (.A1_N(_06186_),
    .A2_N(_06270_),
    .B1(_06186_),
    .B2(_06270_),
    .X(_06271_));
 sky130_fd_sc_hd__o22a_1 _22156_ (.A1(_06072_),
    .A2(_06174_),
    .B1(_06085_),
    .B2(_06175_),
    .X(_06272_));
 sky130_fd_sc_hd__a2bb2o_1 _22157_ (.A1_N(_06271_),
    .A2_N(_06272_),
    .B1(_06271_),
    .B2(_06272_),
    .X(_06273_));
 sky130_fd_sc_hd__a2bb2o_1 _22158_ (.A1_N(_06084_),
    .A2_N(_06273_),
    .B1(_06084_),
    .B2(_06273_),
    .X(_06274_));
 sky130_fd_sc_hd__o22a_1 _22159_ (.A1(_06176_),
    .A2(_06177_),
    .B1(_05994_),
    .B2(_06178_),
    .X(_06275_));
 sky130_fd_sc_hd__or2_1 _22160_ (.A(_06274_),
    .B(_06275_),
    .X(_06276_));
 sky130_fd_sc_hd__a21bo_1 _22161_ (.A1(_06274_),
    .A2(_06275_),
    .B1_N(_06276_),
    .X(_06277_));
 sky130_fd_sc_hd__o21ai_1 _22162_ (.A1(_06082_),
    .A2(_06183_),
    .B1(_06181_),
    .Y(_06278_));
 sky130_fd_sc_hd__a2bb2o_1 _22163_ (.A1_N(_06277_),
    .A2_N(_06278_),
    .B1(_06277_),
    .B2(_06278_),
    .X(_02636_));
 sky130_fd_sc_hd__o22a_1 _22164_ (.A1(_06125_),
    .A2(_06265_),
    .B1(_06215_),
    .B2(_06266_),
    .X(_06279_));
 sky130_fd_sc_hd__o22a_1 _22165_ (.A1(_06242_),
    .A2(_06243_),
    .B1(_06216_),
    .B2(_06244_),
    .X(_06280_));
 sky130_fd_sc_hd__or2_2 _22166_ (.A(_06279_),
    .B(_06280_),
    .X(_06281_));
 sky130_fd_sc_hd__a21bo_1 _22167_ (.A1(_06279_),
    .A2(_06280_),
    .B1_N(_06281_),
    .X(_06282_));
 sky130_vsdinv _22168_ (.A(\pcpi_mul.rs2[18] ),
    .Y(_06283_));
 sky130_fd_sc_hd__clkbuf_2 _22169_ (.A(_06283_),
    .X(_06284_));
 sky130_fd_sc_hd__buf_2 _22170_ (.A(_06284_),
    .X(_06285_));
 sky130_fd_sc_hd__clkbuf_2 _22171_ (.A(_06285_),
    .X(_06286_));
 sky130_fd_sc_hd__buf_4 _22172_ (.A(_06286_),
    .X(_06287_));
 sky130_fd_sc_hd__or2_2 _22173_ (.A(_06287_),
    .B(_05154_),
    .X(_06288_));
 sky130_fd_sc_hd__or2_1 _22174_ (.A(_05996_),
    .B(_05338_),
    .X(_06289_));
 sky130_fd_sc_hd__o22a_1 _22175_ (.A1(_06189_),
    .A2(_05295_),
    .B1(_06086_),
    .B2(_05342_),
    .X(_06290_));
 sky130_fd_sc_hd__and4_1 _22176_ (.A(\pcpi_mul.rs2[17] ),
    .B(_13622_),
    .C(\pcpi_mul.rs2[16] ),
    .D(_05345_),
    .X(_06291_));
 sky130_fd_sc_hd__or2_1 _22177_ (.A(_06290_),
    .B(_06291_),
    .X(_06292_));
 sky130_fd_sc_hd__a2bb2o_1 _22178_ (.A1_N(_06289_),
    .A2_N(_06292_),
    .B1(_06289_),
    .B2(_06292_),
    .X(_06293_));
 sky130_fd_sc_hd__o21ba_1 _22179_ (.A1(_06188_),
    .A2(_06192_),
    .B1_N(_06191_),
    .X(_06294_));
 sky130_fd_sc_hd__or2_2 _22180_ (.A(_06293_),
    .B(_06294_),
    .X(_06295_));
 sky130_fd_sc_hd__a21bo_1 _22181_ (.A1(_06293_),
    .A2(_06294_),
    .B1_N(_06295_),
    .X(_06296_));
 sky130_fd_sc_hd__o2bb2ai_1 _22182_ (.A1_N(_06194_),
    .A2_N(_06296_),
    .B1(_06194_),
    .B2(_06296_),
    .Y(_06297_));
 sky130_fd_sc_hd__clkbuf_4 _22183_ (.A(_05946_),
    .X(_06298_));
 sky130_fd_sc_hd__or2_1 _22184_ (.A(_05711_),
    .B(_06298_),
    .X(_06299_));
 sky130_fd_sc_hd__buf_2 _22185_ (.A(_05713_),
    .X(_06300_));
 sky130_fd_sc_hd__clkbuf_2 _22186_ (.A(_05600_),
    .X(_06301_));
 sky130_fd_sc_hd__o22a_1 _22187_ (.A1(_06300_),
    .A2(_06301_),
    .B1(_05592_),
    .B2(_05963_),
    .X(_06302_));
 sky130_fd_sc_hd__buf_1 _22188_ (.A(_13597_),
    .X(_06303_));
 sky130_fd_sc_hd__buf_1 _22189_ (.A(_13593_),
    .X(_06304_));
 sky130_fd_sc_hd__and4_1 _22190_ (.A(_13136_),
    .B(_06303_),
    .C(_13142_),
    .D(_06304_),
    .X(_06305_));
 sky130_fd_sc_hd__or2_1 _22191_ (.A(_06302_),
    .B(_06305_),
    .X(_06306_));
 sky130_fd_sc_hd__a2bb2o_1 _22192_ (.A1_N(_06299_),
    .A2_N(_06306_),
    .B1(_06299_),
    .B2(_06306_),
    .X(_06307_));
 sky130_fd_sc_hd__clkbuf_2 _22193_ (.A(_05867_),
    .X(_06308_));
 sky130_fd_sc_hd__or2_1 _22194_ (.A(_05707_),
    .B(_06308_),
    .X(_06309_));
 sky130_fd_sc_hd__o22a_1 _22195_ (.A1(_06013_),
    .A2(_06005_),
    .B1(_06014_),
    .B2(_05899_),
    .X(_06310_));
 sky130_fd_sc_hd__buf_1 _22196_ (.A(_13607_),
    .X(_06311_));
 sky130_fd_sc_hd__and4_1 _22197_ (.A(_05916_),
    .B(_05904_),
    .C(_06017_),
    .D(_06311_),
    .X(_06312_));
 sky130_fd_sc_hd__or2_1 _22198_ (.A(_06310_),
    .B(_06312_),
    .X(_06313_));
 sky130_fd_sc_hd__a2bb2o_1 _22199_ (.A1_N(_06309_),
    .A2_N(_06313_),
    .B1(_06309_),
    .B2(_06313_),
    .X(_06314_));
 sky130_fd_sc_hd__o21ba_1 _22200_ (.A1(_06202_),
    .A2(_06206_),
    .B1_N(_06205_),
    .X(_06315_));
 sky130_fd_sc_hd__a2bb2o_1 _22201_ (.A1_N(_06314_),
    .A2_N(_06315_),
    .B1(_06314_),
    .B2(_06315_),
    .X(_06316_));
 sky130_fd_sc_hd__a2bb2o_1 _22202_ (.A1_N(_06307_),
    .A2_N(_06316_),
    .B1(_06307_),
    .B2(_06316_),
    .X(_06317_));
 sky130_fd_sc_hd__o2bb2a_1 _22203_ (.A1_N(_06297_),
    .A2_N(_06317_),
    .B1(_06297_),
    .B2(_06317_),
    .X(_06318_));
 sky130_fd_sc_hd__nand2_1 _22204_ (.A(_06211_),
    .B(_06318_),
    .Y(_06319_));
 sky130_fd_sc_hd__o21ai_1 _22205_ (.A1(_06211_),
    .A2(_06318_),
    .B1(_06319_),
    .Y(_06320_));
 sky130_fd_sc_hd__or2_1 _22206_ (.A(_06288_),
    .B(_06320_),
    .X(_06321_));
 sky130_vsdinv _22207_ (.A(_06321_),
    .Y(_06322_));
 sky130_fd_sc_hd__a21o_1 _22208_ (.A1(_06288_),
    .A2(_06320_),
    .B1(_06322_),
    .X(_06323_));
 sky130_fd_sc_hd__o22a_1 _22209_ (.A1(_06262_),
    .A2(_06263_),
    .B1(_06245_),
    .B2(_06264_),
    .X(_06324_));
 sky130_fd_sc_hd__a21oi_2 _22210_ (.A1(_06222_),
    .A2(_06223_),
    .B1(_06221_),
    .Y(_06325_));
 sky130_fd_sc_hd__buf_1 _22211_ (.A(_06138_),
    .X(_06326_));
 sky130_fd_sc_hd__buf_2 _22212_ (.A(_06326_),
    .X(_06327_));
 sky130_fd_sc_hd__buf_1 _22213_ (.A(_06225_),
    .X(_06328_));
 sky130_fd_sc_hd__buf_1 _22214_ (.A(_06328_),
    .X(_06329_));
 sky130_fd_sc_hd__buf_2 _22215_ (.A(_06329_),
    .X(_06330_));
 sky130_fd_sc_hd__o22a_1 _22216_ (.A1(_06217_),
    .A2(_06327_),
    .B1(_05929_),
    .B2(_06330_),
    .X(_06331_));
 sky130_fd_sc_hd__and4_1 _22217_ (.A(_13174_),
    .B(_13568_),
    .C(_13179_),
    .D(_13565_),
    .X(_06332_));
 sky130_fd_sc_hd__nor2_2 _22218_ (.A(_06331_),
    .B(_06332_),
    .Y(_06333_));
 sky130_fd_sc_hd__buf_2 _22219_ (.A(_06040_),
    .X(_06334_));
 sky130_fd_sc_hd__nor2_2 _22220_ (.A(_05938_),
    .B(_06334_),
    .Y(_06335_));
 sky130_fd_sc_hd__a2bb2o_1 _22221_ (.A1_N(_06333_),
    .A2_N(_06335_),
    .B1(_06333_),
    .B2(_06335_),
    .X(_06336_));
 sky130_vsdinv _22222_ (.A(\pcpi_mul.rs1[18] ),
    .Y(_06337_));
 sky130_fd_sc_hd__buf_1 _22223_ (.A(_06337_),
    .X(_06338_));
 sky130_fd_sc_hd__clkbuf_2 _22224_ (.A(_06338_),
    .X(_06339_));
 sky130_fd_sc_hd__or2_1 _22225_ (.A(_05834_),
    .B(_06339_),
    .X(_06340_));
 sky130_fd_sc_hd__o22a_1 _22226_ (.A1(_06229_),
    .A2(_05836_),
    .B1(_06230_),
    .B2(_06129_),
    .X(_06341_));
 sky130_fd_sc_hd__buf_1 _22227_ (.A(\pcpi_mul.rs1[14] ),
    .X(_06342_));
 sky130_fd_sc_hd__and4_1 _22228_ (.A(_05845_),
    .B(_06236_),
    .C(_05847_),
    .D(_06342_),
    .X(_06343_));
 sky130_fd_sc_hd__or2_1 _22229_ (.A(_06341_),
    .B(_06343_),
    .X(_06344_));
 sky130_fd_sc_hd__a2bb2o_1 _22230_ (.A1_N(_06340_),
    .A2_N(_06344_),
    .B1(_06340_),
    .B2(_06344_),
    .X(_06345_));
 sky130_fd_sc_hd__o21ba_1 _22231_ (.A1(_06228_),
    .A2(_06238_),
    .B1_N(_06237_),
    .X(_06346_));
 sky130_fd_sc_hd__a2bb2o_1 _22232_ (.A1_N(_06345_),
    .A2_N(_06346_),
    .B1(_06345_),
    .B2(_06346_),
    .X(_06347_));
 sky130_fd_sc_hd__a2bb2o_2 _22233_ (.A1_N(_06336_),
    .A2_N(_06347_),
    .B1(_06336_),
    .B2(_06347_),
    .X(_06348_));
 sky130_fd_sc_hd__o22a_1 _22234_ (.A1(_06239_),
    .A2(_06240_),
    .B1(_06224_),
    .B2(_06241_),
    .X(_06349_));
 sky130_fd_sc_hd__a2bb2o_1 _22235_ (.A1_N(_06348_),
    .A2_N(_06349_),
    .B1(_06348_),
    .B2(_06349_),
    .X(_06350_));
 sky130_fd_sc_hd__a2bb2o_1 _22236_ (.A1_N(_06325_),
    .A2_N(_06350_),
    .B1(_06325_),
    .B2(_06350_),
    .X(_06351_));
 sky130_fd_sc_hd__o22a_1 _22237_ (.A1(_06249_),
    .A2(_06258_),
    .B1(_06248_),
    .B2(_06259_),
    .X(_06352_));
 sky130_fd_sc_hd__o22a_1 _22238_ (.A1(_06207_),
    .A2(_06208_),
    .B1(_06200_),
    .B2(_06209_),
    .X(_06353_));
 sky130_fd_sc_hd__o21ba_1 _22239_ (.A1(_06250_),
    .A2(_06257_),
    .B1_N(_06256_),
    .X(_06354_));
 sky130_fd_sc_hd__o21ba_1 _22240_ (.A1(_06196_),
    .A2(_06199_),
    .B1_N(_06198_),
    .X(_06355_));
 sky130_fd_sc_hd__clkbuf_2 _22241_ (.A(_05926_),
    .X(_06356_));
 sky130_fd_sc_hd__or2_1 _22242_ (.A(_05423_),
    .B(_06356_),
    .X(_06357_));
 sky130_fd_sc_hd__o22a_1 _22243_ (.A1(_05965_),
    .A2(_05829_),
    .B1(_06252_),
    .B2(_05724_),
    .X(_06358_));
 sky130_fd_sc_hd__and4_1 _22244_ (.A(_06254_),
    .B(_13587_),
    .C(_06255_),
    .D(_06143_),
    .X(_06359_));
 sky130_fd_sc_hd__or2_1 _22245_ (.A(_06358_),
    .B(_06359_),
    .X(_06360_));
 sky130_fd_sc_hd__a2bb2o_2 _22246_ (.A1_N(_06357_),
    .A2_N(_06360_),
    .B1(_06357_),
    .B2(_06360_),
    .X(_06361_));
 sky130_fd_sc_hd__a2bb2o_1 _22247_ (.A1_N(_06355_),
    .A2_N(_06361_),
    .B1(_06355_),
    .B2(_06361_),
    .X(_06362_));
 sky130_fd_sc_hd__a2bb2o_1 _22248_ (.A1_N(_06354_),
    .A2_N(_06362_),
    .B1(_06354_),
    .B2(_06362_),
    .X(_06363_));
 sky130_fd_sc_hd__a2bb2o_1 _22249_ (.A1_N(_06353_),
    .A2_N(_06363_),
    .B1(_06353_),
    .B2(_06363_),
    .X(_06364_));
 sky130_fd_sc_hd__a2bb2o_1 _22250_ (.A1_N(_06352_),
    .A2_N(_06364_),
    .B1(_06352_),
    .B2(_06364_),
    .X(_06365_));
 sky130_fd_sc_hd__o22a_1 _22251_ (.A1(_06247_),
    .A2(_06260_),
    .B1(_06246_),
    .B2(_06261_),
    .X(_06366_));
 sky130_fd_sc_hd__a2bb2o_1 _22252_ (.A1_N(_06365_),
    .A2_N(_06366_),
    .B1(_06365_),
    .B2(_06366_),
    .X(_06367_));
 sky130_fd_sc_hd__a2bb2o_1 _22253_ (.A1_N(_06351_),
    .A2_N(_06367_),
    .B1(_06351_),
    .B2(_06367_),
    .X(_06368_));
 sky130_fd_sc_hd__a2bb2o_1 _22254_ (.A1_N(_06213_),
    .A2_N(_06368_),
    .B1(_06213_),
    .B2(_06368_),
    .X(_06369_));
 sky130_fd_sc_hd__a2bb2o_1 _22255_ (.A1_N(_06324_),
    .A2_N(_06369_),
    .B1(_06324_),
    .B2(_06369_),
    .X(_06370_));
 sky130_fd_sc_hd__or2_1 _22256_ (.A(_06323_),
    .B(_06370_),
    .X(_06371_));
 sky130_fd_sc_hd__a21bo_1 _22257_ (.A1(_06323_),
    .A2(_06370_),
    .B1_N(_06371_),
    .X(_06372_));
 sky130_fd_sc_hd__a2bb2o_1 _22258_ (.A1_N(_06268_),
    .A2_N(_06372_),
    .B1(_06268_),
    .B2(_06372_),
    .X(_06373_));
 sky130_fd_sc_hd__a2bb2o_1 _22259_ (.A1_N(_06282_),
    .A2_N(_06373_),
    .B1(_06282_),
    .B2(_06373_),
    .X(_06374_));
 sky130_fd_sc_hd__o22a_1 _22260_ (.A1(_06173_),
    .A2(_06269_),
    .B1(_06186_),
    .B2(_06270_),
    .X(_06375_));
 sky130_fd_sc_hd__a2bb2o_1 _22261_ (.A1_N(_06374_),
    .A2_N(_06375_),
    .B1(_06374_),
    .B2(_06375_),
    .X(_06376_));
 sky130_fd_sc_hd__a2bb2o_1 _22262_ (.A1_N(_06185_),
    .A2_N(_06376_),
    .B1(_06185_),
    .B2(_06376_),
    .X(_06377_));
 sky130_fd_sc_hd__o22a_1 _22263_ (.A1(_06271_),
    .A2(_06272_),
    .B1(_06084_),
    .B2(_06273_),
    .X(_06378_));
 sky130_fd_sc_hd__or2_1 _22264_ (.A(_06377_),
    .B(_06378_),
    .X(_06379_));
 sky130_fd_sc_hd__a21bo_2 _22265_ (.A1(_06377_),
    .A2(_06378_),
    .B1_N(_06379_),
    .X(_06380_));
 sky130_fd_sc_hd__a22o_1 _22266_ (.A1(_06274_),
    .A2(_06275_),
    .B1(_06181_),
    .B2(_06276_),
    .X(_06381_));
 sky130_fd_sc_hd__o31a_2 _22267_ (.A1(_06183_),
    .A2(_06277_),
    .A3(_06082_),
    .B1(_06381_),
    .X(_06382_));
 sky130_fd_sc_hd__a2bb2oi_4 _22268_ (.A1_N(_06380_),
    .A2_N(_06382_),
    .B1(_06380_),
    .B2(_06382_),
    .Y(_02637_));
 sky130_fd_sc_hd__o22a_1 _22269_ (.A1(_06374_),
    .A2(_06375_),
    .B1(_06185_),
    .B2(_06376_),
    .X(_06383_));
 sky130_fd_sc_hd__o22a_1 _22270_ (.A1(_06213_),
    .A2(_06368_),
    .B1(_06324_),
    .B2(_06369_),
    .X(_06384_));
 sky130_fd_sc_hd__o22a_1 _22271_ (.A1(_06348_),
    .A2(_06349_),
    .B1(_06325_),
    .B2(_06350_),
    .X(_06385_));
 sky130_fd_sc_hd__or2_1 _22272_ (.A(_06384_),
    .B(_06385_),
    .X(_06386_));
 sky130_fd_sc_hd__a21bo_1 _22273_ (.A1(_06384_),
    .A2(_06385_),
    .B1_N(_06386_),
    .X(_06387_));
 sky130_vsdinv _22274_ (.A(\pcpi_mul.rs2[19] ),
    .Y(_06388_));
 sky130_fd_sc_hd__clkbuf_2 _22275_ (.A(_06388_),
    .X(_06389_));
 sky130_fd_sc_hd__clkbuf_2 _22276_ (.A(_06389_),
    .X(_06390_));
 sky130_fd_sc_hd__clkbuf_2 _22277_ (.A(_06390_),
    .X(_06391_));
 sky130_fd_sc_hd__clkbuf_4 _22278_ (.A(_06391_),
    .X(_06392_));
 sky130_fd_sc_hd__o22a_2 _22279_ (.A1(_06392_),
    .A2(_05590_),
    .B1(_06287_),
    .B2(_05300_),
    .X(_06393_));
 sky130_fd_sc_hd__buf_1 _22280_ (.A(_06388_),
    .X(_06394_));
 sky130_fd_sc_hd__buf_1 _22281_ (.A(_06394_),
    .X(_06395_));
 sky130_fd_sc_hd__clkbuf_2 _22282_ (.A(_06283_),
    .X(_06396_));
 sky130_fd_sc_hd__or4_4 _22283_ (.A(_06395_),
    .B(_05149_),
    .C(_06396_),
    .D(_05319_),
    .X(_06397_));
 sky130_fd_sc_hd__or2b_1 _22284_ (.A(_06393_),
    .B_N(_06397_),
    .X(_06398_));
 sky130_fd_sc_hd__buf_2 _22285_ (.A(_05722_),
    .X(_06399_));
 sky130_fd_sc_hd__or2_1 _22286_ (.A(_05711_),
    .B(_06399_),
    .X(_06400_));
 sky130_fd_sc_hd__o22a_1 _22287_ (.A1(_06300_),
    .A2(_05841_),
    .B1(_05592_),
    .B2(_05843_),
    .X(_06401_));
 sky130_fd_sc_hd__and4_1 _22288_ (.A(_13136_),
    .B(_06304_),
    .C(_13142_),
    .D(_13591_),
    .X(_06402_));
 sky130_fd_sc_hd__or2_1 _22289_ (.A(_06401_),
    .B(_06402_),
    .X(_06403_));
 sky130_fd_sc_hd__a2bb2o_1 _22290_ (.A1_N(_06400_),
    .A2_N(_06403_),
    .B1(_06400_),
    .B2(_06403_),
    .X(_06404_));
 sky130_fd_sc_hd__or2_1 _22291_ (.A(_05790_),
    .B(_06301_),
    .X(_06405_));
 sky130_fd_sc_hd__o22a_1 _22292_ (.A1(_05912_),
    .A2(_05680_),
    .B1(_06014_),
    .B2(_05867_),
    .X(_06406_));
 sky130_fd_sc_hd__and4_1 _22293_ (.A(_06114_),
    .B(_06007_),
    .C(_06017_),
    .D(_05969_),
    .X(_06407_));
 sky130_fd_sc_hd__or2_1 _22294_ (.A(_06406_),
    .B(_06407_),
    .X(_06408_));
 sky130_fd_sc_hd__a2bb2o_1 _22295_ (.A1_N(_06405_),
    .A2_N(_06408_),
    .B1(_06405_),
    .B2(_06408_),
    .X(_06409_));
 sky130_fd_sc_hd__o21ba_1 _22296_ (.A1(_06309_),
    .A2(_06313_),
    .B1_N(_06312_),
    .X(_06410_));
 sky130_fd_sc_hd__a2bb2o_1 _22297_ (.A1_N(_06409_),
    .A2_N(_06410_),
    .B1(_06409_),
    .B2(_06410_),
    .X(_06411_));
 sky130_fd_sc_hd__a2bb2o_1 _22298_ (.A1_N(_06404_),
    .A2_N(_06411_),
    .B1(_06404_),
    .B2(_06411_),
    .X(_06412_));
 sky130_fd_sc_hd__or2_1 _22299_ (.A(_05997_),
    .B(_05366_),
    .X(_06413_));
 sky130_fd_sc_hd__o22a_1 _22300_ (.A1(_06189_),
    .A2(_05342_),
    .B1(_06087_),
    .B2(_05683_),
    .X(_06414_));
 sky130_fd_sc_hd__and4_1 _22301_ (.A(_13116_),
    .B(_13619_),
    .C(\pcpi_mul.rs2[16] ),
    .D(_05376_),
    .X(_06415_));
 sky130_fd_sc_hd__or2_1 _22302_ (.A(_06414_),
    .B(_06415_),
    .X(_06416_));
 sky130_fd_sc_hd__a2bb2o_1 _22303_ (.A1_N(_06413_),
    .A2_N(_06416_),
    .B1(_06413_),
    .B2(_06416_),
    .X(_06417_));
 sky130_fd_sc_hd__o21ba_1 _22304_ (.A1(_06289_),
    .A2(_06292_),
    .B1_N(_06291_),
    .X(_06418_));
 sky130_fd_sc_hd__or2_1 _22305_ (.A(_06417_),
    .B(_06418_),
    .X(_06419_));
 sky130_fd_sc_hd__a21bo_1 _22306_ (.A1(_06417_),
    .A2(_06418_),
    .B1_N(_06419_),
    .X(_06420_));
 sky130_fd_sc_hd__a2bb2o_1 _22307_ (.A1_N(_06295_),
    .A2_N(_06420_),
    .B1(_06295_),
    .B2(_06420_),
    .X(_06421_));
 sky130_fd_sc_hd__a2bb2o_1 _22308_ (.A1_N(_06412_),
    .A2_N(_06421_),
    .B1(_06412_),
    .B2(_06421_),
    .X(_06422_));
 sky130_fd_sc_hd__o22a_1 _22309_ (.A1(_06194_),
    .A2(_06296_),
    .B1(_06297_),
    .B2(_06317_),
    .X(_06423_));
 sky130_fd_sc_hd__or2_1 _22310_ (.A(_06422_),
    .B(_06423_),
    .X(_06424_));
 sky130_fd_sc_hd__a21bo_1 _22311_ (.A1(_06422_),
    .A2(_06423_),
    .B1_N(_06424_),
    .X(_06425_));
 sky130_fd_sc_hd__or2_1 _22312_ (.A(_06398_),
    .B(_06425_),
    .X(_06426_));
 sky130_vsdinv _22313_ (.A(_06426_),
    .Y(_06427_));
 sky130_fd_sc_hd__a21oi_2 _22314_ (.A1(_06398_),
    .A2(_06425_),
    .B1(_06427_),
    .Y(_06428_));
 sky130_vsdinv _22315_ (.A(_06428_),
    .Y(_06429_));
 sky130_fd_sc_hd__a22o_1 _22316_ (.A1(_06321_),
    .A2(_06429_),
    .B1(_06322_),
    .B2(_06428_),
    .X(_06430_));
 sky130_fd_sc_hd__o22a_1 _22317_ (.A1(_06365_),
    .A2(_06366_),
    .B1(_06351_),
    .B2(_06367_),
    .X(_06431_));
 sky130_fd_sc_hd__a21oi_2 _22318_ (.A1(_06333_),
    .A2(_06335_),
    .B1(_06332_),
    .Y(_06432_));
 sky130_fd_sc_hd__clkbuf_2 _22319_ (.A(_06217_),
    .X(_06433_));
 sky130_fd_sc_hd__clkbuf_2 _22320_ (.A(_06328_),
    .X(_06434_));
 sky130_fd_sc_hd__buf_2 _22321_ (.A(_06434_),
    .X(_06435_));
 sky130_fd_sc_hd__clkbuf_2 _22322_ (.A(_05929_),
    .X(_06436_));
 sky130_fd_sc_hd__clkbuf_2 _22323_ (.A(_06337_),
    .X(_06437_));
 sky130_fd_sc_hd__buf_2 _22324_ (.A(_06437_),
    .X(_06438_));
 sky130_fd_sc_hd__clkbuf_4 _22325_ (.A(_06438_),
    .X(_06439_));
 sky130_fd_sc_hd__o22a_1 _22326_ (.A1(_06433_),
    .A2(_06435_),
    .B1(_06436_),
    .B2(_06439_),
    .X(_06440_));
 sky130_fd_sc_hd__buf_1 _22327_ (.A(_05934_),
    .X(_06441_));
 sky130_fd_sc_hd__buf_1 _22328_ (.A(_05935_),
    .X(_06442_));
 sky130_fd_sc_hd__and4_1 _22329_ (.A(_06441_),
    .B(_13565_),
    .C(_06442_),
    .D(_13561_),
    .X(_06443_));
 sky130_fd_sc_hd__nor2_2 _22330_ (.A(_06440_),
    .B(_06443_),
    .Y(_06444_));
 sky130_fd_sc_hd__clkbuf_2 _22331_ (.A(_05828_),
    .X(_06445_));
 sky130_fd_sc_hd__nor2_2 _22332_ (.A(_06445_),
    .B(_06219_),
    .Y(_06446_));
 sky130_fd_sc_hd__a2bb2o_1 _22333_ (.A1_N(_06444_),
    .A2_N(_06446_),
    .B1(_06444_),
    .B2(_06446_),
    .X(_06447_));
 sky130_fd_sc_hd__buf_1 _22334_ (.A(_05834_),
    .X(_06448_));
 sky130_vsdinv _22335_ (.A(\pcpi_mul.rs1[19] ),
    .Y(_06449_));
 sky130_fd_sc_hd__buf_1 _22336_ (.A(_06449_),
    .X(_06450_));
 sky130_fd_sc_hd__buf_1 _22337_ (.A(_06450_),
    .X(_06451_));
 sky130_fd_sc_hd__buf_4 _22338_ (.A(_06451_),
    .X(_06452_));
 sky130_fd_sc_hd__or2_1 _22339_ (.A(_06448_),
    .B(_06452_),
    .X(_06453_));
 sky130_fd_sc_hd__clkbuf_2 _22340_ (.A(_06229_),
    .X(_06454_));
 sky130_fd_sc_hd__clkbuf_2 _22341_ (.A(_06230_),
    .X(_06455_));
 sky130_fd_sc_hd__buf_1 _22342_ (.A(_06038_),
    .X(_06456_));
 sky130_fd_sc_hd__clkbuf_2 _22343_ (.A(_06456_),
    .X(_06457_));
 sky130_fd_sc_hd__o22a_1 _22344_ (.A1(_06454_),
    .A2(_05944_),
    .B1(_06455_),
    .B2(_06457_),
    .X(_06458_));
 sky130_fd_sc_hd__buf_1 _22345_ (.A(_05845_),
    .X(_06459_));
 sky130_fd_sc_hd__clkbuf_2 _22346_ (.A(_06342_),
    .X(_06460_));
 sky130_fd_sc_hd__buf_1 _22347_ (.A(_05847_),
    .X(_06461_));
 sky130_fd_sc_hd__buf_1 _22348_ (.A(\pcpi_mul.rs1[15] ),
    .X(_06462_));
 sky130_fd_sc_hd__buf_1 _22349_ (.A(_06462_),
    .X(_06463_));
 sky130_fd_sc_hd__and4_1 _22350_ (.A(_06459_),
    .B(_06460_),
    .C(_06461_),
    .D(_06463_),
    .X(_06464_));
 sky130_fd_sc_hd__or2_1 _22351_ (.A(_06458_),
    .B(_06464_),
    .X(_06465_));
 sky130_fd_sc_hd__a2bb2o_1 _22352_ (.A1_N(_06453_),
    .A2_N(_06465_),
    .B1(_06453_),
    .B2(_06465_),
    .X(_06466_));
 sky130_fd_sc_hd__o21ba_1 _22353_ (.A1(_06340_),
    .A2(_06344_),
    .B1_N(_06343_),
    .X(_06467_));
 sky130_fd_sc_hd__a2bb2o_1 _22354_ (.A1_N(_06466_),
    .A2_N(_06467_),
    .B1(_06466_),
    .B2(_06467_),
    .X(_06468_));
 sky130_fd_sc_hd__a2bb2o_1 _22355_ (.A1_N(_06447_),
    .A2_N(_06468_),
    .B1(_06447_),
    .B2(_06468_),
    .X(_06469_));
 sky130_fd_sc_hd__o22a_1 _22356_ (.A1(_06345_),
    .A2(_06346_),
    .B1(_06336_),
    .B2(_06347_),
    .X(_06470_));
 sky130_fd_sc_hd__a2bb2o_1 _22357_ (.A1_N(_06469_),
    .A2_N(_06470_),
    .B1(_06469_),
    .B2(_06470_),
    .X(_06471_));
 sky130_fd_sc_hd__a2bb2o_2 _22358_ (.A1_N(_06432_),
    .A2_N(_06471_),
    .B1(_06432_),
    .B2(_06471_),
    .X(_06472_));
 sky130_fd_sc_hd__o22a_1 _22359_ (.A1(_06355_),
    .A2(_06361_),
    .B1(_06354_),
    .B2(_06362_),
    .X(_06473_));
 sky130_fd_sc_hd__o22a_1 _22360_ (.A1(_06314_),
    .A2(_06315_),
    .B1(_06307_),
    .B2(_06316_),
    .X(_06474_));
 sky130_fd_sc_hd__o21ba_1 _22361_ (.A1(_06357_),
    .A2(_06360_),
    .B1_N(_06359_),
    .X(_06475_));
 sky130_fd_sc_hd__o21ba_1 _22362_ (.A1(_06299_),
    .A2(_06306_),
    .B1_N(_06305_),
    .X(_06476_));
 sky130_fd_sc_hd__clkbuf_2 _22363_ (.A(_05962_),
    .X(_06477_));
 sky130_fd_sc_hd__buf_1 _22364_ (.A(_05835_),
    .X(_06478_));
 sky130_fd_sc_hd__clkbuf_2 _22365_ (.A(_06478_),
    .X(_06479_));
 sky130_fd_sc_hd__or2_1 _22366_ (.A(_06477_),
    .B(_06479_),
    .X(_06480_));
 sky130_fd_sc_hd__clkbuf_2 _22367_ (.A(_05965_),
    .X(_06481_));
 sky130_fd_sc_hd__clkbuf_2 _22368_ (.A(_05667_),
    .X(_06482_));
 sky130_fd_sc_hd__clkbuf_2 _22369_ (.A(_05966_),
    .X(_06483_));
 sky130_fd_sc_hd__clkbuf_2 _22370_ (.A(_05926_),
    .X(_06484_));
 sky130_fd_sc_hd__o22a_1 _22371_ (.A1(_06481_),
    .A2(_06482_),
    .B1(_06483_),
    .B2(_06484_),
    .X(_06485_));
 sky130_fd_sc_hd__buf_1 _22372_ (.A(_06143_),
    .X(_06486_));
 sky130_fd_sc_hd__and4_1 _22373_ (.A(_13148_),
    .B(_06486_),
    .C(_13154_),
    .D(_13582_),
    .X(_06487_));
 sky130_fd_sc_hd__or2_1 _22374_ (.A(_06485_),
    .B(_06487_),
    .X(_06488_));
 sky130_fd_sc_hd__a2bb2o_2 _22375_ (.A1_N(_06480_),
    .A2_N(_06488_),
    .B1(_06480_),
    .B2(_06488_),
    .X(_06489_));
 sky130_fd_sc_hd__a2bb2o_1 _22376_ (.A1_N(_06476_),
    .A2_N(_06489_),
    .B1(_06476_),
    .B2(_06489_),
    .X(_06490_));
 sky130_fd_sc_hd__a2bb2o_1 _22377_ (.A1_N(_06475_),
    .A2_N(_06490_),
    .B1(_06475_),
    .B2(_06490_),
    .X(_06491_));
 sky130_fd_sc_hd__a2bb2o_1 _22378_ (.A1_N(_06474_),
    .A2_N(_06491_),
    .B1(_06474_),
    .B2(_06491_),
    .X(_06492_));
 sky130_fd_sc_hd__a2bb2o_1 _22379_ (.A1_N(_06473_),
    .A2_N(_06492_),
    .B1(_06473_),
    .B2(_06492_),
    .X(_06493_));
 sky130_fd_sc_hd__o22a_1 _22380_ (.A1(_06353_),
    .A2(_06363_),
    .B1(_06352_),
    .B2(_06364_),
    .X(_06494_));
 sky130_fd_sc_hd__a2bb2o_1 _22381_ (.A1_N(_06493_),
    .A2_N(_06494_),
    .B1(_06493_),
    .B2(_06494_),
    .X(_06495_));
 sky130_fd_sc_hd__a2bb2o_1 _22382_ (.A1_N(_06472_),
    .A2_N(_06495_),
    .B1(_06472_),
    .B2(_06495_),
    .X(_06496_));
 sky130_fd_sc_hd__a2bb2o_1 _22383_ (.A1_N(_06319_),
    .A2_N(_06496_),
    .B1(_06319_),
    .B2(_06496_),
    .X(_06497_));
 sky130_fd_sc_hd__a2bb2o_1 _22384_ (.A1_N(_06431_),
    .A2_N(_06497_),
    .B1(_06431_),
    .B2(_06497_),
    .X(_06498_));
 sky130_fd_sc_hd__a2bb2o_1 _22385_ (.A1_N(_06430_),
    .A2_N(_06498_),
    .B1(_06430_),
    .B2(_06498_),
    .X(_06499_));
 sky130_fd_sc_hd__a2bb2o_1 _22386_ (.A1_N(_06371_),
    .A2_N(_06499_),
    .B1(_06371_),
    .B2(_06499_),
    .X(_06500_));
 sky130_fd_sc_hd__a2bb2o_1 _22387_ (.A1_N(_06387_),
    .A2_N(_06500_),
    .B1(_06387_),
    .B2(_06500_),
    .X(_06501_));
 sky130_fd_sc_hd__o22a_1 _22388_ (.A1(_06268_),
    .A2(_06372_),
    .B1(_06282_),
    .B2(_06373_),
    .X(_06502_));
 sky130_fd_sc_hd__a2bb2o_1 _22389_ (.A1_N(_06501_),
    .A2_N(_06502_),
    .B1(_06501_),
    .B2(_06502_),
    .X(_06503_));
 sky130_fd_sc_hd__a2bb2o_1 _22390_ (.A1_N(_06281_),
    .A2_N(_06503_),
    .B1(_06281_),
    .B2(_06503_),
    .X(_06504_));
 sky130_fd_sc_hd__and2_1 _22391_ (.A(_06383_),
    .B(_06504_),
    .X(_06505_));
 sky130_fd_sc_hd__or2_1 _22392_ (.A(_06383_),
    .B(_06504_),
    .X(_06506_));
 sky130_fd_sc_hd__or2b_2 _22393_ (.A(_06505_),
    .B_N(_06506_),
    .X(_06507_));
 sky130_fd_sc_hd__o21ai_2 _22394_ (.A1(_06380_),
    .A2(_06382_),
    .B1(_06379_),
    .Y(_06508_));
 sky130_fd_sc_hd__a2bb2o_4 _22395_ (.A1_N(_06507_),
    .A2_N(_06508_),
    .B1(_06507_),
    .B2(_06508_),
    .X(_02638_));
 sky130_fd_sc_hd__o22a_1 _22396_ (.A1(_06319_),
    .A2(_06496_),
    .B1(_06431_),
    .B2(_06497_),
    .X(_06509_));
 sky130_fd_sc_hd__o22a_2 _22397_ (.A1(_06469_),
    .A2(_06470_),
    .B1(_06432_),
    .B2(_06471_),
    .X(_06510_));
 sky130_fd_sc_hd__or2_1 _22398_ (.A(_06509_),
    .B(_06510_),
    .X(_06511_));
 sky130_fd_sc_hd__a21bo_1 _22399_ (.A1(_06509_),
    .A2(_06510_),
    .B1_N(_06511_),
    .X(_06512_));
 sky130_fd_sc_hd__or2_1 _22400_ (.A(_06283_),
    .B(_05908_),
    .X(_06513_));
 sky130_vsdinv _22401_ (.A(\pcpi_mul.rs2[20] ),
    .Y(_06514_));
 sky130_fd_sc_hd__o22a_1 _22402_ (.A1(_06388_),
    .A2(_05296_),
    .B1(_06514_),
    .B2(_05363_),
    .X(_06515_));
 sky130_fd_sc_hd__and4_1 _22403_ (.A(_13110_),
    .B(_13623_),
    .C(\pcpi_mul.rs2[20] ),
    .D(_05917_),
    .X(_06516_));
 sky130_fd_sc_hd__or2_1 _22404_ (.A(_06515_),
    .B(_06516_),
    .X(_06517_));
 sky130_fd_sc_hd__a2bb2o_1 _22405_ (.A1_N(_06513_),
    .A2_N(_06517_),
    .B1(_06513_),
    .B2(_06517_),
    .X(_06518_));
 sky130_fd_sc_hd__buf_2 _22406_ (.A(_05797_),
    .X(_06519_));
 sky130_fd_sc_hd__clkbuf_2 _22407_ (.A(_06482_),
    .X(_06520_));
 sky130_fd_sc_hd__or2_1 _22408_ (.A(_06519_),
    .B(_06520_),
    .X(_06521_));
 sky130_fd_sc_hd__clkbuf_2 _22409_ (.A(_05801_),
    .X(_06522_));
 sky130_fd_sc_hd__clkbuf_2 _22410_ (.A(_05802_),
    .X(_06523_));
 sky130_fd_sc_hd__o22a_1 _22411_ (.A1(_06522_),
    .A2(_05946_),
    .B1(_06523_),
    .B2(_05947_),
    .X(_06524_));
 sky130_fd_sc_hd__clkbuf_2 _22412_ (.A(_05805_),
    .X(_06525_));
 sky130_fd_sc_hd__buf_1 _22413_ (.A(_05654_),
    .X(_06526_));
 sky130_fd_sc_hd__clkbuf_2 _22414_ (.A(_05807_),
    .X(_06527_));
 sky130_fd_sc_hd__buf_1 _22415_ (.A(_05655_),
    .X(_06528_));
 sky130_fd_sc_hd__and4_1 _22416_ (.A(_06525_),
    .B(_06526_),
    .C(_06527_),
    .D(_06528_),
    .X(_06529_));
 sky130_fd_sc_hd__or2_1 _22417_ (.A(_06524_),
    .B(_06529_),
    .X(_06530_));
 sky130_fd_sc_hd__a2bb2o_2 _22418_ (.A1_N(_06521_),
    .A2_N(_06530_),
    .B1(_06521_),
    .B2(_06530_),
    .X(_06531_));
 sky130_fd_sc_hd__or2_1 _22419_ (.A(_05794_),
    .B(_05663_),
    .X(_06532_));
 sky130_fd_sc_hd__clkbuf_4 _22420_ (.A(_05787_),
    .X(_06533_));
 sky130_fd_sc_hd__o22a_1 _22421_ (.A1(_06110_),
    .A2(_06101_),
    .B1(_06533_),
    .B2(_05861_),
    .X(_06534_));
 sky130_fd_sc_hd__buf_2 _22422_ (.A(_13128_),
    .X(_06535_));
 sky130_fd_sc_hd__buf_2 _22423_ (.A(_13131_),
    .X(_06536_));
 sky130_fd_sc_hd__and4_1 _22424_ (.A(_06535_),
    .B(_13603_),
    .C(_06536_),
    .D(_13598_),
    .X(_06537_));
 sky130_fd_sc_hd__or2_1 _22425_ (.A(_06534_),
    .B(_06537_),
    .X(_06538_));
 sky130_fd_sc_hd__a2bb2o_1 _22426_ (.A1_N(_06532_),
    .A2_N(_06538_),
    .B1(_06532_),
    .B2(_06538_),
    .X(_06539_));
 sky130_fd_sc_hd__o21ba_1 _22427_ (.A1(_06405_),
    .A2(_06408_),
    .B1_N(_06407_),
    .X(_06540_));
 sky130_fd_sc_hd__a2bb2o_1 _22428_ (.A1_N(_06539_),
    .A2_N(_06540_),
    .B1(_06539_),
    .B2(_06540_),
    .X(_06541_));
 sky130_fd_sc_hd__a2bb2o_1 _22429_ (.A1_N(_06531_),
    .A2_N(_06541_),
    .B1(_06531_),
    .B2(_06541_),
    .X(_06542_));
 sky130_fd_sc_hd__o21ba_1 _22430_ (.A1(_06413_),
    .A2(_06416_),
    .B1_N(_06415_),
    .X(_06543_));
 sky130_fd_sc_hd__buf_2 _22431_ (.A(_05509_),
    .X(_06544_));
 sky130_fd_sc_hd__or2_1 _22432_ (.A(_05997_),
    .B(_06544_),
    .X(_06545_));
 sky130_fd_sc_hd__buf_1 _22433_ (.A(_06189_),
    .X(_06546_));
 sky130_fd_sc_hd__o22a_1 _22434_ (.A1(_06546_),
    .A2(_05338_),
    .B1(_06087_),
    .B2(_05366_),
    .X(_06547_));
 sky130_fd_sc_hd__and4_1 _22435_ (.A(_13116_),
    .B(_06204_),
    .C(_13120_),
    .D(_05758_),
    .X(_06548_));
 sky130_fd_sc_hd__or2_1 _22436_ (.A(_06547_),
    .B(_06548_),
    .X(_06549_));
 sky130_fd_sc_hd__a2bb2o_1 _22437_ (.A1_N(_06545_),
    .A2_N(_06549_),
    .B1(_06545_),
    .B2(_06549_),
    .X(_06550_));
 sky130_fd_sc_hd__a2bb2o_1 _22438_ (.A1_N(_06397_),
    .A2_N(_06550_),
    .B1(_06397_),
    .B2(_06550_),
    .X(_06551_));
 sky130_fd_sc_hd__a2bb2o_1 _22439_ (.A1_N(_06543_),
    .A2_N(_06551_),
    .B1(_06543_),
    .B2(_06551_),
    .X(_06552_));
 sky130_fd_sc_hd__a2bb2o_1 _22440_ (.A1_N(_06419_),
    .A2_N(_06552_),
    .B1(_06419_),
    .B2(_06552_),
    .X(_06553_));
 sky130_fd_sc_hd__a2bb2o_1 _22441_ (.A1_N(_06542_),
    .A2_N(_06553_),
    .B1(_06542_),
    .B2(_06553_),
    .X(_06554_));
 sky130_fd_sc_hd__o22a_1 _22442_ (.A1(_06295_),
    .A2(_06420_),
    .B1(_06412_),
    .B2(_06421_),
    .X(_06555_));
 sky130_fd_sc_hd__or2_1 _22443_ (.A(_06554_),
    .B(_06555_),
    .X(_06556_));
 sky130_fd_sc_hd__a21bo_1 _22444_ (.A1(_06554_),
    .A2(_06555_),
    .B1_N(_06556_),
    .X(_06557_));
 sky130_fd_sc_hd__or2_2 _22445_ (.A(_06518_),
    .B(_06557_),
    .X(_06558_));
 sky130_fd_sc_hd__a21bo_1 _22446_ (.A1(_06518_),
    .A2(_06557_),
    .B1_N(_06558_),
    .X(_06559_));
 sky130_vsdinv _22447_ (.A(_06559_),
    .Y(_06560_));
 sky130_fd_sc_hd__a22o_1 _22448_ (.A1(_06426_),
    .A2(_06559_),
    .B1(_06427_),
    .B2(_06560_),
    .X(_06561_));
 sky130_fd_sc_hd__o22a_1 _22449_ (.A1(_06493_),
    .A2(_06494_),
    .B1(_06472_),
    .B2(_06495_),
    .X(_06562_));
 sky130_fd_sc_hd__a21oi_2 _22450_ (.A1(_06444_),
    .A2(_06446_),
    .B1(_06443_),
    .Y(_06563_));
 sky130_fd_sc_hd__clkbuf_2 _22451_ (.A(_05925_),
    .X(_06564_));
 sky130_fd_sc_hd__buf_1 _22452_ (.A(_06449_),
    .X(_06565_));
 sky130_fd_sc_hd__clkbuf_2 _22453_ (.A(_06565_),
    .X(_06566_));
 sky130_fd_sc_hd__buf_2 _22454_ (.A(_06566_),
    .X(_06567_));
 sky130_fd_sc_hd__o22a_1 _22455_ (.A1(_06564_),
    .A2(_06439_),
    .B1(_06436_),
    .B2(_06567_),
    .X(_06568_));
 sky130_fd_sc_hd__and4_1 _22456_ (.A(_06441_),
    .B(_13561_),
    .C(_06442_),
    .D(_13557_),
    .X(_06569_));
 sky130_fd_sc_hd__nor2_2 _22457_ (.A(_06568_),
    .B(_06569_),
    .Y(_06570_));
 sky130_fd_sc_hd__nor2_2 _22458_ (.A(_06445_),
    .B(_06435_),
    .Y(_06571_));
 sky130_fd_sc_hd__a2bb2o_1 _22459_ (.A1_N(_06570_),
    .A2_N(_06571_),
    .B1(_06570_),
    .B2(_06571_),
    .X(_06572_));
 sky130_vsdinv _22460_ (.A(\pcpi_mul.rs1[20] ),
    .Y(_06573_));
 sky130_fd_sc_hd__buf_1 _22461_ (.A(_06573_),
    .X(_06574_));
 sky130_fd_sc_hd__buf_1 _22462_ (.A(_06574_),
    .X(_06575_));
 sky130_fd_sc_hd__buf_2 _22463_ (.A(_06575_),
    .X(_06576_));
 sky130_fd_sc_hd__or2_1 _22464_ (.A(_06448_),
    .B(_06576_),
    .X(_06577_));
 sky130_fd_sc_hd__buf_2 _22465_ (.A(_05839_),
    .X(_06578_));
 sky130_fd_sc_hd__buf_2 _22466_ (.A(_05842_),
    .X(_06579_));
 sky130_fd_sc_hd__buf_1 _22467_ (.A(_06138_),
    .X(_06580_));
 sky130_fd_sc_hd__clkbuf_2 _22468_ (.A(_06580_),
    .X(_06581_));
 sky130_fd_sc_hd__o22a_1 _22469_ (.A1(_06578_),
    .A2(_06457_),
    .B1(_06579_),
    .B2(_06581_),
    .X(_06582_));
 sky130_fd_sc_hd__buf_1 _22470_ (.A(\pcpi_mul.rs1[16] ),
    .X(_06583_));
 sky130_fd_sc_hd__buf_1 _22471_ (.A(_06583_),
    .X(_06584_));
 sky130_fd_sc_hd__and4_1 _22472_ (.A(_06459_),
    .B(_06463_),
    .C(_06461_),
    .D(_06584_),
    .X(_06585_));
 sky130_fd_sc_hd__or2_1 _22473_ (.A(_06582_),
    .B(_06585_),
    .X(_06586_));
 sky130_fd_sc_hd__a2bb2o_1 _22474_ (.A1_N(_06577_),
    .A2_N(_06586_),
    .B1(_06577_),
    .B2(_06586_),
    .X(_06587_));
 sky130_fd_sc_hd__o21ba_1 _22475_ (.A1(_06453_),
    .A2(_06465_),
    .B1_N(_06464_),
    .X(_06588_));
 sky130_fd_sc_hd__a2bb2o_1 _22476_ (.A1_N(_06587_),
    .A2_N(_06588_),
    .B1(_06587_),
    .B2(_06588_),
    .X(_06589_));
 sky130_fd_sc_hd__a2bb2o_1 _22477_ (.A1_N(_06572_),
    .A2_N(_06589_),
    .B1(_06572_),
    .B2(_06589_),
    .X(_06590_));
 sky130_fd_sc_hd__o22a_1 _22478_ (.A1(_06466_),
    .A2(_06467_),
    .B1(_06447_),
    .B2(_06468_),
    .X(_06591_));
 sky130_fd_sc_hd__a2bb2o_1 _22479_ (.A1_N(_06590_),
    .A2_N(_06591_),
    .B1(_06590_),
    .B2(_06591_),
    .X(_06592_));
 sky130_fd_sc_hd__a2bb2o_1 _22480_ (.A1_N(_06563_),
    .A2_N(_06592_),
    .B1(_06563_),
    .B2(_06592_),
    .X(_06593_));
 sky130_fd_sc_hd__o22a_1 _22481_ (.A1(_06476_),
    .A2(_06489_),
    .B1(_06475_),
    .B2(_06490_),
    .X(_06594_));
 sky130_fd_sc_hd__o22a_1 _22482_ (.A1(_06409_),
    .A2(_06410_),
    .B1(_06404_),
    .B2(_06411_),
    .X(_06595_));
 sky130_fd_sc_hd__o21ba_2 _22483_ (.A1(_06480_),
    .A2(_06488_),
    .B1_N(_06487_),
    .X(_06596_));
 sky130_fd_sc_hd__o21ba_1 _22484_ (.A1(_06400_),
    .A2(_06403_),
    .B1_N(_06402_),
    .X(_06597_));
 sky130_fd_sc_hd__clkbuf_2 _22485_ (.A(_05942_),
    .X(_06598_));
 sky130_fd_sc_hd__clkbuf_2 _22486_ (.A(_06598_),
    .X(_06599_));
 sky130_fd_sc_hd__or2_1 _22487_ (.A(_06477_),
    .B(_06599_),
    .X(_06600_));
 sky130_fd_sc_hd__o22a_1 _22488_ (.A1(_06481_),
    .A2(_05927_),
    .B1(_06483_),
    .B2(_06028_),
    .X(_06601_));
 sky130_fd_sc_hd__buf_1 _22489_ (.A(_13581_),
    .X(_06602_));
 sky130_fd_sc_hd__buf_1 _22490_ (.A(_13578_),
    .X(_06603_));
 sky130_fd_sc_hd__and4_1 _22491_ (.A(_13148_),
    .B(_06602_),
    .C(_13154_),
    .D(_06603_),
    .X(_06604_));
 sky130_fd_sc_hd__or2_1 _22492_ (.A(_06601_),
    .B(_06604_),
    .X(_06605_));
 sky130_fd_sc_hd__a2bb2o_2 _22493_ (.A1_N(_06600_),
    .A2_N(_06605_),
    .B1(_06600_),
    .B2(_06605_),
    .X(_06606_));
 sky130_fd_sc_hd__a2bb2o_1 _22494_ (.A1_N(_06597_),
    .A2_N(_06606_),
    .B1(_06597_),
    .B2(_06606_),
    .X(_06607_));
 sky130_fd_sc_hd__a2bb2o_1 _22495_ (.A1_N(_06596_),
    .A2_N(_06607_),
    .B1(_06596_),
    .B2(_06607_),
    .X(_06608_));
 sky130_fd_sc_hd__a2bb2o_1 _22496_ (.A1_N(_06595_),
    .A2_N(_06608_),
    .B1(_06595_),
    .B2(_06608_),
    .X(_06609_));
 sky130_fd_sc_hd__a2bb2o_1 _22497_ (.A1_N(_06594_),
    .A2_N(_06609_),
    .B1(_06594_),
    .B2(_06609_),
    .X(_06610_));
 sky130_fd_sc_hd__o22a_2 _22498_ (.A1(_06474_),
    .A2(_06491_),
    .B1(_06473_),
    .B2(_06492_),
    .X(_06611_));
 sky130_fd_sc_hd__a2bb2o_1 _22499_ (.A1_N(_06610_),
    .A2_N(_06611_),
    .B1(_06610_),
    .B2(_06611_),
    .X(_06612_));
 sky130_fd_sc_hd__a2bb2o_2 _22500_ (.A1_N(_06593_),
    .A2_N(_06612_),
    .B1(_06593_),
    .B2(_06612_),
    .X(_06613_));
 sky130_fd_sc_hd__a2bb2o_1 _22501_ (.A1_N(_06424_),
    .A2_N(_06613_),
    .B1(_06424_),
    .B2(_06613_),
    .X(_06614_));
 sky130_fd_sc_hd__a2bb2o_1 _22502_ (.A1_N(_06562_),
    .A2_N(_06614_),
    .B1(_06562_),
    .B2(_06614_),
    .X(_06615_));
 sky130_fd_sc_hd__a2bb2o_1 _22503_ (.A1_N(_06561_),
    .A2_N(_06615_),
    .B1(_06561_),
    .B2(_06615_),
    .X(_06616_));
 sky130_fd_sc_hd__o22a_1 _22504_ (.A1(_06321_),
    .A2(_06429_),
    .B1(_06430_),
    .B2(_06498_),
    .X(_06617_));
 sky130_fd_sc_hd__a2bb2o_1 _22505_ (.A1_N(_06616_),
    .A2_N(_06617_),
    .B1(_06616_),
    .B2(_06617_),
    .X(_06618_));
 sky130_fd_sc_hd__a2bb2o_1 _22506_ (.A1_N(_06512_),
    .A2_N(_06618_),
    .B1(_06512_),
    .B2(_06618_),
    .X(_06619_));
 sky130_fd_sc_hd__o22a_1 _22507_ (.A1(_06371_),
    .A2(_06499_),
    .B1(_06387_),
    .B2(_06500_),
    .X(_06620_));
 sky130_fd_sc_hd__a2bb2o_1 _22508_ (.A1_N(_06619_),
    .A2_N(_06620_),
    .B1(_06619_),
    .B2(_06620_),
    .X(_06621_));
 sky130_fd_sc_hd__a2bb2o_1 _22509_ (.A1_N(_06386_),
    .A2_N(_06621_),
    .B1(_06386_),
    .B2(_06621_),
    .X(_06622_));
 sky130_fd_sc_hd__o22a_1 _22510_ (.A1(_06501_),
    .A2(_06502_),
    .B1(_06281_),
    .B2(_06503_),
    .X(_06623_));
 sky130_fd_sc_hd__or2_2 _22511_ (.A(_06622_),
    .B(_06623_),
    .X(_06624_));
 sky130_fd_sc_hd__a21bo_1 _22512_ (.A1(_06622_),
    .A2(_06623_),
    .B1_N(_06624_),
    .X(_06625_));
 sky130_fd_sc_hd__clkbuf_2 _22513_ (.A(_06625_),
    .X(_06626_));
 sky130_fd_sc_hd__or2_1 _22514_ (.A(_06380_),
    .B(_06507_),
    .X(_06627_));
 sky130_fd_sc_hd__or3_1 _22515_ (.A(_06182_),
    .B(_06277_),
    .C(_06627_),
    .X(_06628_));
 sky130_fd_sc_hd__o221a_1 _22516_ (.A1(_06379_),
    .A2(_06505_),
    .B1(_06381_),
    .B2(_06627_),
    .C1(_06506_),
    .X(_06629_));
 sky130_fd_sc_hd__o21ai_1 _22517_ (.A1(_06081_),
    .A2(_06628_),
    .B1(_06629_),
    .Y(_06630_));
 sky130_vsdinv _22518_ (.A(_06630_),
    .Y(_06631_));
 sky130_vsdinv _22519_ (.A(_06626_),
    .Y(_06632_));
 sky130_fd_sc_hd__o22a_4 _22520_ (.A1(_06626_),
    .A2(_06631_),
    .B1(_06632_),
    .B2(_06630_),
    .X(_02639_));
 sky130_fd_sc_hd__o22a_1 _22521_ (.A1(_06619_),
    .A2(_06620_),
    .B1(_06386_),
    .B2(_06621_),
    .X(_06633_));
 sky130_fd_sc_hd__o22a_1 _22522_ (.A1(_06424_),
    .A2(_06613_),
    .B1(_06562_),
    .B2(_06614_),
    .X(_06634_));
 sky130_fd_sc_hd__o22a_2 _22523_ (.A1(_06590_),
    .A2(_06591_),
    .B1(_06563_),
    .B2(_06592_),
    .X(_06635_));
 sky130_fd_sc_hd__or2_1 _22524_ (.A(_06634_),
    .B(_06635_),
    .X(_06636_));
 sky130_fd_sc_hd__a21bo_1 _22525_ (.A1(_06634_),
    .A2(_06635_),
    .B1_N(_06636_),
    .X(_06637_));
 sky130_fd_sc_hd__o22a_1 _22526_ (.A1(_06610_),
    .A2(_06611_),
    .B1(_06593_),
    .B2(_06612_),
    .X(_06638_));
 sky130_fd_sc_hd__a21oi_2 _22527_ (.A1(_06570_),
    .A2(_06571_),
    .B1(_06569_),
    .Y(_06639_));
 sky130_fd_sc_hd__buf_1 _22528_ (.A(_06573_),
    .X(_06640_));
 sky130_fd_sc_hd__buf_2 _22529_ (.A(_06640_),
    .X(_06641_));
 sky130_fd_sc_hd__buf_4 _22530_ (.A(_06641_),
    .X(_06642_));
 sky130_fd_sc_hd__o22a_1 _22531_ (.A1(_06564_),
    .A2(_06567_),
    .B1(_06436_),
    .B2(_06642_),
    .X(_06643_));
 sky130_fd_sc_hd__and4_1 _22532_ (.A(_06441_),
    .B(_13557_),
    .C(_06442_),
    .D(_13554_),
    .X(_06644_));
 sky130_fd_sc_hd__nor2_2 _22533_ (.A(_06643_),
    .B(_06644_),
    .Y(_06645_));
 sky130_fd_sc_hd__nor2_2 _22534_ (.A(_06445_),
    .B(_06439_),
    .Y(_06646_));
 sky130_fd_sc_hd__a2bb2o_1 _22535_ (.A1_N(_06645_),
    .A2_N(_06646_),
    .B1(_06645_),
    .B2(_06646_),
    .X(_06647_));
 sky130_vsdinv _22536_ (.A(\pcpi_mul.rs1[21] ),
    .Y(_06648_));
 sky130_fd_sc_hd__buf_1 _22537_ (.A(_06648_),
    .X(_06649_));
 sky130_fd_sc_hd__clkbuf_2 _22538_ (.A(_06649_),
    .X(_06650_));
 sky130_fd_sc_hd__clkbuf_4 _22539_ (.A(_06650_),
    .X(_06651_));
 sky130_fd_sc_hd__or2_1 _22540_ (.A(_06448_),
    .B(_06651_),
    .X(_06652_));
 sky130_fd_sc_hd__o22a_1 _22541_ (.A1(_06578_),
    .A2(_06581_),
    .B1(_06579_),
    .B2(_06227_),
    .X(_06653_));
 sky130_fd_sc_hd__buf_1 _22542_ (.A(_13563_),
    .X(_06654_));
 sky130_fd_sc_hd__and4_1 _22543_ (.A(_06459_),
    .B(_06584_),
    .C(_06461_),
    .D(_06654_),
    .X(_06655_));
 sky130_fd_sc_hd__or2_1 _22544_ (.A(_06653_),
    .B(_06655_),
    .X(_06656_));
 sky130_fd_sc_hd__a2bb2o_1 _22545_ (.A1_N(_06652_),
    .A2_N(_06656_),
    .B1(_06652_),
    .B2(_06656_),
    .X(_06657_));
 sky130_fd_sc_hd__o21ba_1 _22546_ (.A1(_06577_),
    .A2(_06586_),
    .B1_N(_06585_),
    .X(_06658_));
 sky130_fd_sc_hd__a2bb2o_1 _22547_ (.A1_N(_06657_),
    .A2_N(_06658_),
    .B1(_06657_),
    .B2(_06658_),
    .X(_06659_));
 sky130_fd_sc_hd__a2bb2o_1 _22548_ (.A1_N(_06647_),
    .A2_N(_06659_),
    .B1(_06647_),
    .B2(_06659_),
    .X(_06660_));
 sky130_fd_sc_hd__o22a_1 _22549_ (.A1(_06587_),
    .A2(_06588_),
    .B1(_06572_),
    .B2(_06589_),
    .X(_06661_));
 sky130_fd_sc_hd__a2bb2o_1 _22550_ (.A1_N(_06660_),
    .A2_N(_06661_),
    .B1(_06660_),
    .B2(_06661_),
    .X(_06662_));
 sky130_fd_sc_hd__a2bb2o_2 _22551_ (.A1_N(_06639_),
    .A2_N(_06662_),
    .B1(_06639_),
    .B2(_06662_),
    .X(_06663_));
 sky130_fd_sc_hd__o22a_1 _22552_ (.A1(_06597_),
    .A2(_06606_),
    .B1(_06596_),
    .B2(_06607_),
    .X(_06664_));
 sky130_fd_sc_hd__o22a_1 _22553_ (.A1(_06539_),
    .A2(_06540_),
    .B1(_06531_),
    .B2(_06541_),
    .X(_06665_));
 sky130_fd_sc_hd__o21ba_1 _22554_ (.A1(_06600_),
    .A2(_06605_),
    .B1_N(_06604_),
    .X(_06666_));
 sky130_fd_sc_hd__o21ba_1 _22555_ (.A1(_06521_),
    .A2(_06530_),
    .B1_N(_06529_),
    .X(_06667_));
 sky130_fd_sc_hd__buf_1 _22556_ (.A(_06039_),
    .X(_06668_));
 sky130_fd_sc_hd__buf_2 _22557_ (.A(_06668_),
    .X(_06669_));
 sky130_fd_sc_hd__or2_1 _22558_ (.A(_06477_),
    .B(_06669_),
    .X(_06670_));
 sky130_fd_sc_hd__buf_2 _22559_ (.A(_05864_),
    .X(_06671_));
 sky130_fd_sc_hd__o22a_1 _22560_ (.A1(_06671_),
    .A2(_06478_),
    .B1(_06483_),
    .B2(_06129_),
    .X(_06672_));
 sky130_fd_sc_hd__buf_1 _22561_ (.A(_13574_),
    .X(_06673_));
 sky130_fd_sc_hd__and4_1 _22562_ (.A(_05870_),
    .B(_06603_),
    .C(_05871_),
    .D(_06673_),
    .X(_06674_));
 sky130_fd_sc_hd__or2_1 _22563_ (.A(_06672_),
    .B(_06674_),
    .X(_06675_));
 sky130_fd_sc_hd__a2bb2o_1 _22564_ (.A1_N(_06670_),
    .A2_N(_06675_),
    .B1(_06670_),
    .B2(_06675_),
    .X(_06676_));
 sky130_fd_sc_hd__a2bb2o_1 _22565_ (.A1_N(_06667_),
    .A2_N(_06676_),
    .B1(_06667_),
    .B2(_06676_),
    .X(_06677_));
 sky130_fd_sc_hd__a2bb2o_1 _22566_ (.A1_N(_06666_),
    .A2_N(_06677_),
    .B1(_06666_),
    .B2(_06677_),
    .X(_06678_));
 sky130_fd_sc_hd__a2bb2o_1 _22567_ (.A1_N(_06665_),
    .A2_N(_06678_),
    .B1(_06665_),
    .B2(_06678_),
    .X(_06679_));
 sky130_fd_sc_hd__a2bb2o_1 _22568_ (.A1_N(_06664_),
    .A2_N(_06679_),
    .B1(_06664_),
    .B2(_06679_),
    .X(_06680_));
 sky130_fd_sc_hd__o22a_1 _22569_ (.A1(_06595_),
    .A2(_06608_),
    .B1(_06594_),
    .B2(_06609_),
    .X(_06681_));
 sky130_fd_sc_hd__a2bb2o_1 _22570_ (.A1_N(_06680_),
    .A2_N(_06681_),
    .B1(_06680_),
    .B2(_06681_),
    .X(_06682_));
 sky130_fd_sc_hd__a2bb2o_1 _22571_ (.A1_N(_06663_),
    .A2_N(_06682_),
    .B1(_06663_),
    .B2(_06682_),
    .X(_06683_));
 sky130_fd_sc_hd__a2bb2o_1 _22572_ (.A1_N(_06556_),
    .A2_N(_06683_),
    .B1(_06556_),
    .B2(_06683_),
    .X(_06684_));
 sky130_fd_sc_hd__a2bb2o_1 _22573_ (.A1_N(_06638_),
    .A2_N(_06684_),
    .B1(_06638_),
    .B2(_06684_),
    .X(_06685_));
 sky130_vsdinv _22574_ (.A(\pcpi_mul.rs2[21] ),
    .Y(_06686_));
 sky130_fd_sc_hd__clkbuf_2 _22575_ (.A(_06686_),
    .X(_06687_));
 sky130_fd_sc_hd__clkbuf_4 _22576_ (.A(_06687_),
    .X(_06688_));
 sky130_fd_sc_hd__clkbuf_2 _22577_ (.A(_06688_),
    .X(_06689_));
 sky130_fd_sc_hd__buf_4 _22578_ (.A(_06689_),
    .X(_06690_));
 sky130_fd_sc_hd__or2_2 _22579_ (.A(_06690_),
    .B(_05152_),
    .X(_06691_));
 sky130_fd_sc_hd__or2_1 _22580_ (.A(_06283_),
    .B(_06011_),
    .X(_06692_));
 sky130_fd_sc_hd__o22a_1 _22581_ (.A1(_06514_),
    .A2(_05296_),
    .B1(_06388_),
    .B2(_06187_),
    .X(_06693_));
 sky130_fd_sc_hd__buf_1 _22582_ (.A(\pcpi_mul.rs2[20] ),
    .X(_06694_));
 sky130_fd_sc_hd__buf_1 _22583_ (.A(_05647_),
    .X(_06695_));
 sky130_fd_sc_hd__and4_1 _22584_ (.A(_06694_),
    .B(_06695_),
    .C(_13110_),
    .D(_05346_),
    .X(_06696_));
 sky130_fd_sc_hd__or2_1 _22585_ (.A(_06693_),
    .B(_06696_),
    .X(_06697_));
 sky130_fd_sc_hd__a2bb2o_2 _22586_ (.A1_N(_06692_),
    .A2_N(_06697_),
    .B1(_06692_),
    .B2(_06697_),
    .X(_06698_));
 sky130_fd_sc_hd__nor2_2 _22587_ (.A(_06691_),
    .B(_06698_),
    .Y(_06699_));
 sky130_fd_sc_hd__a21o_1 _22588_ (.A1(_06691_),
    .A2(_06698_),
    .B1(_06699_),
    .X(_06700_));
 sky130_fd_sc_hd__o22a_1 _22589_ (.A1(_06419_),
    .A2(_06552_),
    .B1(_06542_),
    .B2(_06553_),
    .X(_06701_));
 sky130_fd_sc_hd__buf_2 _22590_ (.A(_05819_),
    .X(_06702_));
 sky130_fd_sc_hd__or2_1 _22591_ (.A(_06519_),
    .B(_06702_),
    .X(_06703_));
 sky130_fd_sc_hd__clkbuf_2 _22592_ (.A(_05667_),
    .X(_06704_));
 sky130_fd_sc_hd__o22a_1 _22593_ (.A1(_06300_),
    .A2(_06042_),
    .B1(_06523_),
    .B2(_06704_),
    .X(_06705_));
 sky130_fd_sc_hd__and4_1 _22594_ (.A(_06525_),
    .B(_06528_),
    .C(_06527_),
    .D(_06144_),
    .X(_06706_));
 sky130_fd_sc_hd__or2_1 _22595_ (.A(_06705_),
    .B(_06706_),
    .X(_06707_));
 sky130_fd_sc_hd__a2bb2o_2 _22596_ (.A1_N(_06703_),
    .A2_N(_06707_),
    .B1(_06703_),
    .B2(_06707_),
    .X(_06708_));
 sky130_fd_sc_hd__or2_1 _22597_ (.A(_05708_),
    .B(_06298_),
    .X(_06709_));
 sky130_fd_sc_hd__buf_2 _22598_ (.A(_06013_),
    .X(_06710_));
 sky130_fd_sc_hd__o22a_1 _22599_ (.A1(_06710_),
    .A2(_05861_),
    .B1(_05788_),
    .B2(_05841_),
    .X(_06711_));
 sky130_fd_sc_hd__and4_1 _22600_ (.A(_13129_),
    .B(_06303_),
    .C(_13132_),
    .D(_06304_),
    .X(_06712_));
 sky130_fd_sc_hd__or2_1 _22601_ (.A(_06711_),
    .B(_06712_),
    .X(_06713_));
 sky130_fd_sc_hd__a2bb2o_1 _22602_ (.A1_N(_06709_),
    .A2_N(_06713_),
    .B1(_06709_),
    .B2(_06713_),
    .X(_06714_));
 sky130_fd_sc_hd__o21ba_1 _22603_ (.A1(_06532_),
    .A2(_06538_),
    .B1_N(_06537_),
    .X(_06715_));
 sky130_fd_sc_hd__a2bb2o_1 _22604_ (.A1_N(_06714_),
    .A2_N(_06715_),
    .B1(_06714_),
    .B2(_06715_),
    .X(_06716_));
 sky130_fd_sc_hd__a2bb2o_1 _22605_ (.A1_N(_06708_),
    .A2_N(_06716_),
    .B1(_06708_),
    .B2(_06716_),
    .X(_06717_));
 sky130_fd_sc_hd__o21ba_1 _22606_ (.A1(_06545_),
    .A2(_06549_),
    .B1_N(_06548_),
    .X(_06718_));
 sky130_fd_sc_hd__o21ba_1 _22607_ (.A1(_06513_),
    .A2(_06517_),
    .B1_N(_06516_),
    .X(_06719_));
 sky130_fd_sc_hd__or2_1 _22608_ (.A(_06095_),
    .B(_06308_),
    .X(_06720_));
 sky130_fd_sc_hd__o22a_1 _22609_ (.A1(_06546_),
    .A2(_06005_),
    .B1(_06092_),
    .B2(_05680_),
    .X(_06721_));
 sky130_fd_sc_hd__buf_1 _22610_ (.A(_13116_),
    .X(_06722_));
 sky130_fd_sc_hd__buf_1 _22611_ (.A(_13120_),
    .X(_06723_));
 sky130_fd_sc_hd__and4_1 _22612_ (.A(_06722_),
    .B(_05758_),
    .C(_06723_),
    .D(_06311_),
    .X(_06724_));
 sky130_fd_sc_hd__or2_1 _22613_ (.A(_06721_),
    .B(_06724_),
    .X(_06725_));
 sky130_fd_sc_hd__a2bb2o_1 _22614_ (.A1_N(_06720_),
    .A2_N(_06725_),
    .B1(_06720_),
    .B2(_06725_),
    .X(_06726_));
 sky130_fd_sc_hd__a2bb2o_1 _22615_ (.A1_N(_06719_),
    .A2_N(_06726_),
    .B1(_06719_),
    .B2(_06726_),
    .X(_06727_));
 sky130_fd_sc_hd__a2bb2o_1 _22616_ (.A1_N(_06718_),
    .A2_N(_06727_),
    .B1(_06718_),
    .B2(_06727_),
    .X(_06728_));
 sky130_fd_sc_hd__o22a_1 _22617_ (.A1(_06397_),
    .A2(_06550_),
    .B1(_06543_),
    .B2(_06551_),
    .X(_06729_));
 sky130_fd_sc_hd__a2bb2o_1 _22618_ (.A1_N(_06728_),
    .A2_N(_06729_),
    .B1(_06728_),
    .B2(_06729_),
    .X(_06730_));
 sky130_fd_sc_hd__a2bb2o_1 _22619_ (.A1_N(_06717_),
    .A2_N(_06730_),
    .B1(_06717_),
    .B2(_06730_),
    .X(_06731_));
 sky130_fd_sc_hd__or2_2 _22620_ (.A(_06701_),
    .B(_06731_),
    .X(_06732_));
 sky130_fd_sc_hd__a21bo_1 _22621_ (.A1(_06701_),
    .A2(_06731_),
    .B1_N(_06732_),
    .X(_06733_));
 sky130_fd_sc_hd__or2_1 _22622_ (.A(_06700_),
    .B(_06733_),
    .X(_06734_));
 sky130_fd_sc_hd__a21bo_1 _22623_ (.A1(_06700_),
    .A2(_06733_),
    .B1_N(_06734_),
    .X(_06735_));
 sky130_fd_sc_hd__a2bb2o_1 _22624_ (.A1_N(_06558_),
    .A2_N(_06735_),
    .B1(_06558_),
    .B2(_06735_),
    .X(_06736_));
 sky130_fd_sc_hd__a2bb2o_2 _22625_ (.A1_N(_06685_),
    .A2_N(_06736_),
    .B1(_06685_),
    .B2(_06736_),
    .X(_06737_));
 sky130_fd_sc_hd__o22a_1 _22626_ (.A1(_06426_),
    .A2(_06559_),
    .B1(_06561_),
    .B2(_06615_),
    .X(_06738_));
 sky130_fd_sc_hd__a2bb2o_1 _22627_ (.A1_N(_06737_),
    .A2_N(_06738_),
    .B1(_06737_),
    .B2(_06738_),
    .X(_06739_));
 sky130_fd_sc_hd__a2bb2o_1 _22628_ (.A1_N(_06637_),
    .A2_N(_06739_),
    .B1(_06637_),
    .B2(_06739_),
    .X(_06740_));
 sky130_fd_sc_hd__o22a_1 _22629_ (.A1(_06616_),
    .A2(_06617_),
    .B1(_06512_),
    .B2(_06618_),
    .X(_06741_));
 sky130_fd_sc_hd__a2bb2o_1 _22630_ (.A1_N(_06740_),
    .A2_N(_06741_),
    .B1(_06740_),
    .B2(_06741_),
    .X(_06742_));
 sky130_fd_sc_hd__a2bb2o_1 _22631_ (.A1_N(_06511_),
    .A2_N(_06742_),
    .B1(_06511_),
    .B2(_06742_),
    .X(_06743_));
 sky130_fd_sc_hd__or2_1 _22632_ (.A(_06633_),
    .B(_06743_),
    .X(_06744_));
 sky130_fd_sc_hd__a21bo_1 _22633_ (.A1(_06633_),
    .A2(_06743_),
    .B1_N(_06744_),
    .X(_06745_));
 sky130_fd_sc_hd__o21ai_2 _22634_ (.A1(_06626_),
    .A2(_06631_),
    .B1(_06624_),
    .Y(_06746_));
 sky130_fd_sc_hd__a2bb2o_4 _22635_ (.A1_N(_06745_),
    .A2_N(_06746_),
    .B1(_06745_),
    .B2(_06746_),
    .X(_02640_));
 sky130_fd_sc_hd__o22a_1 _22636_ (.A1(_06556_),
    .A2(_06683_),
    .B1(_06638_),
    .B2(_06684_),
    .X(_06747_));
 sky130_fd_sc_hd__o22a_1 _22637_ (.A1(_06660_),
    .A2(_06661_),
    .B1(_06639_),
    .B2(_06662_),
    .X(_06748_));
 sky130_fd_sc_hd__or2_1 _22638_ (.A(_06747_),
    .B(_06748_),
    .X(_06749_));
 sky130_fd_sc_hd__a21bo_1 _22639_ (.A1(_06747_),
    .A2(_06748_),
    .B1_N(_06749_),
    .X(_06750_));
 sky130_fd_sc_hd__o22a_1 _22640_ (.A1(_06680_),
    .A2(_06681_),
    .B1(_06663_),
    .B2(_06682_),
    .X(_06751_));
 sky130_fd_sc_hd__a21oi_2 _22641_ (.A1(_06645_),
    .A2(_06646_),
    .B1(_06644_),
    .Y(_06752_));
 sky130_fd_sc_hd__clkbuf_2 _22642_ (.A(_05306_),
    .X(_06753_));
 sky130_fd_sc_hd__buf_1 _22643_ (.A(_06649_),
    .X(_06754_));
 sky130_fd_sc_hd__clkbuf_4 _22644_ (.A(_06754_),
    .X(_06755_));
 sky130_fd_sc_hd__o22a_1 _22645_ (.A1(_06564_),
    .A2(_06576_),
    .B1(_06753_),
    .B2(_06755_),
    .X(_06756_));
 sky130_fd_sc_hd__and4_1 _22646_ (.A(_06441_),
    .B(_13554_),
    .C(_06442_),
    .D(_13551_),
    .X(_06757_));
 sky130_fd_sc_hd__nor2_2 _22647_ (.A(_06756_),
    .B(_06757_),
    .Y(_06758_));
 sky130_fd_sc_hd__nor2_2 _22648_ (.A(_06445_),
    .B(_06567_),
    .Y(_06759_));
 sky130_fd_sc_hd__a2bb2o_1 _22649_ (.A1_N(_06758_),
    .A2_N(_06759_),
    .B1(_06758_),
    .B2(_06759_),
    .X(_06760_));
 sky130_vsdinv _22650_ (.A(\pcpi_mul.rs1[22] ),
    .Y(_06761_));
 sky130_fd_sc_hd__clkbuf_2 _22651_ (.A(_06761_),
    .X(_06762_));
 sky130_fd_sc_hd__buf_2 _22652_ (.A(_06762_),
    .X(_06763_));
 sky130_fd_sc_hd__or2_1 _22653_ (.A(_05142_),
    .B(_06763_),
    .X(_06764_));
 sky130_fd_sc_hd__clkbuf_2 _22654_ (.A(_06337_),
    .X(_06765_));
 sky130_fd_sc_hd__clkbuf_2 _22655_ (.A(_06765_),
    .X(_06766_));
 sky130_fd_sc_hd__o22a_1 _22656_ (.A1(_06578_),
    .A2(_06434_),
    .B1(_06579_),
    .B2(_06766_),
    .X(_06767_));
 sky130_fd_sc_hd__buf_1 _22657_ (.A(_13563_),
    .X(_06768_));
 sky130_fd_sc_hd__buf_1 _22658_ (.A(_13559_),
    .X(_06769_));
 sky130_fd_sc_hd__and4_1 _22659_ (.A(_13161_),
    .B(_06768_),
    .C(_13167_),
    .D(_06769_),
    .X(_06770_));
 sky130_fd_sc_hd__or2_1 _22660_ (.A(_06767_),
    .B(_06770_),
    .X(_06771_));
 sky130_fd_sc_hd__a2bb2o_1 _22661_ (.A1_N(_06764_),
    .A2_N(_06771_),
    .B1(_06764_),
    .B2(_06771_),
    .X(_06772_));
 sky130_fd_sc_hd__o21ba_1 _22662_ (.A1(_06652_),
    .A2(_06656_),
    .B1_N(_06655_),
    .X(_06773_));
 sky130_fd_sc_hd__a2bb2o_1 _22663_ (.A1_N(_06772_),
    .A2_N(_06773_),
    .B1(_06772_),
    .B2(_06773_),
    .X(_06774_));
 sky130_fd_sc_hd__a2bb2o_1 _22664_ (.A1_N(_06760_),
    .A2_N(_06774_),
    .B1(_06760_),
    .B2(_06774_),
    .X(_06775_));
 sky130_fd_sc_hd__o22a_1 _22665_ (.A1(_06657_),
    .A2(_06658_),
    .B1(_06647_),
    .B2(_06659_),
    .X(_06776_));
 sky130_fd_sc_hd__a2bb2o_1 _22666_ (.A1_N(_06775_),
    .A2_N(_06776_),
    .B1(_06775_),
    .B2(_06776_),
    .X(_06777_));
 sky130_fd_sc_hd__a2bb2o_1 _22667_ (.A1_N(_06752_),
    .A2_N(_06777_),
    .B1(_06752_),
    .B2(_06777_),
    .X(_06778_));
 sky130_fd_sc_hd__o22a_2 _22668_ (.A1(_06667_),
    .A2(_06676_),
    .B1(_06666_),
    .B2(_06677_),
    .X(_06779_));
 sky130_fd_sc_hd__o22a_1 _22669_ (.A1(_06714_),
    .A2(_06715_),
    .B1(_06708_),
    .B2(_06716_),
    .X(_06780_));
 sky130_fd_sc_hd__o21ba_1 _22670_ (.A1(_06670_),
    .A2(_06675_),
    .B1_N(_06674_),
    .X(_06781_));
 sky130_fd_sc_hd__o21ba_1 _22671_ (.A1(_06703_),
    .A2(_06707_),
    .B1_N(_06706_),
    .X(_06782_));
 sky130_fd_sc_hd__buf_2 _22672_ (.A(_06326_),
    .X(_06783_));
 sky130_fd_sc_hd__or2_1 _22673_ (.A(_05460_),
    .B(_06783_),
    .X(_06784_));
 sky130_fd_sc_hd__o22a_1 _22674_ (.A1(_06671_),
    .A2(_06598_),
    .B1(_05457_),
    .B2(_06668_),
    .X(_06785_));
 sky130_fd_sc_hd__buf_1 _22675_ (.A(_13569_),
    .X(_06786_));
 sky130_fd_sc_hd__and4_1 _22676_ (.A(_05870_),
    .B(_06673_),
    .C(_05871_),
    .D(_06786_),
    .X(_06787_));
 sky130_fd_sc_hd__or2_1 _22677_ (.A(_06785_),
    .B(_06787_),
    .X(_06788_));
 sky130_fd_sc_hd__a2bb2o_1 _22678_ (.A1_N(_06784_),
    .A2_N(_06788_),
    .B1(_06784_),
    .B2(_06788_),
    .X(_06789_));
 sky130_fd_sc_hd__a2bb2o_1 _22679_ (.A1_N(_06782_),
    .A2_N(_06789_),
    .B1(_06782_),
    .B2(_06789_),
    .X(_06790_));
 sky130_fd_sc_hd__a2bb2o_1 _22680_ (.A1_N(_06781_),
    .A2_N(_06790_),
    .B1(_06781_),
    .B2(_06790_),
    .X(_06791_));
 sky130_fd_sc_hd__a2bb2o_1 _22681_ (.A1_N(_06780_),
    .A2_N(_06791_),
    .B1(_06780_),
    .B2(_06791_),
    .X(_06792_));
 sky130_fd_sc_hd__a2bb2o_1 _22682_ (.A1_N(_06779_),
    .A2_N(_06792_),
    .B1(_06779_),
    .B2(_06792_),
    .X(_06793_));
 sky130_fd_sc_hd__o22a_1 _22683_ (.A1(_06665_),
    .A2(_06678_),
    .B1(_06664_),
    .B2(_06679_),
    .X(_06794_));
 sky130_fd_sc_hd__a2bb2o_1 _22684_ (.A1_N(_06793_),
    .A2_N(_06794_),
    .B1(_06793_),
    .B2(_06794_),
    .X(_06795_));
 sky130_fd_sc_hd__a2bb2o_1 _22685_ (.A1_N(_06778_),
    .A2_N(_06795_),
    .B1(_06778_),
    .B2(_06795_),
    .X(_06796_));
 sky130_fd_sc_hd__a2bb2o_1 _22686_ (.A1_N(_06732_),
    .A2_N(_06796_),
    .B1(_06732_),
    .B2(_06796_),
    .X(_06797_));
 sky130_fd_sc_hd__a2bb2o_1 _22687_ (.A1_N(_06751_),
    .A2_N(_06797_),
    .B1(_06751_),
    .B2(_06797_),
    .X(_06798_));
 sky130_vsdinv _22688_ (.A(\pcpi_mul.rs2[22] ),
    .Y(_06799_));
 sky130_fd_sc_hd__buf_1 _22689_ (.A(_06799_),
    .X(_06800_));
 sky130_fd_sc_hd__clkbuf_4 _22690_ (.A(_06800_),
    .X(_06801_));
 sky130_fd_sc_hd__clkbuf_2 _22691_ (.A(_06801_),
    .X(_06802_));
 sky130_fd_sc_hd__clkbuf_4 _22692_ (.A(_06687_),
    .X(_06803_));
 sky130_fd_sc_hd__o22a_1 _22693_ (.A1(_06802_),
    .A2(_05150_),
    .B1(_06803_),
    .B2(_05298_),
    .X(_06804_));
 sky130_fd_sc_hd__clkbuf_2 _22694_ (.A(_06799_),
    .X(_06805_));
 sky130_fd_sc_hd__clkbuf_2 _22695_ (.A(_06805_),
    .X(_06806_));
 sky130_fd_sc_hd__or4_4 _22696_ (.A(_06806_),
    .B(_05325_),
    .C(_06687_),
    .D(_05319_),
    .X(_06807_));
 sky130_fd_sc_hd__or2b_1 _22697_ (.A(_06804_),
    .B_N(_06807_),
    .X(_06808_));
 sky130_fd_sc_hd__or2_1 _22698_ (.A(_06396_),
    .B(_05799_),
    .X(_06809_));
 sky130_fd_sc_hd__clkbuf_2 _22699_ (.A(_06514_),
    .X(_06810_));
 sky130_fd_sc_hd__o22a_1 _22700_ (.A1(_06810_),
    .A2(_05645_),
    .B1(_06394_),
    .B2(_05803_),
    .X(_06811_));
 sky130_fd_sc_hd__and4_1 _22701_ (.A(_06694_),
    .B(_06115_),
    .C(_13110_),
    .D(_05808_),
    .X(_06812_));
 sky130_fd_sc_hd__or2_1 _22702_ (.A(_06811_),
    .B(_06812_),
    .X(_06813_));
 sky130_fd_sc_hd__a2bb2o_1 _22703_ (.A1_N(_06809_),
    .A2_N(_06813_),
    .B1(_06809_),
    .B2(_06813_),
    .X(_06814_));
 sky130_fd_sc_hd__or2_1 _22704_ (.A(_06808_),
    .B(_06814_),
    .X(_06815_));
 sky130_fd_sc_hd__a21boi_1 _22705_ (.A1(_06808_),
    .A2(_06814_),
    .B1_N(_06815_),
    .Y(_06816_));
 sky130_fd_sc_hd__nand2_1 _22706_ (.A(_06699_),
    .B(_06816_),
    .Y(_06817_));
 sky130_fd_sc_hd__o21ai_1 _22707_ (.A1(_06699_),
    .A2(_06816_),
    .B1(_06817_),
    .Y(_06818_));
 sky130_fd_sc_hd__o22a_1 _22708_ (.A1(_06728_),
    .A2(_06729_),
    .B1(_06717_),
    .B2(_06730_),
    .X(_06819_));
 sky130_fd_sc_hd__clkbuf_2 _22709_ (.A(_05536_),
    .X(_06820_));
 sky130_fd_sc_hd__or2_1 _22710_ (.A(_06820_),
    .B(_06029_),
    .X(_06821_));
 sky130_fd_sc_hd__clkbuf_2 _22711_ (.A(_05714_),
    .X(_06822_));
 sky130_fd_sc_hd__o22a_1 _22712_ (.A1(_06822_),
    .A2(_06482_),
    .B1(_05588_),
    .B2(_06484_),
    .X(_06823_));
 sky130_fd_sc_hd__buf_1 _22713_ (.A(_06103_),
    .X(_06824_));
 sky130_fd_sc_hd__buf_1 _22714_ (.A(_06104_),
    .X(_06825_));
 sky130_fd_sc_hd__and4_1 _22715_ (.A(_06824_),
    .B(_06486_),
    .C(_06825_),
    .D(_06602_),
    .X(_06826_));
 sky130_fd_sc_hd__or2_1 _22716_ (.A(_06823_),
    .B(_06826_),
    .X(_06827_));
 sky130_fd_sc_hd__a2bb2o_2 _22717_ (.A1_N(_06821_),
    .A2_N(_06827_),
    .B1(_06821_),
    .B2(_06827_),
    .X(_06828_));
 sky130_fd_sc_hd__or2_1 _22718_ (.A(_05708_),
    .B(_06399_),
    .X(_06829_));
 sky130_fd_sc_hd__buf_2 _22719_ (.A(_06013_),
    .X(_06830_));
 sky130_fd_sc_hd__buf_2 _22720_ (.A(_05597_),
    .X(_06831_));
 sky130_fd_sc_hd__o22a_1 _22721_ (.A1(_06830_),
    .A2(_06831_),
    .B1(_05788_),
    .B2(_05946_),
    .X(_06832_));
 sky130_fd_sc_hd__and4_1 _22722_ (.A(_13129_),
    .B(_06304_),
    .C(_13132_),
    .D(_13591_),
    .X(_06833_));
 sky130_fd_sc_hd__or2_1 _22723_ (.A(_06832_),
    .B(_06833_),
    .X(_06834_));
 sky130_fd_sc_hd__a2bb2o_1 _22724_ (.A1_N(_06829_),
    .A2_N(_06834_),
    .B1(_06829_),
    .B2(_06834_),
    .X(_06835_));
 sky130_fd_sc_hd__o21ba_1 _22725_ (.A1(_06709_),
    .A2(_06713_),
    .B1_N(_06712_),
    .X(_06836_));
 sky130_fd_sc_hd__a2bb2o_1 _22726_ (.A1_N(_06835_),
    .A2_N(_06836_),
    .B1(_06835_),
    .B2(_06836_),
    .X(_06837_));
 sky130_fd_sc_hd__a2bb2o_1 _22727_ (.A1_N(_06828_),
    .A2_N(_06837_),
    .B1(_06828_),
    .B2(_06837_),
    .X(_06838_));
 sky130_fd_sc_hd__o21ba_1 _22728_ (.A1(_06720_),
    .A2(_06725_),
    .B1_N(_06724_),
    .X(_06839_));
 sky130_fd_sc_hd__o21ba_1 _22729_ (.A1(_06692_),
    .A2(_06697_),
    .B1_N(_06696_),
    .X(_06840_));
 sky130_fd_sc_hd__or2_1 _22730_ (.A(_06095_),
    .B(_06301_),
    .X(_06841_));
 sky130_fd_sc_hd__clkbuf_2 _22731_ (.A(_06546_),
    .X(_06842_));
 sky130_fd_sc_hd__o22a_1 _22732_ (.A1(_06842_),
    .A2(_05509_),
    .B1(_06092_),
    .B2(_05867_),
    .X(_06843_));
 sky130_fd_sc_hd__and4_1 _22733_ (.A(_06722_),
    .B(_06311_),
    .C(_06723_),
    .D(_13602_),
    .X(_06844_));
 sky130_fd_sc_hd__or2_1 _22734_ (.A(_06843_),
    .B(_06844_),
    .X(_06845_));
 sky130_fd_sc_hd__a2bb2o_1 _22735_ (.A1_N(_06841_),
    .A2_N(_06845_),
    .B1(_06841_),
    .B2(_06845_),
    .X(_06846_));
 sky130_fd_sc_hd__a2bb2o_1 _22736_ (.A1_N(_06840_),
    .A2_N(_06846_),
    .B1(_06840_),
    .B2(_06846_),
    .X(_06847_));
 sky130_fd_sc_hd__a2bb2o_1 _22737_ (.A1_N(_06839_),
    .A2_N(_06847_),
    .B1(_06839_),
    .B2(_06847_),
    .X(_06848_));
 sky130_fd_sc_hd__o22a_1 _22738_ (.A1(_06719_),
    .A2(_06726_),
    .B1(_06718_),
    .B2(_06727_),
    .X(_06849_));
 sky130_fd_sc_hd__a2bb2o_1 _22739_ (.A1_N(_06848_),
    .A2_N(_06849_),
    .B1(_06848_),
    .B2(_06849_),
    .X(_06850_));
 sky130_fd_sc_hd__a2bb2o_1 _22740_ (.A1_N(_06838_),
    .A2_N(_06850_),
    .B1(_06838_),
    .B2(_06850_),
    .X(_06851_));
 sky130_fd_sc_hd__or2_1 _22741_ (.A(_06819_),
    .B(_06851_),
    .X(_06852_));
 sky130_fd_sc_hd__a21bo_1 _22742_ (.A1(_06819_),
    .A2(_06851_),
    .B1_N(_06852_),
    .X(_06853_));
 sky130_fd_sc_hd__or2_2 _22743_ (.A(_06818_),
    .B(_06853_),
    .X(_06854_));
 sky130_fd_sc_hd__a21bo_1 _22744_ (.A1(_06818_),
    .A2(_06853_),
    .B1_N(_06854_),
    .X(_06855_));
 sky130_fd_sc_hd__a2bb2o_1 _22745_ (.A1_N(_06734_),
    .A2_N(_06855_),
    .B1(_06734_),
    .B2(_06855_),
    .X(_06856_));
 sky130_fd_sc_hd__a2bb2o_1 _22746_ (.A1_N(_06798_),
    .A2_N(_06856_),
    .B1(_06798_),
    .B2(_06856_),
    .X(_06857_));
 sky130_fd_sc_hd__o22a_1 _22747_ (.A1(_06558_),
    .A2(_06735_),
    .B1(_06685_),
    .B2(_06736_),
    .X(_06858_));
 sky130_fd_sc_hd__a2bb2o_1 _22748_ (.A1_N(_06857_),
    .A2_N(_06858_),
    .B1(_06857_),
    .B2(_06858_),
    .X(_06859_));
 sky130_fd_sc_hd__a2bb2o_2 _22749_ (.A1_N(_06750_),
    .A2_N(_06859_),
    .B1(_06750_),
    .B2(_06859_),
    .X(_06860_));
 sky130_fd_sc_hd__o22a_1 _22750_ (.A1(_06737_),
    .A2(_06738_),
    .B1(_06637_),
    .B2(_06739_),
    .X(_06861_));
 sky130_fd_sc_hd__a2bb2o_1 _22751_ (.A1_N(_06860_),
    .A2_N(_06861_),
    .B1(_06860_),
    .B2(_06861_),
    .X(_06862_));
 sky130_fd_sc_hd__a2bb2o_1 _22752_ (.A1_N(_06636_),
    .A2_N(_06862_),
    .B1(_06636_),
    .B2(_06862_),
    .X(_06863_));
 sky130_fd_sc_hd__o22a_1 _22753_ (.A1(_06740_),
    .A2(_06741_),
    .B1(_06511_),
    .B2(_06742_),
    .X(_06864_));
 sky130_fd_sc_hd__or2_1 _22754_ (.A(_06863_),
    .B(_06864_),
    .X(_06865_));
 sky130_fd_sc_hd__a21bo_2 _22755_ (.A1(_06863_),
    .A2(_06864_),
    .B1_N(_06865_),
    .X(_06866_));
 sky130_fd_sc_hd__a22o_1 _22756_ (.A1(_06633_),
    .A2(_06743_),
    .B1(_06624_),
    .B2(_06744_),
    .X(_06867_));
 sky130_fd_sc_hd__o31a_2 _22757_ (.A1(_06626_),
    .A2(_06745_),
    .A3(_06631_),
    .B1(_06867_),
    .X(_06868_));
 sky130_fd_sc_hd__a2bb2oi_4 _22758_ (.A1_N(_06866_),
    .A2_N(_06868_),
    .B1(_06866_),
    .B2(_06868_),
    .Y(_02641_));
 sky130_fd_sc_hd__o22a_1 _22759_ (.A1(_06860_),
    .A2(_06861_),
    .B1(_06636_),
    .B2(_06862_),
    .X(_06869_));
 sky130_fd_sc_hd__o22a_1 _22760_ (.A1(_06732_),
    .A2(_06796_),
    .B1(_06751_),
    .B2(_06797_),
    .X(_06870_));
 sky130_fd_sc_hd__o22a_1 _22761_ (.A1(_06775_),
    .A2(_06776_),
    .B1(_06752_),
    .B2(_06777_),
    .X(_06871_));
 sky130_fd_sc_hd__or2_1 _22762_ (.A(_06870_),
    .B(_06871_),
    .X(_06872_));
 sky130_fd_sc_hd__a21bo_1 _22763_ (.A1(_06870_),
    .A2(_06871_),
    .B1_N(_06872_),
    .X(_06873_));
 sky130_fd_sc_hd__o22a_1 _22764_ (.A1(_06793_),
    .A2(_06794_),
    .B1(_06778_),
    .B2(_06795_),
    .X(_06874_));
 sky130_fd_sc_hd__a21oi_2 _22765_ (.A1(_06758_),
    .A2(_06759_),
    .B1(_06757_),
    .Y(_06875_));
 sky130_fd_sc_hd__buf_1 _22766_ (.A(_05816_),
    .X(_06876_));
 sky130_fd_sc_hd__clkbuf_2 _22767_ (.A(_06648_),
    .X(_06877_));
 sky130_fd_sc_hd__buf_2 _22768_ (.A(_06877_),
    .X(_06878_));
 sky130_fd_sc_hd__clkbuf_4 _22769_ (.A(_06878_),
    .X(_06879_));
 sky130_fd_sc_hd__buf_1 _22770_ (.A(_06761_),
    .X(_06880_));
 sky130_fd_sc_hd__clkbuf_2 _22771_ (.A(_06880_),
    .X(_06881_));
 sky130_fd_sc_hd__buf_1 _22772_ (.A(_06881_),
    .X(_06882_));
 sky130_fd_sc_hd__o22a_1 _22773_ (.A1(_06876_),
    .A2(_06879_),
    .B1(_05308_),
    .B2(_06882_),
    .X(_06883_));
 sky130_fd_sc_hd__clkbuf_2 _22774_ (.A(_13546_),
    .X(_06884_));
 sky130_fd_sc_hd__and4_1 _22775_ (.A(_13175_),
    .B(_13551_),
    .C(_13180_),
    .D(_06884_),
    .X(_06885_));
 sky130_fd_sc_hd__nor2_2 _22776_ (.A(_06883_),
    .B(_06885_),
    .Y(_06886_));
 sky130_fd_sc_hd__clkbuf_4 _22777_ (.A(_05828_),
    .X(_06887_));
 sky130_fd_sc_hd__nor2_4 _22778_ (.A(_06887_),
    .B(_06642_),
    .Y(_06888_));
 sky130_fd_sc_hd__a2bb2o_1 _22779_ (.A1_N(_06886_),
    .A2_N(_06888_),
    .B1(_06886_),
    .B2(_06888_),
    .X(_06889_));
 sky130_vsdinv _22780_ (.A(\pcpi_mul.rs1[23] ),
    .Y(_06890_));
 sky130_fd_sc_hd__clkbuf_2 _22781_ (.A(_06890_),
    .X(_06891_));
 sky130_fd_sc_hd__clkbuf_4 _22782_ (.A(_06891_),
    .X(_06892_));
 sky130_fd_sc_hd__or2_1 _22783_ (.A(_05311_),
    .B(_06892_),
    .X(_06893_));
 sky130_fd_sc_hd__clkbuf_2 _22784_ (.A(_06229_),
    .X(_06894_));
 sky130_fd_sc_hd__clkbuf_2 _22785_ (.A(_06230_),
    .X(_06895_));
 sky130_fd_sc_hd__o22a_1 _22786_ (.A1(_06894_),
    .A2(_06339_),
    .B1(_06895_),
    .B2(_06566_),
    .X(_06896_));
 sky130_fd_sc_hd__buf_1 _22787_ (.A(_06233_),
    .X(_06897_));
 sky130_fd_sc_hd__buf_1 _22788_ (.A(\pcpi_mul.rs1[18] ),
    .X(_06898_));
 sky130_fd_sc_hd__clkbuf_2 _22789_ (.A(_06898_),
    .X(_06899_));
 sky130_fd_sc_hd__buf_1 _22790_ (.A(_06235_),
    .X(_06900_));
 sky130_fd_sc_hd__clkbuf_2 _22791_ (.A(_13555_),
    .X(_06901_));
 sky130_fd_sc_hd__and4_1 _22792_ (.A(_06897_),
    .B(_06899_),
    .C(_06900_),
    .D(_06901_),
    .X(_06902_));
 sky130_fd_sc_hd__or2_1 _22793_ (.A(_06896_),
    .B(_06902_),
    .X(_06903_));
 sky130_fd_sc_hd__a2bb2o_1 _22794_ (.A1_N(_06893_),
    .A2_N(_06903_),
    .B1(_06893_),
    .B2(_06903_),
    .X(_06904_));
 sky130_fd_sc_hd__o21ba_1 _22795_ (.A1(_06764_),
    .A2(_06771_),
    .B1_N(_06770_),
    .X(_06905_));
 sky130_fd_sc_hd__a2bb2o_1 _22796_ (.A1_N(_06904_),
    .A2_N(_06905_),
    .B1(_06904_),
    .B2(_06905_),
    .X(_06906_));
 sky130_fd_sc_hd__a2bb2o_1 _22797_ (.A1_N(_06889_),
    .A2_N(_06906_),
    .B1(_06889_),
    .B2(_06906_),
    .X(_06907_));
 sky130_fd_sc_hd__o22a_1 _22798_ (.A1(_06772_),
    .A2(_06773_),
    .B1(_06760_),
    .B2(_06774_),
    .X(_06908_));
 sky130_fd_sc_hd__a2bb2o_1 _22799_ (.A1_N(_06907_),
    .A2_N(_06908_),
    .B1(_06907_),
    .B2(_06908_),
    .X(_06909_));
 sky130_fd_sc_hd__a2bb2o_1 _22800_ (.A1_N(_06875_),
    .A2_N(_06909_),
    .B1(_06875_),
    .B2(_06909_),
    .X(_06910_));
 sky130_fd_sc_hd__o22a_1 _22801_ (.A1(_06782_),
    .A2(_06789_),
    .B1(_06781_),
    .B2(_06790_),
    .X(_06911_));
 sky130_fd_sc_hd__o22a_1 _22802_ (.A1(_06835_),
    .A2(_06836_),
    .B1(_06828_),
    .B2(_06837_),
    .X(_06912_));
 sky130_fd_sc_hd__o21ba_1 _22803_ (.A1(_06784_),
    .A2(_06788_),
    .B1_N(_06787_),
    .X(_06913_));
 sky130_fd_sc_hd__o21ba_1 _22804_ (.A1(_06821_),
    .A2(_06827_),
    .B1_N(_06826_),
    .X(_06914_));
 sky130_fd_sc_hd__clkbuf_2 _22805_ (.A(_05423_),
    .X(_06915_));
 sky130_fd_sc_hd__clkbuf_2 _22806_ (.A(_06225_),
    .X(_06916_));
 sky130_fd_sc_hd__clkbuf_2 _22807_ (.A(_06916_),
    .X(_06917_));
 sky130_fd_sc_hd__or2_1 _22808_ (.A(_06915_),
    .B(_06917_),
    .X(_06918_));
 sky130_fd_sc_hd__clkbuf_2 _22809_ (.A(_05865_),
    .X(_06919_));
 sky130_fd_sc_hd__clkbuf_2 _22810_ (.A(_06252_),
    .X(_06920_));
 sky130_fd_sc_hd__clkbuf_2 _22811_ (.A(_06139_),
    .X(_06921_));
 sky130_fd_sc_hd__o22a_1 _22812_ (.A1(_06919_),
    .A2(_06131_),
    .B1(_06920_),
    .B2(_06921_),
    .X(_06922_));
 sky130_fd_sc_hd__clkbuf_2 _22813_ (.A(_06254_),
    .X(_06923_));
 sky130_fd_sc_hd__clkbuf_2 _22814_ (.A(_06255_),
    .X(_06924_));
 sky130_fd_sc_hd__buf_1 _22815_ (.A(_13566_),
    .X(_06925_));
 sky130_fd_sc_hd__and4_1 _22816_ (.A(_06923_),
    .B(_13570_),
    .C(_06924_),
    .D(_06925_),
    .X(_06926_));
 sky130_fd_sc_hd__or2_1 _22817_ (.A(_06922_),
    .B(_06926_),
    .X(_06927_));
 sky130_fd_sc_hd__a2bb2o_2 _22818_ (.A1_N(_06918_),
    .A2_N(_06927_),
    .B1(_06918_),
    .B2(_06927_),
    .X(_06928_));
 sky130_fd_sc_hd__a2bb2o_1 _22819_ (.A1_N(_06914_),
    .A2_N(_06928_),
    .B1(_06914_),
    .B2(_06928_),
    .X(_06929_));
 sky130_fd_sc_hd__a2bb2o_1 _22820_ (.A1_N(_06913_),
    .A2_N(_06929_),
    .B1(_06913_),
    .B2(_06929_),
    .X(_06930_));
 sky130_fd_sc_hd__a2bb2o_1 _22821_ (.A1_N(_06912_),
    .A2_N(_06930_),
    .B1(_06912_),
    .B2(_06930_),
    .X(_06931_));
 sky130_fd_sc_hd__a2bb2o_1 _22822_ (.A1_N(_06911_),
    .A2_N(_06931_),
    .B1(_06911_),
    .B2(_06931_),
    .X(_06932_));
 sky130_fd_sc_hd__o22a_1 _22823_ (.A1(_06780_),
    .A2(_06791_),
    .B1(_06779_),
    .B2(_06792_),
    .X(_06933_));
 sky130_fd_sc_hd__a2bb2o_1 _22824_ (.A1_N(_06932_),
    .A2_N(_06933_),
    .B1(_06932_),
    .B2(_06933_),
    .X(_06934_));
 sky130_fd_sc_hd__a2bb2o_1 _22825_ (.A1_N(_06910_),
    .A2_N(_06934_),
    .B1(_06910_),
    .B2(_06934_),
    .X(_06935_));
 sky130_fd_sc_hd__a2bb2o_1 _22826_ (.A1_N(_06852_),
    .A2_N(_06935_),
    .B1(_06852_),
    .B2(_06935_),
    .X(_06936_));
 sky130_fd_sc_hd__a2bb2o_1 _22827_ (.A1_N(_06874_),
    .A2_N(_06936_),
    .B1(_06874_),
    .B2(_06936_),
    .X(_06937_));
 sky130_fd_sc_hd__or2_1 _22828_ (.A(_06284_),
    .B(_05900_),
    .X(_06938_));
 sky130_fd_sc_hd__clkbuf_2 _22829_ (.A(_05684_),
    .X(_06939_));
 sky130_fd_sc_hd__o22a_1 _22830_ (.A1(_06810_),
    .A2(_06112_),
    .B1(_06394_),
    .B2(_06939_),
    .X(_06940_));
 sky130_fd_sc_hd__buf_2 _22831_ (.A(\pcpi_mul.rs2[19] ),
    .X(_06941_));
 sky130_fd_sc_hd__and4_1 _22832_ (.A(_13105_),
    .B(_06116_),
    .C(_06941_),
    .D(_13612_),
    .X(_06942_));
 sky130_fd_sc_hd__or2_1 _22833_ (.A(_06940_),
    .B(_06942_),
    .X(_06943_));
 sky130_fd_sc_hd__a2bb2o_1 _22834_ (.A1_N(_06938_),
    .A2_N(_06943_),
    .B1(_06938_),
    .B2(_06943_),
    .X(_06944_));
 sky130_fd_sc_hd__clkbuf_2 _22835_ (.A(_06686_),
    .X(_06945_));
 sky130_fd_sc_hd__or2_1 _22836_ (.A(_06945_),
    .B(_05908_),
    .X(_06946_));
 sky130_vsdinv _22837_ (.A(\pcpi_mul.rs2[23] ),
    .Y(_06947_));
 sky130_fd_sc_hd__clkbuf_2 _22838_ (.A(_06947_),
    .X(_06948_));
 sky130_fd_sc_hd__o22a_1 _22839_ (.A1(_06799_),
    .A2(_05380_),
    .B1(_06948_),
    .B2(_05363_),
    .X(_06949_));
 sky130_fd_sc_hd__buf_1 _22840_ (.A(\pcpi_mul.rs2[22] ),
    .X(_06950_));
 sky130_fd_sc_hd__and4_1 _22841_ (.A(_06950_),
    .B(_06695_),
    .C(\pcpi_mul.rs2[23] ),
    .D(_05917_),
    .X(_06951_));
 sky130_fd_sc_hd__or2_1 _22842_ (.A(_06949_),
    .B(_06951_),
    .X(_06952_));
 sky130_fd_sc_hd__a2bb2o_2 _22843_ (.A1_N(_06946_),
    .A2_N(_06952_),
    .B1(_06946_),
    .B2(_06952_),
    .X(_06953_));
 sky130_fd_sc_hd__a2bb2o_1 _22844_ (.A1_N(_06807_),
    .A2_N(_06953_),
    .B1(_06807_),
    .B2(_06953_),
    .X(_06954_));
 sky130_fd_sc_hd__a2bb2o_1 _22845_ (.A1_N(_06944_),
    .A2_N(_06954_),
    .B1(_06944_),
    .B2(_06954_),
    .X(_06955_));
 sky130_fd_sc_hd__or2_1 _22846_ (.A(_06815_),
    .B(_06955_),
    .X(_06956_));
 sky130_fd_sc_hd__a21bo_1 _22847_ (.A1(_06815_),
    .A2(_06955_),
    .B1_N(_06956_),
    .X(_06957_));
 sky130_fd_sc_hd__o22a_1 _22848_ (.A1(_06848_),
    .A2(_06849_),
    .B1(_06838_),
    .B2(_06850_),
    .X(_06958_));
 sky130_fd_sc_hd__or2_1 _22849_ (.A(_06820_),
    .B(_06130_),
    .X(_06959_));
 sky130_fd_sc_hd__clkbuf_2 _22850_ (.A(_05587_),
    .X(_06960_));
 sky130_fd_sc_hd__o22a_1 _22851_ (.A1(_06822_),
    .A2(_05927_),
    .B1(_06960_),
    .B2(_06231_),
    .X(_06961_));
 sky130_fd_sc_hd__clkbuf_2 _22852_ (.A(_06103_),
    .X(_06962_));
 sky130_fd_sc_hd__clkbuf_2 _22853_ (.A(_06104_),
    .X(_06963_));
 sky130_fd_sc_hd__and4_1 _22854_ (.A(_06962_),
    .B(_06602_),
    .C(_06963_),
    .D(_06603_),
    .X(_06964_));
 sky130_fd_sc_hd__or2_1 _22855_ (.A(_06961_),
    .B(_06964_),
    .X(_06965_));
 sky130_fd_sc_hd__a2bb2o_2 _22856_ (.A1_N(_06959_),
    .A2_N(_06965_),
    .B1(_06959_),
    .B2(_06965_),
    .X(_06966_));
 sky130_fd_sc_hd__buf_1 _22857_ (.A(_06108_),
    .X(_06967_));
 sky130_fd_sc_hd__or2_1 _22858_ (.A(_06967_),
    .B(_05725_),
    .X(_06968_));
 sky130_fd_sc_hd__clkbuf_2 _22859_ (.A(_06110_),
    .X(_06969_));
 sky130_fd_sc_hd__buf_1 _22860_ (.A(_06111_),
    .X(_06970_));
 sky130_fd_sc_hd__o22a_1 _22861_ (.A1(_06969_),
    .A2(_05843_),
    .B1(_06970_),
    .B2(_05830_),
    .X(_06971_));
 sky130_fd_sc_hd__buf_1 _22862_ (.A(_06114_),
    .X(_06972_));
 sky130_fd_sc_hd__buf_1 _22863_ (.A(_05914_),
    .X(_06973_));
 sky130_fd_sc_hd__buf_1 _22864_ (.A(_05655_),
    .X(_06974_));
 sky130_fd_sc_hd__and4_1 _22865_ (.A(_06972_),
    .B(_06526_),
    .C(_06973_),
    .D(_06974_),
    .X(_06975_));
 sky130_fd_sc_hd__or2_1 _22866_ (.A(_06971_),
    .B(_06975_),
    .X(_06976_));
 sky130_fd_sc_hd__a2bb2o_1 _22867_ (.A1_N(_06968_),
    .A2_N(_06976_),
    .B1(_06968_),
    .B2(_06976_),
    .X(_06977_));
 sky130_fd_sc_hd__o21ba_1 _22868_ (.A1(_06829_),
    .A2(_06834_),
    .B1_N(_06833_),
    .X(_06978_));
 sky130_fd_sc_hd__a2bb2o_1 _22869_ (.A1_N(_06977_),
    .A2_N(_06978_),
    .B1(_06977_),
    .B2(_06978_),
    .X(_06979_));
 sky130_fd_sc_hd__a2bb2o_1 _22870_ (.A1_N(_06966_),
    .A2_N(_06979_),
    .B1(_06966_),
    .B2(_06979_),
    .X(_06980_));
 sky130_fd_sc_hd__o21ba_1 _22871_ (.A1(_06841_),
    .A2(_06845_),
    .B1_N(_06844_),
    .X(_06981_));
 sky130_fd_sc_hd__o21ba_1 _22872_ (.A1(_06809_),
    .A2(_06813_),
    .B1_N(_06812_),
    .X(_06982_));
 sky130_fd_sc_hd__clkbuf_2 _22873_ (.A(_05840_),
    .X(_06983_));
 sky130_fd_sc_hd__or2_1 _22874_ (.A(_06095_),
    .B(_06983_),
    .X(_06984_));
 sky130_fd_sc_hd__o22a_1 _22875_ (.A1(_06842_),
    .A2(_06101_),
    .B1(_06088_),
    .B2(_05967_),
    .X(_06985_));
 sky130_fd_sc_hd__and4_1 _22876_ (.A(_06722_),
    .B(_13603_),
    .C(_06723_),
    .D(_05741_),
    .X(_06986_));
 sky130_fd_sc_hd__or2_1 _22877_ (.A(_06985_),
    .B(_06986_),
    .X(_06987_));
 sky130_fd_sc_hd__a2bb2o_1 _22878_ (.A1_N(_06984_),
    .A2_N(_06987_),
    .B1(_06984_),
    .B2(_06987_),
    .X(_06988_));
 sky130_fd_sc_hd__a2bb2o_1 _22879_ (.A1_N(_06982_),
    .A2_N(_06988_),
    .B1(_06982_),
    .B2(_06988_),
    .X(_06989_));
 sky130_fd_sc_hd__a2bb2o_1 _22880_ (.A1_N(_06981_),
    .A2_N(_06989_),
    .B1(_06981_),
    .B2(_06989_),
    .X(_06990_));
 sky130_fd_sc_hd__o22a_1 _22881_ (.A1(_06840_),
    .A2(_06846_),
    .B1(_06839_),
    .B2(_06847_),
    .X(_06991_));
 sky130_fd_sc_hd__a2bb2o_1 _22882_ (.A1_N(_06990_),
    .A2_N(_06991_),
    .B1(_06990_),
    .B2(_06991_),
    .X(_06992_));
 sky130_fd_sc_hd__a2bb2o_1 _22883_ (.A1_N(_06980_),
    .A2_N(_06992_),
    .B1(_06980_),
    .B2(_06992_),
    .X(_06993_));
 sky130_fd_sc_hd__a2bb2o_1 _22884_ (.A1_N(_06817_),
    .A2_N(_06993_),
    .B1(_06817_),
    .B2(_06993_),
    .X(_06994_));
 sky130_fd_sc_hd__a2bb2o_1 _22885_ (.A1_N(_06958_),
    .A2_N(_06994_),
    .B1(_06958_),
    .B2(_06994_),
    .X(_06995_));
 sky130_fd_sc_hd__or2_1 _22886_ (.A(_06957_),
    .B(_06995_),
    .X(_06996_));
 sky130_fd_sc_hd__a21bo_1 _22887_ (.A1(_06957_),
    .A2(_06995_),
    .B1_N(_06996_),
    .X(_06997_));
 sky130_fd_sc_hd__a2bb2o_1 _22888_ (.A1_N(_06854_),
    .A2_N(_06997_),
    .B1(_06854_),
    .B2(_06997_),
    .X(_06998_));
 sky130_fd_sc_hd__a2bb2o_1 _22889_ (.A1_N(_06937_),
    .A2_N(_06998_),
    .B1(_06937_),
    .B2(_06998_),
    .X(_06999_));
 sky130_fd_sc_hd__o22a_1 _22890_ (.A1(_06734_),
    .A2(_06855_),
    .B1(_06798_),
    .B2(_06856_),
    .X(_07000_));
 sky130_fd_sc_hd__a2bb2o_1 _22891_ (.A1_N(_06999_),
    .A2_N(_07000_),
    .B1(_06999_),
    .B2(_07000_),
    .X(_07001_));
 sky130_fd_sc_hd__a2bb2o_1 _22892_ (.A1_N(_06873_),
    .A2_N(_07001_),
    .B1(_06873_),
    .B2(_07001_),
    .X(_07002_));
 sky130_fd_sc_hd__o22a_1 _22893_ (.A1(_06857_),
    .A2(_06858_),
    .B1(_06750_),
    .B2(_06859_),
    .X(_07003_));
 sky130_fd_sc_hd__a2bb2o_1 _22894_ (.A1_N(_07002_),
    .A2_N(_07003_),
    .B1(_07002_),
    .B2(_07003_),
    .X(_07004_));
 sky130_fd_sc_hd__a2bb2o_2 _22895_ (.A1_N(_06749_),
    .A2_N(_07004_),
    .B1(_06749_),
    .B2(_07004_),
    .X(_07005_));
 sky130_fd_sc_hd__and2_1 _22896_ (.A(_06869_),
    .B(_07005_),
    .X(_07006_));
 sky130_fd_sc_hd__or2_1 _22897_ (.A(_06869_),
    .B(_07005_),
    .X(_07007_));
 sky130_fd_sc_hd__or2b_1 _22898_ (.A(_07006_),
    .B_N(_07007_),
    .X(_07008_));
 sky130_fd_sc_hd__o21ai_1 _22899_ (.A1(_06866_),
    .A2(_06868_),
    .B1(_06865_),
    .Y(_07009_));
 sky130_fd_sc_hd__a2bb2o_2 _22900_ (.A1_N(_07008_),
    .A2_N(_07009_),
    .B1(_07008_),
    .B2(_07009_),
    .X(_02642_));
 sky130_fd_sc_hd__o22a_1 _22901_ (.A1(_06852_),
    .A2(_06935_),
    .B1(_06874_),
    .B2(_06936_),
    .X(_07010_));
 sky130_fd_sc_hd__o22a_1 _22902_ (.A1(_06907_),
    .A2(_06908_),
    .B1(_06875_),
    .B2(_06909_),
    .X(_07011_));
 sky130_fd_sc_hd__or2_1 _22903_ (.A(_07010_),
    .B(_07011_),
    .X(_07012_));
 sky130_fd_sc_hd__a21bo_1 _22904_ (.A1(_07010_),
    .A2(_07011_),
    .B1_N(_07012_),
    .X(_07013_));
 sky130_fd_sc_hd__o22a_1 _22905_ (.A1(_06932_),
    .A2(_06933_),
    .B1(_06910_),
    .B2(_06934_),
    .X(_07014_));
 sky130_fd_sc_hd__o22a_1 _22906_ (.A1(_06817_),
    .A2(_06993_),
    .B1(_06958_),
    .B2(_06994_),
    .X(_07015_));
 sky130_fd_sc_hd__a21oi_4 _22907_ (.A1(_06886_),
    .A2(_06888_),
    .B1(_06885_),
    .Y(_07016_));
 sky130_fd_sc_hd__buf_1 _22908_ (.A(_05307_),
    .X(_07017_));
 sky130_fd_sc_hd__buf_1 _22909_ (.A(_06890_),
    .X(_07018_));
 sky130_fd_sc_hd__buf_2 _22910_ (.A(_07018_),
    .X(_07019_));
 sky130_fd_sc_hd__buf_1 _22911_ (.A(_07019_),
    .X(_07020_));
 sky130_fd_sc_hd__o22a_1 _22912_ (.A1(_06876_),
    .A2(_06882_),
    .B1(_07017_),
    .B2(_07020_),
    .X(_07021_));
 sky130_fd_sc_hd__buf_1 _22913_ (.A(_13174_),
    .X(_07022_));
 sky130_fd_sc_hd__buf_1 _22914_ (.A(_13179_),
    .X(_07023_));
 sky130_fd_sc_hd__buf_1 _22915_ (.A(_13542_),
    .X(_07024_));
 sky130_fd_sc_hd__and4_2 _22916_ (.A(_07022_),
    .B(_06884_),
    .C(_07023_),
    .D(_07024_),
    .X(_07025_));
 sky130_fd_sc_hd__nor2_2 _22917_ (.A(_07021_),
    .B(_07025_),
    .Y(_07026_));
 sky130_fd_sc_hd__buf_2 _22918_ (.A(_05828_),
    .X(_07027_));
 sky130_fd_sc_hd__nor2_4 _22919_ (.A(_07027_),
    .B(_06879_),
    .Y(_07028_));
 sky130_fd_sc_hd__a2bb2o_1 _22920_ (.A1_N(_07026_),
    .A2_N(_07028_),
    .B1(_07026_),
    .B2(_07028_),
    .X(_07029_));
 sky130_fd_sc_hd__buf_1 _22921_ (.A(_05142_),
    .X(_07030_));
 sky130_vsdinv _22922_ (.A(\pcpi_mul.rs1[24] ),
    .Y(_07031_));
 sky130_fd_sc_hd__buf_1 _22923_ (.A(_07031_),
    .X(_07032_));
 sky130_fd_sc_hd__clkbuf_2 _22924_ (.A(_07032_),
    .X(_07033_));
 sky130_fd_sc_hd__clkbuf_4 _22925_ (.A(_07033_),
    .X(_07034_));
 sky130_fd_sc_hd__or2_1 _22926_ (.A(_07030_),
    .B(_07034_),
    .X(_07035_));
 sky130_fd_sc_hd__clkbuf_2 _22927_ (.A(_06450_),
    .X(_07036_));
 sky130_fd_sc_hd__clkbuf_2 _22928_ (.A(_06640_),
    .X(_07037_));
 sky130_fd_sc_hd__o22a_1 _22929_ (.A1(_06894_),
    .A2(_07036_),
    .B1(_06895_),
    .B2(_07037_),
    .X(_07038_));
 sky130_fd_sc_hd__buf_1 _22930_ (.A(\pcpi_mul.rs1[20] ),
    .X(_07039_));
 sky130_fd_sc_hd__clkbuf_2 _22931_ (.A(_07039_),
    .X(_07040_));
 sky130_fd_sc_hd__and4_1 _22932_ (.A(_06897_),
    .B(_06901_),
    .C(_06900_),
    .D(_07040_),
    .X(_07041_));
 sky130_fd_sc_hd__or2_1 _22933_ (.A(_07038_),
    .B(_07041_),
    .X(_07042_));
 sky130_fd_sc_hd__a2bb2o_1 _22934_ (.A1_N(_07035_),
    .A2_N(_07042_),
    .B1(_07035_),
    .B2(_07042_),
    .X(_07043_));
 sky130_fd_sc_hd__o21ba_1 _22935_ (.A1(_06893_),
    .A2(_06903_),
    .B1_N(_06902_),
    .X(_07044_));
 sky130_fd_sc_hd__a2bb2o_1 _22936_ (.A1_N(_07043_),
    .A2_N(_07044_),
    .B1(_07043_),
    .B2(_07044_),
    .X(_07045_));
 sky130_fd_sc_hd__a2bb2o_1 _22937_ (.A1_N(_07029_),
    .A2_N(_07045_),
    .B1(_07029_),
    .B2(_07045_),
    .X(_07046_));
 sky130_fd_sc_hd__o22a_1 _22938_ (.A1(_06904_),
    .A2(_06905_),
    .B1(_06889_),
    .B2(_06906_),
    .X(_07047_));
 sky130_fd_sc_hd__a2bb2o_1 _22939_ (.A1_N(_07046_),
    .A2_N(_07047_),
    .B1(_07046_),
    .B2(_07047_),
    .X(_07048_));
 sky130_fd_sc_hd__a2bb2o_2 _22940_ (.A1_N(_07016_),
    .A2_N(_07048_),
    .B1(_07016_),
    .B2(_07048_),
    .X(_07049_));
 sky130_fd_sc_hd__o22a_1 _22941_ (.A1(_06914_),
    .A2(_06928_),
    .B1(_06913_),
    .B2(_06929_),
    .X(_07050_));
 sky130_fd_sc_hd__o22a_1 _22942_ (.A1(_06977_),
    .A2(_06978_),
    .B1(_06966_),
    .B2(_06979_),
    .X(_07051_));
 sky130_fd_sc_hd__o21ba_1 _22943_ (.A1(_06918_),
    .A2(_06927_),
    .B1_N(_06926_),
    .X(_07052_));
 sky130_fd_sc_hd__o21ba_1 _22944_ (.A1(_06959_),
    .A2(_06965_),
    .B1_N(_06964_),
    .X(_07053_));
 sky130_fd_sc_hd__or2_1 _22945_ (.A(_05424_),
    .B(_06438_),
    .X(_07054_));
 sky130_fd_sc_hd__clkbuf_2 _22946_ (.A(_05865_),
    .X(_07055_));
 sky130_fd_sc_hd__o22a_1 _22947_ (.A1(_07055_),
    .A2(_06326_),
    .B1(_06920_),
    .B2(_06916_),
    .X(_07056_));
 sky130_fd_sc_hd__buf_1 _22948_ (.A(_06254_),
    .X(_07057_));
 sky130_fd_sc_hd__buf_1 _22949_ (.A(_06255_),
    .X(_07058_));
 sky130_fd_sc_hd__clkbuf_2 _22950_ (.A(_13563_),
    .X(_07059_));
 sky130_fd_sc_hd__and4_1 _22951_ (.A(_07057_),
    .B(_06925_),
    .C(_07058_),
    .D(_07059_),
    .X(_07060_));
 sky130_fd_sc_hd__or2_1 _22952_ (.A(_07056_),
    .B(_07060_),
    .X(_07061_));
 sky130_fd_sc_hd__a2bb2o_1 _22953_ (.A1_N(_07054_),
    .A2_N(_07061_),
    .B1(_07054_),
    .B2(_07061_),
    .X(_07062_));
 sky130_fd_sc_hd__a2bb2o_1 _22954_ (.A1_N(_07053_),
    .A2_N(_07062_),
    .B1(_07053_),
    .B2(_07062_),
    .X(_07063_));
 sky130_fd_sc_hd__a2bb2o_1 _22955_ (.A1_N(_07052_),
    .A2_N(_07063_),
    .B1(_07052_),
    .B2(_07063_),
    .X(_07064_));
 sky130_fd_sc_hd__a2bb2o_1 _22956_ (.A1_N(_07051_),
    .A2_N(_07064_),
    .B1(_07051_),
    .B2(_07064_),
    .X(_07065_));
 sky130_fd_sc_hd__a2bb2o_1 _22957_ (.A1_N(_07050_),
    .A2_N(_07065_),
    .B1(_07050_),
    .B2(_07065_),
    .X(_07066_));
 sky130_fd_sc_hd__o22a_1 _22958_ (.A1(_06912_),
    .A2(_06930_),
    .B1(_06911_),
    .B2(_06931_),
    .X(_07067_));
 sky130_fd_sc_hd__a2bb2o_1 _22959_ (.A1_N(_07066_),
    .A2_N(_07067_),
    .B1(_07066_),
    .B2(_07067_),
    .X(_07068_));
 sky130_fd_sc_hd__a2bb2o_1 _22960_ (.A1_N(_07049_),
    .A2_N(_07068_),
    .B1(_07049_),
    .B2(_07068_),
    .X(_07069_));
 sky130_fd_sc_hd__a2bb2o_1 _22961_ (.A1_N(_07015_),
    .A2_N(_07069_),
    .B1(_07015_),
    .B2(_07069_),
    .X(_07070_));
 sky130_fd_sc_hd__a2bb2o_1 _22962_ (.A1_N(_07014_),
    .A2_N(_07070_),
    .B1(_07014_),
    .B2(_07070_),
    .X(_07071_));
 sky130_vsdinv _22963_ (.A(\pcpi_mul.rs2[24] ),
    .Y(_07072_));
 sky130_fd_sc_hd__buf_1 _22964_ (.A(_07072_),
    .X(_07073_));
 sky130_fd_sc_hd__clkbuf_4 _22965_ (.A(_07073_),
    .X(_07074_));
 sky130_fd_sc_hd__clkbuf_2 _22966_ (.A(_07074_),
    .X(_07075_));
 sky130_fd_sc_hd__clkbuf_4 _22967_ (.A(_07075_),
    .X(_07076_));
 sky130_fd_sc_hd__or2_1 _22968_ (.A(_07076_),
    .B(_05590_),
    .X(_07077_));
 sky130_fd_sc_hd__buf_1 _22969_ (.A(_06396_),
    .X(_07078_));
 sky130_fd_sc_hd__clkbuf_2 _22970_ (.A(_05868_),
    .X(_07079_));
 sky130_fd_sc_hd__or2_1 _22971_ (.A(_07078_),
    .B(_07079_),
    .X(_07080_));
 sky130_fd_sc_hd__buf_2 _22972_ (.A(_06514_),
    .X(_07081_));
 sky130_fd_sc_hd__buf_2 _22973_ (.A(_05366_),
    .X(_07082_));
 sky130_fd_sc_hd__o22a_1 _22974_ (.A1(_07081_),
    .A2(_07082_),
    .B1(_06389_),
    .B2(_06201_),
    .X(_07083_));
 sky130_fd_sc_hd__buf_1 _22975_ (.A(_06694_),
    .X(_07084_));
 sky130_fd_sc_hd__clkbuf_2 _22976_ (.A(_05758_),
    .X(_07085_));
 sky130_fd_sc_hd__clkbuf_2 _22977_ (.A(_06311_),
    .X(_07086_));
 sky130_fd_sc_hd__and4_1 _22978_ (.A(_07084_),
    .B(_07085_),
    .C(_13111_),
    .D(_07086_),
    .X(_07087_));
 sky130_fd_sc_hd__or2_1 _22979_ (.A(_07083_),
    .B(_07087_),
    .X(_07088_));
 sky130_fd_sc_hd__a2bb2o_1 _22980_ (.A1_N(_07080_),
    .A2_N(_07088_),
    .B1(_07080_),
    .B2(_07088_),
    .X(_07089_));
 sky130_fd_sc_hd__or2_1 _22981_ (.A(_06945_),
    .B(_06011_),
    .X(_07090_));
 sky130_fd_sc_hd__o22a_1 _22982_ (.A1(_06947_),
    .A2(_05380_),
    .B1(_06800_),
    .B2(_05645_),
    .X(_07091_));
 sky130_fd_sc_hd__buf_1 _22983_ (.A(\pcpi_mul.rs2[23] ),
    .X(_07092_));
 sky130_fd_sc_hd__and4_1 _22984_ (.A(_07092_),
    .B(_06695_),
    .C(\pcpi_mul.rs2[22] ),
    .D(_05346_),
    .X(_07093_));
 sky130_fd_sc_hd__or2_1 _22985_ (.A(_07091_),
    .B(_07093_),
    .X(_07094_));
 sky130_fd_sc_hd__a2bb2o_1 _22986_ (.A1_N(_07090_),
    .A2_N(_07094_),
    .B1(_07090_),
    .B2(_07094_),
    .X(_07095_));
 sky130_fd_sc_hd__o21ba_1 _22987_ (.A1(_06946_),
    .A2(_06952_),
    .B1_N(_06951_),
    .X(_07096_));
 sky130_fd_sc_hd__a2bb2o_1 _22988_ (.A1_N(_07095_),
    .A2_N(_07096_),
    .B1(_07095_),
    .B2(_07096_),
    .X(_07097_));
 sky130_fd_sc_hd__a2bb2o_1 _22989_ (.A1_N(_07089_),
    .A2_N(_07097_),
    .B1(_07089_),
    .B2(_07097_),
    .X(_07098_));
 sky130_fd_sc_hd__o22a_1 _22990_ (.A1(_06807_),
    .A2(_06953_),
    .B1(_06944_),
    .B2(_06954_),
    .X(_07099_));
 sky130_fd_sc_hd__or2_1 _22991_ (.A(_07098_),
    .B(_07099_),
    .X(_07100_));
 sky130_fd_sc_hd__a21bo_1 _22992_ (.A1(_07098_),
    .A2(_07099_),
    .B1_N(_07100_),
    .X(_07101_));
 sky130_fd_sc_hd__or2_1 _22993_ (.A(_07077_),
    .B(_07101_),
    .X(_07102_));
 sky130_fd_sc_hd__a21bo_1 _22994_ (.A1(_07077_),
    .A2(_07101_),
    .B1_N(_07102_),
    .X(_07103_));
 sky130_fd_sc_hd__o22a_1 _22995_ (.A1(_06990_),
    .A2(_06991_),
    .B1(_06980_),
    .B2(_06992_),
    .X(_07104_));
 sky130_fd_sc_hd__buf_1 _22996_ (.A(_05536_),
    .X(_07105_));
 sky130_fd_sc_hd__or2_1 _22997_ (.A(_07105_),
    .B(_06669_),
    .X(_07106_));
 sky130_fd_sc_hd__clkbuf_2 _22998_ (.A(_05714_),
    .X(_07107_));
 sky130_fd_sc_hd__buf_2 _22999_ (.A(_05802_),
    .X(_07108_));
 sky130_fd_sc_hd__o22a_1 _23000_ (.A1(_07107_),
    .A2(_06478_),
    .B1(_07108_),
    .B2(_06129_),
    .X(_07109_));
 sky130_fd_sc_hd__and4_1 _23001_ (.A(_06962_),
    .B(_06236_),
    .C(_06963_),
    .D(_06673_),
    .X(_07110_));
 sky130_fd_sc_hd__or2_1 _23002_ (.A(_07109_),
    .B(_07110_),
    .X(_07111_));
 sky130_fd_sc_hd__a2bb2o_1 _23003_ (.A1_N(_07106_),
    .A2_N(_07111_),
    .B1(_07106_),
    .B2(_07111_),
    .X(_07112_));
 sky130_fd_sc_hd__or2_1 _23004_ (.A(_06967_),
    .B(_06702_),
    .X(_07113_));
 sky130_fd_sc_hd__o22a_1 _23005_ (.A1(_06969_),
    .A2(_06042_),
    .B1(_06970_),
    .B2(_06482_),
    .X(_07114_));
 sky130_fd_sc_hd__clkbuf_2 _23006_ (.A(_06114_),
    .X(_07115_));
 sky130_fd_sc_hd__clkbuf_2 _23007_ (.A(_05914_),
    .X(_07116_));
 sky130_fd_sc_hd__buf_1 _23008_ (.A(_06143_),
    .X(_07117_));
 sky130_fd_sc_hd__and4_1 _23009_ (.A(_07115_),
    .B(_06974_),
    .C(_07116_),
    .D(_07117_),
    .X(_07118_));
 sky130_fd_sc_hd__or2_1 _23010_ (.A(_07114_),
    .B(_07118_),
    .X(_07119_));
 sky130_fd_sc_hd__a2bb2o_1 _23011_ (.A1_N(_07113_),
    .A2_N(_07119_),
    .B1(_07113_),
    .B2(_07119_),
    .X(_07120_));
 sky130_fd_sc_hd__o21ba_1 _23012_ (.A1(_06968_),
    .A2(_06976_),
    .B1_N(_06975_),
    .X(_07121_));
 sky130_fd_sc_hd__a2bb2o_1 _23013_ (.A1_N(_07120_),
    .A2_N(_07121_),
    .B1(_07120_),
    .B2(_07121_),
    .X(_07122_));
 sky130_fd_sc_hd__a2bb2o_1 _23014_ (.A1_N(_07112_),
    .A2_N(_07122_),
    .B1(_07112_),
    .B2(_07122_),
    .X(_07123_));
 sky130_fd_sc_hd__o21ba_1 _23015_ (.A1(_06984_),
    .A2(_06987_),
    .B1_N(_06986_),
    .X(_07124_));
 sky130_fd_sc_hd__o21ba_1 _23016_ (.A1(_06938_),
    .A2(_06943_),
    .B1_N(_06942_),
    .X(_07125_));
 sky130_fd_sc_hd__clkbuf_2 _23017_ (.A(_06251_),
    .X(_07126_));
 sky130_fd_sc_hd__or2_1 _23018_ (.A(_05998_),
    .B(_07126_),
    .X(_07127_));
 sky130_fd_sc_hd__buf_2 _23019_ (.A(_06546_),
    .X(_07128_));
 sky130_fd_sc_hd__o22a_1 _23020_ (.A1(_07128_),
    .A2(_05967_),
    .B1(_06088_),
    .B2(_05662_),
    .X(_07129_));
 sky130_fd_sc_hd__and4_1 _23021_ (.A(_13117_),
    .B(_13598_),
    .C(_13121_),
    .D(_13594_),
    .X(_07130_));
 sky130_fd_sc_hd__or2_1 _23022_ (.A(_07129_),
    .B(_07130_),
    .X(_07131_));
 sky130_fd_sc_hd__a2bb2o_1 _23023_ (.A1_N(_07127_),
    .A2_N(_07131_),
    .B1(_07127_),
    .B2(_07131_),
    .X(_07132_));
 sky130_fd_sc_hd__a2bb2o_1 _23024_ (.A1_N(_07125_),
    .A2_N(_07132_),
    .B1(_07125_),
    .B2(_07132_),
    .X(_07133_));
 sky130_fd_sc_hd__a2bb2o_1 _23025_ (.A1_N(_07124_),
    .A2_N(_07133_),
    .B1(_07124_),
    .B2(_07133_),
    .X(_07134_));
 sky130_fd_sc_hd__o22a_1 _23026_ (.A1(_06982_),
    .A2(_06988_),
    .B1(_06981_),
    .B2(_06989_),
    .X(_07135_));
 sky130_fd_sc_hd__a2bb2o_1 _23027_ (.A1_N(_07134_),
    .A2_N(_07135_),
    .B1(_07134_),
    .B2(_07135_),
    .X(_07136_));
 sky130_fd_sc_hd__a2bb2o_1 _23028_ (.A1_N(_07123_),
    .A2_N(_07136_),
    .B1(_07123_),
    .B2(_07136_),
    .X(_07137_));
 sky130_fd_sc_hd__a2bb2o_1 _23029_ (.A1_N(_06956_),
    .A2_N(_07137_),
    .B1(_06956_),
    .B2(_07137_),
    .X(_07138_));
 sky130_fd_sc_hd__a2bb2o_1 _23030_ (.A1_N(_07104_),
    .A2_N(_07138_),
    .B1(_07104_),
    .B2(_07138_),
    .X(_07139_));
 sky130_fd_sc_hd__or2_1 _23031_ (.A(_07103_),
    .B(_07139_),
    .X(_07140_));
 sky130_fd_sc_hd__a21bo_1 _23032_ (.A1(_07103_),
    .A2(_07139_),
    .B1_N(_07140_),
    .X(_07141_));
 sky130_fd_sc_hd__a2bb2o_1 _23033_ (.A1_N(_06996_),
    .A2_N(_07141_),
    .B1(_06996_),
    .B2(_07141_),
    .X(_07142_));
 sky130_fd_sc_hd__a2bb2o_1 _23034_ (.A1_N(_07071_),
    .A2_N(_07142_),
    .B1(_07071_),
    .B2(_07142_),
    .X(_07143_));
 sky130_fd_sc_hd__o22a_1 _23035_ (.A1(_06854_),
    .A2(_06997_),
    .B1(_06937_),
    .B2(_06998_),
    .X(_07144_));
 sky130_fd_sc_hd__a2bb2o_1 _23036_ (.A1_N(_07143_),
    .A2_N(_07144_),
    .B1(_07143_),
    .B2(_07144_),
    .X(_07145_));
 sky130_fd_sc_hd__a2bb2o_1 _23037_ (.A1_N(_07013_),
    .A2_N(_07145_),
    .B1(_07013_),
    .B2(_07145_),
    .X(_07146_));
 sky130_fd_sc_hd__o22a_1 _23038_ (.A1(_06999_),
    .A2(_07000_),
    .B1(_06873_),
    .B2(_07001_),
    .X(_07147_));
 sky130_fd_sc_hd__a2bb2o_1 _23039_ (.A1_N(_07146_),
    .A2_N(_07147_),
    .B1(_07146_),
    .B2(_07147_),
    .X(_07148_));
 sky130_fd_sc_hd__a2bb2o_1 _23040_ (.A1_N(_06872_),
    .A2_N(_07148_),
    .B1(_06872_),
    .B2(_07148_),
    .X(_07149_));
 sky130_fd_sc_hd__o22a_1 _23041_ (.A1(_07002_),
    .A2(_07003_),
    .B1(_06749_),
    .B2(_07004_),
    .X(_07150_));
 sky130_fd_sc_hd__or2_1 _23042_ (.A(_07149_),
    .B(_07150_),
    .X(_07151_));
 sky130_fd_sc_hd__a21bo_1 _23043_ (.A1(_07149_),
    .A2(_07150_),
    .B1_N(_07151_),
    .X(_07152_));
 sky130_fd_sc_hd__buf_1 _23044_ (.A(_07152_),
    .X(_07153_));
 sky130_fd_sc_hd__or2_1 _23045_ (.A(_06866_),
    .B(_07008_),
    .X(_07154_));
 sky130_fd_sc_hd__or3_1 _23046_ (.A(_06625_),
    .B(_06745_),
    .C(_07154_),
    .X(_07155_));
 sky130_fd_sc_hd__or3_4 _23047_ (.A(_06628_),
    .B(_07155_),
    .C(_06081_),
    .X(_07156_));
 sky130_fd_sc_hd__o21a_1 _23048_ (.A1(_06865_),
    .A2(_07006_),
    .B1(_07007_),
    .X(_07157_));
 sky130_fd_sc_hd__o221a_4 _23049_ (.A1(_06867_),
    .A2(_07154_),
    .B1(_06629_),
    .B2(_07155_),
    .C1(_07157_),
    .X(_07158_));
 sky130_fd_sc_hd__nand2_1 _23050_ (.A(_07156_),
    .B(_07158_),
    .Y(_07159_));
 sky130_vsdinv _23051_ (.A(_07159_),
    .Y(_07160_));
 sky130_vsdinv _23052_ (.A(_07153_),
    .Y(_07161_));
 sky130_fd_sc_hd__o22a_1 _23053_ (.A1(_07153_),
    .A2(_07160_),
    .B1(_07161_),
    .B2(_07159_),
    .X(_02643_));
 sky130_fd_sc_hd__o22a_1 _23054_ (.A1(_07146_),
    .A2(_07147_),
    .B1(_06872_),
    .B2(_07148_),
    .X(_07162_));
 sky130_fd_sc_hd__o22a_1 _23055_ (.A1(_07015_),
    .A2(_07069_),
    .B1(_07014_),
    .B2(_07070_),
    .X(_07163_));
 sky130_fd_sc_hd__o22a_1 _23056_ (.A1(_07046_),
    .A2(_07047_),
    .B1(_07016_),
    .B2(_07048_),
    .X(_07164_));
 sky130_fd_sc_hd__or2_1 _23057_ (.A(_07163_),
    .B(_07164_),
    .X(_07165_));
 sky130_fd_sc_hd__a21bo_1 _23058_ (.A1(_07163_),
    .A2(_07164_),
    .B1_N(_07165_),
    .X(_07166_));
 sky130_fd_sc_hd__o22a_1 _23059_ (.A1(_07066_),
    .A2(_07067_),
    .B1(_07049_),
    .B2(_07068_),
    .X(_07167_));
 sky130_fd_sc_hd__o22a_1 _23060_ (.A1(_06956_),
    .A2(_07137_),
    .B1(_07104_),
    .B2(_07138_),
    .X(_07168_));
 sky130_fd_sc_hd__a21oi_4 _23061_ (.A1(_07026_),
    .A2(_07028_),
    .B1(_07025_),
    .Y(_07169_));
 sky130_fd_sc_hd__buf_1 _23062_ (.A(_07018_),
    .X(_07170_));
 sky130_fd_sc_hd__clkbuf_4 _23063_ (.A(_07170_),
    .X(_07171_));
 sky130_fd_sc_hd__clkbuf_2 _23064_ (.A(_07032_),
    .X(_07172_));
 sky130_fd_sc_hd__clkbuf_2 _23065_ (.A(_07172_),
    .X(_07173_));
 sky130_fd_sc_hd__o22a_1 _23066_ (.A1(_06433_),
    .A2(_07171_),
    .B1(_07017_),
    .B2(_07173_),
    .X(_07174_));
 sky130_fd_sc_hd__buf_1 _23067_ (.A(_13539_),
    .X(_07175_));
 sky130_fd_sc_hd__and4_2 _23068_ (.A(_07022_),
    .B(_07024_),
    .C(_07023_),
    .D(_07175_),
    .X(_07176_));
 sky130_fd_sc_hd__nor2_2 _23069_ (.A(_07174_),
    .B(_07176_),
    .Y(_07177_));
 sky130_fd_sc_hd__clkbuf_4 _23070_ (.A(_06763_),
    .X(_07178_));
 sky130_fd_sc_hd__nor2_4 _23071_ (.A(_07027_),
    .B(_07178_),
    .Y(_07179_));
 sky130_fd_sc_hd__a2bb2o_1 _23072_ (.A1_N(_07177_),
    .A2_N(_07179_),
    .B1(_07177_),
    .B2(_07179_),
    .X(_07180_));
 sky130_fd_sc_hd__buf_1 _23073_ (.A(_05737_),
    .X(_07181_));
 sky130_fd_sc_hd__buf_1 _23074_ (.A(_07181_),
    .X(_07182_));
 sky130_fd_sc_hd__buf_1 _23075_ (.A(_05739_),
    .X(_07183_));
 sky130_fd_sc_hd__buf_1 _23076_ (.A(_07183_),
    .X(_07184_));
 sky130_fd_sc_hd__o22a_1 _23077_ (.A1(_07182_),
    .A2(_06641_),
    .B1(_07184_),
    .B2(_06878_),
    .X(_07185_));
 sky130_fd_sc_hd__buf_1 _23078_ (.A(_06233_),
    .X(_07186_));
 sky130_fd_sc_hd__clkbuf_2 _23079_ (.A(_07039_),
    .X(_07187_));
 sky130_fd_sc_hd__buf_1 _23080_ (.A(_07187_),
    .X(_07188_));
 sky130_fd_sc_hd__buf_1 _23081_ (.A(_06235_),
    .X(_07189_));
 sky130_fd_sc_hd__buf_1 _23082_ (.A(\pcpi_mul.rs1[21] ),
    .X(_07190_));
 sky130_fd_sc_hd__clkbuf_2 _23083_ (.A(_07190_),
    .X(_07191_));
 sky130_fd_sc_hd__buf_1 _23084_ (.A(_07191_),
    .X(_07192_));
 sky130_fd_sc_hd__and4_1 _23085_ (.A(_07186_),
    .B(_07188_),
    .C(_07189_),
    .D(_07192_),
    .X(_07193_));
 sky130_fd_sc_hd__nor2_2 _23086_ (.A(_07185_),
    .B(_07193_),
    .Y(_07194_));
 sky130_vsdinv _23087_ (.A(\pcpi_mul.rs1[25] ),
    .Y(_07195_));
 sky130_fd_sc_hd__buf_1 _23088_ (.A(_07195_),
    .X(_07196_));
 sky130_fd_sc_hd__clkbuf_2 _23089_ (.A(_07196_),
    .X(_07197_));
 sky130_fd_sc_hd__clkbuf_2 _23090_ (.A(_07197_),
    .X(_07198_));
 sky130_fd_sc_hd__nor2_2 _23091_ (.A(_05311_),
    .B(_07198_),
    .Y(_07199_));
 sky130_fd_sc_hd__a2bb2o_1 _23092_ (.A1_N(_07194_),
    .A2_N(_07199_),
    .B1(_07194_),
    .B2(_07199_),
    .X(_07200_));
 sky130_fd_sc_hd__o21ba_1 _23093_ (.A1(_07035_),
    .A2(_07042_),
    .B1_N(_07041_),
    .X(_07201_));
 sky130_fd_sc_hd__a2bb2o_1 _23094_ (.A1_N(_07200_),
    .A2_N(_07201_),
    .B1(_07200_),
    .B2(_07201_),
    .X(_07202_));
 sky130_fd_sc_hd__a2bb2o_1 _23095_ (.A1_N(_07180_),
    .A2_N(_07202_),
    .B1(_07180_),
    .B2(_07202_),
    .X(_07203_));
 sky130_fd_sc_hd__o22a_1 _23096_ (.A1(_07043_),
    .A2(_07044_),
    .B1(_07029_),
    .B2(_07045_),
    .X(_07204_));
 sky130_fd_sc_hd__a2bb2o_1 _23097_ (.A1_N(_07203_),
    .A2_N(_07204_),
    .B1(_07203_),
    .B2(_07204_),
    .X(_07205_));
 sky130_fd_sc_hd__a2bb2o_1 _23098_ (.A1_N(_07169_),
    .A2_N(_07205_),
    .B1(_07169_),
    .B2(_07205_),
    .X(_07206_));
 sky130_fd_sc_hd__o22a_1 _23099_ (.A1(_07053_),
    .A2(_07062_),
    .B1(_07052_),
    .B2(_07063_),
    .X(_07207_));
 sky130_fd_sc_hd__o22a_1 _23100_ (.A1(_07120_),
    .A2(_07121_),
    .B1(_07112_),
    .B2(_07122_),
    .X(_07208_));
 sky130_fd_sc_hd__o21ba_1 _23101_ (.A1(_07054_),
    .A2(_07061_),
    .B1_N(_07060_),
    .X(_07209_));
 sky130_fd_sc_hd__o21ba_1 _23102_ (.A1(_07106_),
    .A2(_07111_),
    .B1_N(_07110_),
    .X(_07210_));
 sky130_fd_sc_hd__or2_1 _23103_ (.A(_05424_),
    .B(_06566_),
    .X(_07211_));
 sky130_fd_sc_hd__buf_1 _23104_ (.A(_13559_),
    .X(_07212_));
 sky130_fd_sc_hd__and4_1 _23105_ (.A(_07057_),
    .B(_07059_),
    .C(_07058_),
    .D(_07212_),
    .X(_07213_));
 sky130_fd_sc_hd__clkbuf_2 _23106_ (.A(_06252_),
    .X(_07214_));
 sky130_fd_sc_hd__o22a_1 _23107_ (.A1(_06481_),
    .A2(_06226_),
    .B1(_07214_),
    .B2(_06437_),
    .X(_07215_));
 sky130_fd_sc_hd__or2_1 _23108_ (.A(_07213_),
    .B(_07215_),
    .X(_07216_));
 sky130_fd_sc_hd__a2bb2o_1 _23109_ (.A1_N(_07211_),
    .A2_N(_07216_),
    .B1(_07211_),
    .B2(_07216_),
    .X(_07217_));
 sky130_fd_sc_hd__a2bb2o_1 _23110_ (.A1_N(_07210_),
    .A2_N(_07217_),
    .B1(_07210_),
    .B2(_07217_),
    .X(_07218_));
 sky130_fd_sc_hd__a2bb2o_1 _23111_ (.A1_N(_07209_),
    .A2_N(_07218_),
    .B1(_07209_),
    .B2(_07218_),
    .X(_07219_));
 sky130_fd_sc_hd__a2bb2o_1 _23112_ (.A1_N(_07208_),
    .A2_N(_07219_),
    .B1(_07208_),
    .B2(_07219_),
    .X(_07220_));
 sky130_fd_sc_hd__a2bb2o_1 _23113_ (.A1_N(_07207_),
    .A2_N(_07220_),
    .B1(_07207_),
    .B2(_07220_),
    .X(_07221_));
 sky130_fd_sc_hd__o22a_1 _23114_ (.A1(_07051_),
    .A2(_07064_),
    .B1(_07050_),
    .B2(_07065_),
    .X(_07222_));
 sky130_fd_sc_hd__a2bb2o_1 _23115_ (.A1_N(_07221_),
    .A2_N(_07222_),
    .B1(_07221_),
    .B2(_07222_),
    .X(_07223_));
 sky130_fd_sc_hd__a2bb2o_1 _23116_ (.A1_N(_07206_),
    .A2_N(_07223_),
    .B1(_07206_),
    .B2(_07223_),
    .X(_07224_));
 sky130_fd_sc_hd__a2bb2o_1 _23117_ (.A1_N(_07168_),
    .A2_N(_07224_),
    .B1(_07168_),
    .B2(_07224_),
    .X(_07225_));
 sky130_fd_sc_hd__a2bb2o_1 _23118_ (.A1_N(_07167_),
    .A2_N(_07225_),
    .B1(_07167_),
    .B2(_07225_),
    .X(_07226_));
 sky130_fd_sc_hd__o22a_1 _23119_ (.A1(_07134_),
    .A2(_07135_),
    .B1(_07123_),
    .B2(_07136_),
    .X(_07227_));
 sky130_fd_sc_hd__or2_1 _23120_ (.A(_06519_),
    .B(_06783_),
    .X(_07228_));
 sky130_fd_sc_hd__and4_1 _23121_ (.A(_06824_),
    .B(_06673_),
    .C(_06825_),
    .D(_06786_),
    .X(_07229_));
 sky130_fd_sc_hd__o22a_1 _23122_ (.A1(_06522_),
    .A2(_05943_),
    .B1(_06523_),
    .B2(_06668_),
    .X(_07230_));
 sky130_fd_sc_hd__or2_1 _23123_ (.A(_07229_),
    .B(_07230_),
    .X(_07231_));
 sky130_fd_sc_hd__a2bb2o_1 _23124_ (.A1_N(_07228_),
    .A2_N(_07231_),
    .B1(_07228_),
    .B2(_07231_),
    .X(_07232_));
 sky130_fd_sc_hd__or2_1 _23125_ (.A(_05791_),
    .B(_05837_),
    .X(_07233_));
 sky130_fd_sc_hd__buf_1 _23126_ (.A(_06535_),
    .X(_07234_));
 sky130_fd_sc_hd__buf_1 _23127_ (.A(_06536_),
    .X(_07235_));
 sky130_fd_sc_hd__and4_1 _23128_ (.A(_07234_),
    .B(_07117_),
    .C(_07235_),
    .D(_06145_),
    .X(_07236_));
 sky130_fd_sc_hd__clkbuf_2 _23129_ (.A(_05912_),
    .X(_07237_));
 sky130_fd_sc_hd__buf_2 _23130_ (.A(_06111_),
    .X(_07238_));
 sky130_fd_sc_hd__o22a_1 _23131_ (.A1(_07237_),
    .A2(_06043_),
    .B1(_07238_),
    .B2(_05927_),
    .X(_07239_));
 sky130_fd_sc_hd__or2_1 _23132_ (.A(_07236_),
    .B(_07239_),
    .X(_07240_));
 sky130_fd_sc_hd__a2bb2o_1 _23133_ (.A1_N(_07233_),
    .A2_N(_07240_),
    .B1(_07233_),
    .B2(_07240_),
    .X(_07241_));
 sky130_fd_sc_hd__o21ba_1 _23134_ (.A1(_07113_),
    .A2(_07119_),
    .B1_N(_07118_),
    .X(_07242_));
 sky130_fd_sc_hd__a2bb2o_1 _23135_ (.A1_N(_07241_),
    .A2_N(_07242_),
    .B1(_07241_),
    .B2(_07242_),
    .X(_07243_));
 sky130_fd_sc_hd__a2bb2o_1 _23136_ (.A1_N(_07232_),
    .A2_N(_07243_),
    .B1(_07232_),
    .B2(_07243_),
    .X(_07244_));
 sky130_fd_sc_hd__o21ba_1 _23137_ (.A1(_07127_),
    .A2(_07131_),
    .B1_N(_07130_),
    .X(_07245_));
 sky130_fd_sc_hd__o21ba_1 _23138_ (.A1(_07080_),
    .A2(_07088_),
    .B1_N(_07087_),
    .X(_07246_));
 sky130_fd_sc_hd__or2_1 _23139_ (.A(_06096_),
    .B(_05831_),
    .X(_07247_));
 sky130_fd_sc_hd__buf_1 _23140_ (.A(_13117_),
    .X(_07248_));
 sky130_fd_sc_hd__buf_1 _23141_ (.A(_13594_),
    .X(_07249_));
 sky130_fd_sc_hd__buf_1 _23142_ (.A(_13121_),
    .X(_07250_));
 sky130_fd_sc_hd__buf_1 _23143_ (.A(_05654_),
    .X(_07251_));
 sky130_fd_sc_hd__and4_1 _23144_ (.A(_07248_),
    .B(_07249_),
    .C(_07250_),
    .D(_07251_),
    .X(_07252_));
 sky130_fd_sc_hd__clkbuf_4 _23145_ (.A(_06842_),
    .X(_07253_));
 sky130_fd_sc_hd__buf_1 _23146_ (.A(_06092_),
    .X(_07254_));
 sky130_fd_sc_hd__clkbuf_2 _23147_ (.A(_05729_),
    .X(_07255_));
 sky130_fd_sc_hd__o22a_1 _23148_ (.A1(_07253_),
    .A2(_05963_),
    .B1(_07254_),
    .B2(_07255_),
    .X(_07256_));
 sky130_fd_sc_hd__or2_1 _23149_ (.A(_07252_),
    .B(_07256_),
    .X(_07257_));
 sky130_fd_sc_hd__a2bb2o_1 _23150_ (.A1_N(_07247_),
    .A2_N(_07257_),
    .B1(_07247_),
    .B2(_07257_),
    .X(_07258_));
 sky130_fd_sc_hd__a2bb2o_1 _23151_ (.A1_N(_07246_),
    .A2_N(_07258_),
    .B1(_07246_),
    .B2(_07258_),
    .X(_07259_));
 sky130_fd_sc_hd__a2bb2o_2 _23152_ (.A1_N(_07245_),
    .A2_N(_07259_),
    .B1(_07245_),
    .B2(_07259_),
    .X(_07260_));
 sky130_fd_sc_hd__o22a_1 _23153_ (.A1(_07125_),
    .A2(_07132_),
    .B1(_07124_),
    .B2(_07133_),
    .X(_07261_));
 sky130_fd_sc_hd__a2bb2o_1 _23154_ (.A1_N(_07260_),
    .A2_N(_07261_),
    .B1(_07260_),
    .B2(_07261_),
    .X(_07262_));
 sky130_fd_sc_hd__a2bb2o_1 _23155_ (.A1_N(_07244_),
    .A2_N(_07262_),
    .B1(_07244_),
    .B2(_07262_),
    .X(_07263_));
 sky130_fd_sc_hd__a2bb2o_1 _23156_ (.A1_N(_07100_),
    .A2_N(_07263_),
    .B1(_07100_),
    .B2(_07263_),
    .X(_07264_));
 sky130_fd_sc_hd__a2bb2o_1 _23157_ (.A1_N(_07227_),
    .A2_N(_07264_),
    .B1(_07227_),
    .B2(_07264_),
    .X(_07265_));
 sky130_vsdinv _23158_ (.A(\pcpi_mul.rs2[25] ),
    .Y(_07266_));
 sky130_fd_sc_hd__clkbuf_2 _23159_ (.A(_07266_),
    .X(_07267_));
 sky130_fd_sc_hd__clkbuf_2 _23160_ (.A(_07267_),
    .X(_07268_));
 sky130_fd_sc_hd__buf_2 _23161_ (.A(_07268_),
    .X(_07269_));
 sky130_fd_sc_hd__clkbuf_4 _23162_ (.A(_07269_),
    .X(_07270_));
 sky130_fd_sc_hd__o22a_1 _23163_ (.A1(_07270_),
    .A2(_05153_),
    .B1(_07076_),
    .B2(_05300_),
    .X(_07271_));
 sky130_fd_sc_hd__clkbuf_4 _23164_ (.A(_07267_),
    .X(_07272_));
 sky130_fd_sc_hd__clkbuf_2 _23165_ (.A(_07073_),
    .X(_07273_));
 sky130_fd_sc_hd__or4_4 _23166_ (.A(_07272_),
    .B(_05150_),
    .C(_07273_),
    .D(_05298_),
    .X(_07274_));
 sky130_fd_sc_hd__or2b_1 _23167_ (.A(_07271_),
    .B_N(_07274_),
    .X(_07275_));
 sky130_fd_sc_hd__o22a_1 _23168_ (.A1(_07095_),
    .A2(_07096_),
    .B1(_07089_),
    .B2(_07097_),
    .X(_07276_));
 sky130_fd_sc_hd__buf_1 _23169_ (.A(_05738_),
    .X(_07277_));
 sky130_fd_sc_hd__clkbuf_2 _23170_ (.A(_07277_),
    .X(_07278_));
 sky130_fd_sc_hd__or2_1 _23171_ (.A(_07078_),
    .B(_07278_),
    .X(_07279_));
 sky130_fd_sc_hd__and4_1 _23172_ (.A(_07084_),
    .B(_07086_),
    .C(_13111_),
    .D(_05872_),
    .X(_07280_));
 sky130_fd_sc_hd__buf_1 _23173_ (.A(_06810_),
    .X(_07281_));
 sky130_fd_sc_hd__buf_1 _23174_ (.A(_06394_),
    .X(_07282_));
 sky130_fd_sc_hd__o22a_1 _23175_ (.A1(_07281_),
    .A2(_05866_),
    .B1(_07282_),
    .B2(_06308_),
    .X(_07283_));
 sky130_fd_sc_hd__or2_1 _23176_ (.A(_07280_),
    .B(_07283_),
    .X(_07284_));
 sky130_fd_sc_hd__a2bb2o_1 _23177_ (.A1_N(_07279_),
    .A2_N(_07284_),
    .B1(_07279_),
    .B2(_07284_),
    .X(_07285_));
 sky130_fd_sc_hd__or2_1 _23178_ (.A(_06945_),
    .B(_07082_),
    .X(_07286_));
 sky130_fd_sc_hd__and4_1 _23179_ (.A(_07092_),
    .B(_05806_),
    .C(_06950_),
    .D(_06204_),
    .X(_07287_));
 sky130_fd_sc_hd__o22a_1 _23180_ (.A1(_06947_),
    .A2(_05343_),
    .B1(_06800_),
    .B2(_05803_),
    .X(_07288_));
 sky130_fd_sc_hd__or2_1 _23181_ (.A(_07287_),
    .B(_07288_),
    .X(_07289_));
 sky130_fd_sc_hd__a2bb2o_1 _23182_ (.A1_N(_07286_),
    .A2_N(_07289_),
    .B1(_07286_),
    .B2(_07289_),
    .X(_07290_));
 sky130_fd_sc_hd__o21ba_1 _23183_ (.A1(_07090_),
    .A2(_07094_),
    .B1_N(_07093_),
    .X(_07291_));
 sky130_fd_sc_hd__a2bb2o_1 _23184_ (.A1_N(_07290_),
    .A2_N(_07291_),
    .B1(_07290_),
    .B2(_07291_),
    .X(_07292_));
 sky130_fd_sc_hd__a2bb2o_1 _23185_ (.A1_N(_07285_),
    .A2_N(_07292_),
    .B1(_07285_),
    .B2(_07292_),
    .X(_07293_));
 sky130_fd_sc_hd__or2_1 _23186_ (.A(_07276_),
    .B(_07293_),
    .X(_07294_));
 sky130_fd_sc_hd__a21bo_1 _23187_ (.A1(_07276_),
    .A2(_07293_),
    .B1_N(_07294_),
    .X(_07295_));
 sky130_fd_sc_hd__or2_1 _23188_ (.A(_07275_),
    .B(_07295_),
    .X(_07296_));
 sky130_fd_sc_hd__a21bo_1 _23189_ (.A1(_07275_),
    .A2(_07295_),
    .B1_N(_07296_),
    .X(_07297_));
 sky130_fd_sc_hd__a2bb2o_1 _23190_ (.A1_N(_07102_),
    .A2_N(_07297_),
    .B1(_07102_),
    .B2(_07297_),
    .X(_07298_));
 sky130_fd_sc_hd__a2bb2o_1 _23191_ (.A1_N(_07265_),
    .A2_N(_07298_),
    .B1(_07265_),
    .B2(_07298_),
    .X(_07299_));
 sky130_fd_sc_hd__a2bb2o_1 _23192_ (.A1_N(_07140_),
    .A2_N(_07299_),
    .B1(_07140_),
    .B2(_07299_),
    .X(_07300_));
 sky130_fd_sc_hd__a2bb2o_1 _23193_ (.A1_N(_07226_),
    .A2_N(_07300_),
    .B1(_07226_),
    .B2(_07300_),
    .X(_07301_));
 sky130_fd_sc_hd__o22a_1 _23194_ (.A1(_06996_),
    .A2(_07141_),
    .B1(_07071_),
    .B2(_07142_),
    .X(_07302_));
 sky130_fd_sc_hd__a2bb2o_1 _23195_ (.A1_N(_07301_),
    .A2_N(_07302_),
    .B1(_07301_),
    .B2(_07302_),
    .X(_07303_));
 sky130_fd_sc_hd__a2bb2o_1 _23196_ (.A1_N(_07166_),
    .A2_N(_07303_),
    .B1(_07166_),
    .B2(_07303_),
    .X(_07304_));
 sky130_fd_sc_hd__o22a_1 _23197_ (.A1(_07143_),
    .A2(_07144_),
    .B1(_07013_),
    .B2(_07145_),
    .X(_07305_));
 sky130_fd_sc_hd__a2bb2o_1 _23198_ (.A1_N(_07304_),
    .A2_N(_07305_),
    .B1(_07304_),
    .B2(_07305_),
    .X(_07306_));
 sky130_fd_sc_hd__a2bb2o_1 _23199_ (.A1_N(_07012_),
    .A2_N(_07306_),
    .B1(_07012_),
    .B2(_07306_),
    .X(_07307_));
 sky130_fd_sc_hd__or2_1 _23200_ (.A(_07162_),
    .B(_07307_),
    .X(_07308_));
 sky130_fd_sc_hd__a21bo_1 _23201_ (.A1(_07162_),
    .A2(_07307_),
    .B1_N(_07308_),
    .X(_07309_));
 sky130_fd_sc_hd__o21ai_1 _23202_ (.A1(_07153_),
    .A2(_07160_),
    .B1(_07151_),
    .Y(_07310_));
 sky130_fd_sc_hd__a2bb2o_1 _23203_ (.A1_N(_07309_),
    .A2_N(_07310_),
    .B1(_07309_),
    .B2(_07310_),
    .X(_02644_));
 sky130_fd_sc_hd__o22a_1 _23204_ (.A1(_07168_),
    .A2(_07224_),
    .B1(_07167_),
    .B2(_07225_),
    .X(_07311_));
 sky130_fd_sc_hd__o22a_1 _23205_ (.A1(_07203_),
    .A2(_07204_),
    .B1(_07169_),
    .B2(_07205_),
    .X(_07312_));
 sky130_fd_sc_hd__or2_1 _23206_ (.A(_07311_),
    .B(_07312_),
    .X(_07313_));
 sky130_fd_sc_hd__a21bo_1 _23207_ (.A1(_07311_),
    .A2(_07312_),
    .B1_N(_07313_),
    .X(_07314_));
 sky130_fd_sc_hd__o22a_1 _23208_ (.A1(_07221_),
    .A2(_07222_),
    .B1(_07206_),
    .B2(_07223_),
    .X(_07315_));
 sky130_fd_sc_hd__o22a_1 _23209_ (.A1(_07100_),
    .A2(_07263_),
    .B1(_07227_),
    .B2(_07264_),
    .X(_07316_));
 sky130_fd_sc_hd__a21oi_4 _23210_ (.A1(_07177_),
    .A2(_07179_),
    .B1(_07176_),
    .Y(_07317_));
 sky130_fd_sc_hd__o22a_1 _23211_ (.A1(_06433_),
    .A2(_07173_),
    .B1(_07017_),
    .B2(_07198_),
    .X(_07318_));
 sky130_fd_sc_hd__and4_1 _23212_ (.A(_07022_),
    .B(_07175_),
    .C(_07023_),
    .D(_13536_),
    .X(_07319_));
 sky130_fd_sc_hd__nor2_2 _23213_ (.A(_07318_),
    .B(_07319_),
    .Y(_07320_));
 sky130_fd_sc_hd__clkbuf_4 _23214_ (.A(_07019_),
    .X(_07321_));
 sky130_fd_sc_hd__nor2_2 _23215_ (.A(_07027_),
    .B(_07321_),
    .Y(_07322_));
 sky130_fd_sc_hd__a2bb2o_1 _23216_ (.A1_N(_07320_),
    .A2_N(_07322_),
    .B1(_07320_),
    .B2(_07322_),
    .X(_07323_));
 sky130_vsdinv _23217_ (.A(\pcpi_mul.rs1[26] ),
    .Y(_07324_));
 sky130_fd_sc_hd__buf_1 _23218_ (.A(_07324_),
    .X(_07325_));
 sky130_fd_sc_hd__clkbuf_2 _23219_ (.A(_07325_),
    .X(_07326_));
 sky130_fd_sc_hd__buf_2 _23220_ (.A(_07326_),
    .X(_07327_));
 sky130_fd_sc_hd__or2_1 _23221_ (.A(_06448_),
    .B(_07327_),
    .X(_07328_));
 sky130_fd_sc_hd__buf_1 _23222_ (.A(_07190_),
    .X(_07329_));
 sky130_fd_sc_hd__buf_1 _23223_ (.A(_13545_),
    .X(_07330_));
 sky130_fd_sc_hd__and4_1 _23224_ (.A(_06897_),
    .B(_07329_),
    .C(_06900_),
    .D(_07330_),
    .X(_07331_));
 sky130_fd_sc_hd__clkbuf_2 _23225_ (.A(_06880_),
    .X(_07332_));
 sky130_fd_sc_hd__o22a_1 _23226_ (.A1(_06454_),
    .A2(_06650_),
    .B1(_06455_),
    .B2(_07332_),
    .X(_07333_));
 sky130_fd_sc_hd__or2_1 _23227_ (.A(_07331_),
    .B(_07333_),
    .X(_07334_));
 sky130_fd_sc_hd__a2bb2o_1 _23228_ (.A1_N(_07328_),
    .A2_N(_07334_),
    .B1(_07328_),
    .B2(_07334_),
    .X(_07335_));
 sky130_fd_sc_hd__a21oi_2 _23229_ (.A1(_07194_),
    .A2(_07199_),
    .B1(_07193_),
    .Y(_07336_));
 sky130_fd_sc_hd__a2bb2o_1 _23230_ (.A1_N(_07335_),
    .A2_N(_07336_),
    .B1(_07335_),
    .B2(_07336_),
    .X(_07337_));
 sky130_fd_sc_hd__a2bb2o_1 _23231_ (.A1_N(_07323_),
    .A2_N(_07337_),
    .B1(_07323_),
    .B2(_07337_),
    .X(_07338_));
 sky130_fd_sc_hd__o22a_1 _23232_ (.A1(_07200_),
    .A2(_07201_),
    .B1(_07180_),
    .B2(_07202_),
    .X(_07339_));
 sky130_fd_sc_hd__a2bb2o_1 _23233_ (.A1_N(_07338_),
    .A2_N(_07339_),
    .B1(_07338_),
    .B2(_07339_),
    .X(_07340_));
 sky130_fd_sc_hd__a2bb2o_1 _23234_ (.A1_N(_07317_),
    .A2_N(_07340_),
    .B1(_07317_),
    .B2(_07340_),
    .X(_07341_));
 sky130_fd_sc_hd__o22a_1 _23235_ (.A1(_07210_),
    .A2(_07217_),
    .B1(_07209_),
    .B2(_07218_),
    .X(_07342_));
 sky130_fd_sc_hd__o22a_1 _23236_ (.A1(_07241_),
    .A2(_07242_),
    .B1(_07232_),
    .B2(_07243_),
    .X(_07343_));
 sky130_fd_sc_hd__o21ba_1 _23237_ (.A1(_07211_),
    .A2(_07216_),
    .B1_N(_07213_),
    .X(_07344_));
 sky130_fd_sc_hd__o21ba_1 _23238_ (.A1(_07228_),
    .A2(_07231_),
    .B1_N(_07229_),
    .X(_07345_));
 sky130_fd_sc_hd__or2_1 _23239_ (.A(_06477_),
    .B(_07037_),
    .X(_07346_));
 sky130_fd_sc_hd__and4_1 _23240_ (.A(_07057_),
    .B(_07212_),
    .C(_07058_),
    .D(_13555_),
    .X(_07347_));
 sky130_fd_sc_hd__clkbuf_2 _23241_ (.A(_06449_),
    .X(_07348_));
 sky130_fd_sc_hd__o22a_1 _23242_ (.A1(_06481_),
    .A2(_06338_),
    .B1(_06483_),
    .B2(_07348_),
    .X(_07349_));
 sky130_fd_sc_hd__or2_1 _23243_ (.A(_07347_),
    .B(_07349_),
    .X(_07350_));
 sky130_fd_sc_hd__a2bb2o_1 _23244_ (.A1_N(_07346_),
    .A2_N(_07350_),
    .B1(_07346_),
    .B2(_07350_),
    .X(_07351_));
 sky130_fd_sc_hd__a2bb2o_1 _23245_ (.A1_N(_07345_),
    .A2_N(_07351_),
    .B1(_07345_),
    .B2(_07351_),
    .X(_07352_));
 sky130_fd_sc_hd__a2bb2o_1 _23246_ (.A1_N(_07344_),
    .A2_N(_07352_),
    .B1(_07344_),
    .B2(_07352_),
    .X(_07353_));
 sky130_fd_sc_hd__a2bb2o_1 _23247_ (.A1_N(_07343_),
    .A2_N(_07353_),
    .B1(_07343_),
    .B2(_07353_),
    .X(_07354_));
 sky130_fd_sc_hd__a2bb2o_1 _23248_ (.A1_N(_07342_),
    .A2_N(_07354_),
    .B1(_07342_),
    .B2(_07354_),
    .X(_07355_));
 sky130_fd_sc_hd__o22a_1 _23249_ (.A1(_07208_),
    .A2(_07219_),
    .B1(_07207_),
    .B2(_07220_),
    .X(_07356_));
 sky130_fd_sc_hd__a2bb2o_1 _23250_ (.A1_N(_07355_),
    .A2_N(_07356_),
    .B1(_07355_),
    .B2(_07356_),
    .X(_07357_));
 sky130_fd_sc_hd__a2bb2o_1 _23251_ (.A1_N(_07341_),
    .A2_N(_07357_),
    .B1(_07341_),
    .B2(_07357_),
    .X(_07358_));
 sky130_fd_sc_hd__a2bb2o_1 _23252_ (.A1_N(_07316_),
    .A2_N(_07358_),
    .B1(_07316_),
    .B2(_07358_),
    .X(_07359_));
 sky130_fd_sc_hd__a2bb2o_1 _23253_ (.A1_N(_07315_),
    .A2_N(_07359_),
    .B1(_07315_),
    .B2(_07359_),
    .X(_07360_));
 sky130_fd_sc_hd__o22a_1 _23254_ (.A1(_07260_),
    .A2(_07261_),
    .B1(_07244_),
    .B2(_07262_),
    .X(_07361_));
 sky130_fd_sc_hd__or2_1 _23255_ (.A(_06820_),
    .B(_06917_),
    .X(_07362_));
 sky130_fd_sc_hd__clkbuf_2 _23256_ (.A(_06103_),
    .X(_07363_));
 sky130_fd_sc_hd__clkbuf_2 _23257_ (.A(_06104_),
    .X(_07364_));
 sky130_fd_sc_hd__and4_1 _23258_ (.A(_07363_),
    .B(_06786_),
    .C(_07364_),
    .D(_06925_),
    .X(_07365_));
 sky130_fd_sc_hd__o22a_1 _23259_ (.A1(_07107_),
    .A2(_06456_),
    .B1(_06960_),
    .B2(_06326_),
    .X(_07366_));
 sky130_fd_sc_hd__or2_1 _23260_ (.A(_07365_),
    .B(_07366_),
    .X(_07367_));
 sky130_fd_sc_hd__a2bb2o_1 _23261_ (.A1_N(_07362_),
    .A2_N(_07367_),
    .B1(_07362_),
    .B2(_07367_),
    .X(_07368_));
 sky130_fd_sc_hd__clkbuf_2 _23262_ (.A(_06108_),
    .X(_07369_));
 sky130_fd_sc_hd__or2_1 _23263_ (.A(_07369_),
    .B(_06599_),
    .X(_07370_));
 sky130_fd_sc_hd__buf_1 _23264_ (.A(\pcpi_mul.rs1[13] ),
    .X(_07371_));
 sky130_fd_sc_hd__and4_1 _23265_ (.A(_07234_),
    .B(_06234_),
    .C(_07235_),
    .D(_07371_),
    .X(_07372_));
 sky130_fd_sc_hd__o22a_1 _23266_ (.A1(_07237_),
    .A2(_05819_),
    .B1(_06970_),
    .B2(_06231_),
    .X(_07373_));
 sky130_fd_sc_hd__or2_1 _23267_ (.A(_07372_),
    .B(_07373_),
    .X(_07374_));
 sky130_fd_sc_hd__a2bb2o_1 _23268_ (.A1_N(_07370_),
    .A2_N(_07374_),
    .B1(_07370_),
    .B2(_07374_),
    .X(_07375_));
 sky130_fd_sc_hd__o21ba_1 _23269_ (.A1(_07233_),
    .A2(_07240_),
    .B1_N(_07236_),
    .X(_07376_));
 sky130_fd_sc_hd__a2bb2o_1 _23270_ (.A1_N(_07375_),
    .A2_N(_07376_),
    .B1(_07375_),
    .B2(_07376_),
    .X(_07377_));
 sky130_fd_sc_hd__a2bb2o_1 _23271_ (.A1_N(_07368_),
    .A2_N(_07377_),
    .B1(_07368_),
    .B2(_07377_),
    .X(_07378_));
 sky130_fd_sc_hd__o21ba_1 _23272_ (.A1(_07247_),
    .A2(_07257_),
    .B1_N(_07252_),
    .X(_07379_));
 sky130_fd_sc_hd__o21ba_1 _23273_ (.A1(_07279_),
    .A2(_07284_),
    .B1_N(_07280_),
    .X(_07380_));
 sky130_fd_sc_hd__or2_1 _23274_ (.A(_05999_),
    .B(_06520_),
    .X(_07381_));
 sky130_fd_sc_hd__and4_1 _23275_ (.A(_13118_),
    .B(_07251_),
    .C(_13122_),
    .D(_06974_),
    .X(_07382_));
 sky130_fd_sc_hd__clkbuf_2 _23276_ (.A(_06842_),
    .X(_07383_));
 sky130_fd_sc_hd__o22a_1 _23277_ (.A1(_07383_),
    .A2(_05730_),
    .B1(_06089_),
    .B2(_05830_),
    .X(_07384_));
 sky130_fd_sc_hd__or2_1 _23278_ (.A(_07382_),
    .B(_07384_),
    .X(_07385_));
 sky130_fd_sc_hd__a2bb2o_1 _23279_ (.A1_N(_07381_),
    .A2_N(_07385_),
    .B1(_07381_),
    .B2(_07385_),
    .X(_07386_));
 sky130_fd_sc_hd__a2bb2o_1 _23280_ (.A1_N(_07380_),
    .A2_N(_07386_),
    .B1(_07380_),
    .B2(_07386_),
    .X(_07387_));
 sky130_fd_sc_hd__a2bb2o_1 _23281_ (.A1_N(_07379_),
    .A2_N(_07387_),
    .B1(_07379_),
    .B2(_07387_),
    .X(_07388_));
 sky130_fd_sc_hd__o22a_1 _23282_ (.A1(_07246_),
    .A2(_07258_),
    .B1(_07245_),
    .B2(_07259_),
    .X(_07389_));
 sky130_fd_sc_hd__a2bb2o_1 _23283_ (.A1_N(_07388_),
    .A2_N(_07389_),
    .B1(_07388_),
    .B2(_07389_),
    .X(_07390_));
 sky130_fd_sc_hd__a2bb2o_1 _23284_ (.A1_N(_07378_),
    .A2_N(_07390_),
    .B1(_07378_),
    .B2(_07390_),
    .X(_07391_));
 sky130_fd_sc_hd__a2bb2o_1 _23285_ (.A1_N(_07294_),
    .A2_N(_07391_),
    .B1(_07294_),
    .B2(_07391_),
    .X(_07392_));
 sky130_fd_sc_hd__a2bb2o_1 _23286_ (.A1_N(_07361_),
    .A2_N(_07392_),
    .B1(_07361_),
    .B2(_07392_),
    .X(_07393_));
 sky130_fd_sc_hd__or2_1 _23287_ (.A(_07072_),
    .B(_05908_),
    .X(_07394_));
 sky130_fd_sc_hd__clkbuf_2 _23288_ (.A(\pcpi_mul.rs2[25] ),
    .X(_07395_));
 sky130_fd_sc_hd__and4_1 _23289_ (.A(_07395_),
    .B(_13623_),
    .C(\pcpi_mul.rs2[26] ),
    .D(_05917_),
    .X(_07396_));
 sky130_vsdinv _23290_ (.A(\pcpi_mul.rs2[26] ),
    .Y(_07397_));
 sky130_fd_sc_hd__o22a_1 _23291_ (.A1(_07266_),
    .A2(_05317_),
    .B1(_07397_),
    .B2(_05363_),
    .X(_07398_));
 sky130_fd_sc_hd__or2_1 _23292_ (.A(_07396_),
    .B(_07398_),
    .X(_07399_));
 sky130_fd_sc_hd__a2bb2o_1 _23293_ (.A1_N(_07394_),
    .A2_N(_07399_),
    .B1(_07394_),
    .B2(_07399_),
    .X(_07400_));
 sky130_fd_sc_hd__or2_2 _23294_ (.A(_07274_),
    .B(_07400_),
    .X(_07401_));
 sky130_fd_sc_hd__a21bo_1 _23295_ (.A1(_07274_),
    .A2(_07400_),
    .B1_N(_07401_),
    .X(_07402_));
 sky130_fd_sc_hd__clkbuf_2 _23296_ (.A(_05963_),
    .X(_07403_));
 sky130_fd_sc_hd__or2_1 _23297_ (.A(_07078_),
    .B(_07403_),
    .X(_07404_));
 sky130_fd_sc_hd__clkbuf_2 _23298_ (.A(_05969_),
    .X(_07405_));
 sky130_fd_sc_hd__buf_1 _23299_ (.A(_06941_),
    .X(_07406_));
 sky130_fd_sc_hd__and4_1 _23300_ (.A(_07084_),
    .B(_07405_),
    .C(_07406_),
    .D(_06303_),
    .X(_07407_));
 sky130_fd_sc_hd__o22a_1 _23301_ (.A1(_07281_),
    .A2(_06308_),
    .B1(_07282_),
    .B2(_07277_),
    .X(_07408_));
 sky130_fd_sc_hd__or2_1 _23302_ (.A(_07407_),
    .B(_07408_),
    .X(_07409_));
 sky130_fd_sc_hd__a2bb2o_1 _23303_ (.A1_N(_07404_),
    .A2_N(_07409_),
    .B1(_07404_),
    .B2(_07409_),
    .X(_07410_));
 sky130_fd_sc_hd__or2_1 _23304_ (.A(_06945_),
    .B(_06201_),
    .X(_07411_));
 sky130_fd_sc_hd__and4_1 _23305_ (.A(_07092_),
    .B(_05808_),
    .C(_06950_),
    .D(_13612_),
    .X(_07412_));
 sky130_fd_sc_hd__o22a_1 _23306_ (.A1(_06948_),
    .A2(_05902_),
    .B1(_06800_),
    .B2(_05798_),
    .X(_07413_));
 sky130_fd_sc_hd__or2_1 _23307_ (.A(_07412_),
    .B(_07413_),
    .X(_07414_));
 sky130_fd_sc_hd__a2bb2o_1 _23308_ (.A1_N(_07411_),
    .A2_N(_07414_),
    .B1(_07411_),
    .B2(_07414_),
    .X(_07415_));
 sky130_fd_sc_hd__o21ba_1 _23309_ (.A1(_07286_),
    .A2(_07289_),
    .B1_N(_07287_),
    .X(_07416_));
 sky130_fd_sc_hd__a2bb2o_1 _23310_ (.A1_N(_07415_),
    .A2_N(_07416_),
    .B1(_07415_),
    .B2(_07416_),
    .X(_07417_));
 sky130_fd_sc_hd__a2bb2o_1 _23311_ (.A1_N(_07410_),
    .A2_N(_07417_),
    .B1(_07410_),
    .B2(_07417_),
    .X(_07418_));
 sky130_fd_sc_hd__o22a_1 _23312_ (.A1(_07290_),
    .A2(_07291_),
    .B1(_07285_),
    .B2(_07292_),
    .X(_07419_));
 sky130_fd_sc_hd__or2_1 _23313_ (.A(_07418_),
    .B(_07419_),
    .X(_07420_));
 sky130_fd_sc_hd__a21bo_1 _23314_ (.A1(_07418_),
    .A2(_07419_),
    .B1_N(_07420_),
    .X(_07421_));
 sky130_fd_sc_hd__or2_1 _23315_ (.A(_07402_),
    .B(_07421_),
    .X(_07422_));
 sky130_fd_sc_hd__a21bo_2 _23316_ (.A1(_07402_),
    .A2(_07421_),
    .B1_N(_07422_),
    .X(_07423_));
 sky130_fd_sc_hd__a2bb2o_1 _23317_ (.A1_N(_07296_),
    .A2_N(_07423_),
    .B1(_07296_),
    .B2(_07423_),
    .X(_07424_));
 sky130_fd_sc_hd__a2bb2o_1 _23318_ (.A1_N(_07393_),
    .A2_N(_07424_),
    .B1(_07393_),
    .B2(_07424_),
    .X(_07425_));
 sky130_fd_sc_hd__o22a_1 _23319_ (.A1(_07102_),
    .A2(_07297_),
    .B1(_07265_),
    .B2(_07298_),
    .X(_07426_));
 sky130_fd_sc_hd__a2bb2o_1 _23320_ (.A1_N(_07425_),
    .A2_N(_07426_),
    .B1(_07425_),
    .B2(_07426_),
    .X(_07427_));
 sky130_fd_sc_hd__a2bb2o_1 _23321_ (.A1_N(_07360_),
    .A2_N(_07427_),
    .B1(_07360_),
    .B2(_07427_),
    .X(_07428_));
 sky130_fd_sc_hd__o22a_1 _23322_ (.A1(_07140_),
    .A2(_07299_),
    .B1(_07226_),
    .B2(_07300_),
    .X(_07429_));
 sky130_fd_sc_hd__a2bb2o_1 _23323_ (.A1_N(_07428_),
    .A2_N(_07429_),
    .B1(_07428_),
    .B2(_07429_),
    .X(_07430_));
 sky130_fd_sc_hd__a2bb2o_1 _23324_ (.A1_N(_07314_),
    .A2_N(_07430_),
    .B1(_07314_),
    .B2(_07430_),
    .X(_07431_));
 sky130_fd_sc_hd__o22a_1 _23325_ (.A1(_07301_),
    .A2(_07302_),
    .B1(_07166_),
    .B2(_07303_),
    .X(_07432_));
 sky130_fd_sc_hd__a2bb2o_1 _23326_ (.A1_N(_07431_),
    .A2_N(_07432_),
    .B1(_07431_),
    .B2(_07432_),
    .X(_07433_));
 sky130_fd_sc_hd__a2bb2o_1 _23327_ (.A1_N(_07165_),
    .A2_N(_07433_),
    .B1(_07165_),
    .B2(_07433_),
    .X(_07434_));
 sky130_fd_sc_hd__o22a_1 _23328_ (.A1(_07304_),
    .A2(_07305_),
    .B1(_07012_),
    .B2(_07306_),
    .X(_07435_));
 sky130_fd_sc_hd__or2_1 _23329_ (.A(_07434_),
    .B(_07435_),
    .X(_07436_));
 sky130_fd_sc_hd__a21bo_1 _23330_ (.A1(_07434_),
    .A2(_07435_),
    .B1_N(_07436_),
    .X(_07437_));
 sky130_fd_sc_hd__a22o_1 _23331_ (.A1(_07162_),
    .A2(_07307_),
    .B1(_07151_),
    .B2(_07308_),
    .X(_07438_));
 sky130_fd_sc_hd__o31a_1 _23332_ (.A1(_07153_),
    .A2(_07309_),
    .A3(_07160_),
    .B1(_07438_),
    .X(_07439_));
 sky130_fd_sc_hd__a2bb2oi_2 _23333_ (.A1_N(_07437_),
    .A2_N(_07439_),
    .B1(_07437_),
    .B2(_07439_),
    .Y(_02645_));
 sky130_fd_sc_hd__o22a_1 _23334_ (.A1(_07431_),
    .A2(_07432_),
    .B1(_07165_),
    .B2(_07433_),
    .X(_07440_));
 sky130_fd_sc_hd__o22a_1 _23335_ (.A1(_07316_),
    .A2(_07358_),
    .B1(_07315_),
    .B2(_07359_),
    .X(_07441_));
 sky130_fd_sc_hd__o22a_1 _23336_ (.A1(_07338_),
    .A2(_07339_),
    .B1(_07317_),
    .B2(_07340_),
    .X(_07442_));
 sky130_fd_sc_hd__or2_1 _23337_ (.A(_07441_),
    .B(_07442_),
    .X(_07443_));
 sky130_fd_sc_hd__a21bo_1 _23338_ (.A1(_07441_),
    .A2(_07442_),
    .B1_N(_07443_),
    .X(_07444_));
 sky130_fd_sc_hd__o22a_1 _23339_ (.A1(_07355_),
    .A2(_07356_),
    .B1(_07341_),
    .B2(_07357_),
    .X(_07445_));
 sky130_fd_sc_hd__o22a_1 _23340_ (.A1(_07294_),
    .A2(_07391_),
    .B1(_07361_),
    .B2(_07392_),
    .X(_07446_));
 sky130_fd_sc_hd__a21oi_2 _23341_ (.A1(_07320_),
    .A2(_07322_),
    .B1(_07319_),
    .Y(_07447_));
 sky130_fd_sc_hd__buf_1 _23342_ (.A(\pcpi_mul.rs1[26] ),
    .X(_07448_));
 sky130_fd_sc_hd__clkbuf_2 _23343_ (.A(_07448_),
    .X(_07449_));
 sky130_fd_sc_hd__clkbuf_2 _23344_ (.A(_07449_),
    .X(_07450_));
 sky130_fd_sc_hd__and4_1 _23345_ (.A(_05823_),
    .B(_13535_),
    .C(_05824_),
    .D(_07450_),
    .X(_07451_));
 sky130_fd_sc_hd__clkbuf_2 _23346_ (.A(_07196_),
    .X(_07452_));
 sky130_fd_sc_hd__buf_2 _23347_ (.A(_07452_),
    .X(_07453_));
 sky130_fd_sc_hd__o22a_1 _23348_ (.A1(_06564_),
    .A2(_07453_),
    .B1(_06753_),
    .B2(_07327_),
    .X(_07454_));
 sky130_fd_sc_hd__or2_1 _23349_ (.A(_07451_),
    .B(_07454_),
    .X(_07455_));
 sky130_fd_sc_hd__buf_1 _23350_ (.A(_05827_),
    .X(_07456_));
 sky130_fd_sc_hd__buf_1 _23351_ (.A(_07031_),
    .X(_07457_));
 sky130_fd_sc_hd__clkbuf_2 _23352_ (.A(_07457_),
    .X(_07458_));
 sky130_fd_sc_hd__clkbuf_2 _23353_ (.A(_07458_),
    .X(_07459_));
 sky130_fd_sc_hd__or2_1 _23354_ (.A(_07456_),
    .B(_07459_),
    .X(_07460_));
 sky130_fd_sc_hd__a2bb2o_1 _23355_ (.A1_N(_07455_),
    .A2_N(_07460_),
    .B1(_07455_),
    .B2(_07460_),
    .X(_07461_));
 sky130_vsdinv _23356_ (.A(\pcpi_mul.rs1[27] ),
    .Y(_07462_));
 sky130_fd_sc_hd__buf_1 _23357_ (.A(_07462_),
    .X(_07463_));
 sky130_fd_sc_hd__buf_2 _23358_ (.A(_07463_),
    .X(_07464_));
 sky130_fd_sc_hd__or2_1 _23359_ (.A(_07030_),
    .B(_07464_),
    .X(_07465_));
 sky130_fd_sc_hd__clkbuf_2 _23360_ (.A(_13541_),
    .X(_07466_));
 sky130_fd_sc_hd__and4_1 _23361_ (.A(_07186_),
    .B(_07330_),
    .C(_07189_),
    .D(_07466_),
    .X(_07467_));
 sky130_fd_sc_hd__clkbuf_2 _23362_ (.A(_07018_),
    .X(_07468_));
 sky130_fd_sc_hd__o22a_1 _23363_ (.A1(_06454_),
    .A2(_07332_),
    .B1(_06455_),
    .B2(_07468_),
    .X(_07469_));
 sky130_fd_sc_hd__or2_1 _23364_ (.A(_07467_),
    .B(_07469_),
    .X(_07470_));
 sky130_fd_sc_hd__a2bb2o_1 _23365_ (.A1_N(_07465_),
    .A2_N(_07470_),
    .B1(_07465_),
    .B2(_07470_),
    .X(_07471_));
 sky130_fd_sc_hd__o21ba_1 _23366_ (.A1(_07328_),
    .A2(_07334_),
    .B1_N(_07331_),
    .X(_07472_));
 sky130_fd_sc_hd__a2bb2o_1 _23367_ (.A1_N(_07471_),
    .A2_N(_07472_),
    .B1(_07471_),
    .B2(_07472_),
    .X(_07473_));
 sky130_fd_sc_hd__a2bb2o_1 _23368_ (.A1_N(_07461_),
    .A2_N(_07473_),
    .B1(_07461_),
    .B2(_07473_),
    .X(_07474_));
 sky130_fd_sc_hd__o22a_1 _23369_ (.A1(_07335_),
    .A2(_07336_),
    .B1(_07323_),
    .B2(_07337_),
    .X(_07475_));
 sky130_fd_sc_hd__a2bb2o_1 _23370_ (.A1_N(_07474_),
    .A2_N(_07475_),
    .B1(_07474_),
    .B2(_07475_),
    .X(_07476_));
 sky130_fd_sc_hd__a2bb2o_1 _23371_ (.A1_N(_07447_),
    .A2_N(_07476_),
    .B1(_07447_),
    .B2(_07476_),
    .X(_07477_));
 sky130_fd_sc_hd__o22a_1 _23372_ (.A1(_07345_),
    .A2(_07351_),
    .B1(_07344_),
    .B2(_07352_),
    .X(_07478_));
 sky130_fd_sc_hd__o22a_1 _23373_ (.A1(_07375_),
    .A2(_07376_),
    .B1(_07368_),
    .B2(_07377_),
    .X(_07479_));
 sky130_fd_sc_hd__o21ba_1 _23374_ (.A1(_07346_),
    .A2(_07350_),
    .B1_N(_07347_),
    .X(_07480_));
 sky130_fd_sc_hd__o21ba_1 _23375_ (.A1(_07362_),
    .A2(_07367_),
    .B1_N(_07365_),
    .X(_07481_));
 sky130_fd_sc_hd__buf_1 _23376_ (.A(_06877_),
    .X(_07482_));
 sky130_fd_sc_hd__or2_1 _23377_ (.A(_06915_),
    .B(_07482_),
    .X(_07483_));
 sky130_fd_sc_hd__buf_1 _23378_ (.A(\pcpi_mul.rs1[19] ),
    .X(_07484_));
 sky130_fd_sc_hd__buf_1 _23379_ (.A(_07484_),
    .X(_07485_));
 sky130_fd_sc_hd__and4_1 _23380_ (.A(_06923_),
    .B(_07485_),
    .C(_06924_),
    .D(_13552_),
    .X(_07486_));
 sky130_fd_sc_hd__o22a_1 _23381_ (.A1(_07055_),
    .A2(_06565_),
    .B1(_07214_),
    .B2(_06640_),
    .X(_07487_));
 sky130_fd_sc_hd__or2_1 _23382_ (.A(_07486_),
    .B(_07487_),
    .X(_07488_));
 sky130_fd_sc_hd__a2bb2o_1 _23383_ (.A1_N(_07483_),
    .A2_N(_07488_),
    .B1(_07483_),
    .B2(_07488_),
    .X(_07489_));
 sky130_fd_sc_hd__a2bb2o_1 _23384_ (.A1_N(_07481_),
    .A2_N(_07489_),
    .B1(_07481_),
    .B2(_07489_),
    .X(_07490_));
 sky130_fd_sc_hd__a2bb2o_1 _23385_ (.A1_N(_07480_),
    .A2_N(_07490_),
    .B1(_07480_),
    .B2(_07490_),
    .X(_07491_));
 sky130_fd_sc_hd__a2bb2o_1 _23386_ (.A1_N(_07479_),
    .A2_N(_07491_),
    .B1(_07479_),
    .B2(_07491_),
    .X(_07492_));
 sky130_fd_sc_hd__a2bb2o_1 _23387_ (.A1_N(_07478_),
    .A2_N(_07492_),
    .B1(_07478_),
    .B2(_07492_),
    .X(_07493_));
 sky130_fd_sc_hd__o22a_1 _23388_ (.A1(_07343_),
    .A2(_07353_),
    .B1(_07342_),
    .B2(_07354_),
    .X(_07494_));
 sky130_fd_sc_hd__a2bb2o_1 _23389_ (.A1_N(_07493_),
    .A2_N(_07494_),
    .B1(_07493_),
    .B2(_07494_),
    .X(_07495_));
 sky130_fd_sc_hd__a2bb2o_1 _23390_ (.A1_N(_07477_),
    .A2_N(_07495_),
    .B1(_07477_),
    .B2(_07495_),
    .X(_07496_));
 sky130_fd_sc_hd__a2bb2o_1 _23391_ (.A1_N(_07446_),
    .A2_N(_07496_),
    .B1(_07446_),
    .B2(_07496_),
    .X(_07497_));
 sky130_fd_sc_hd__a2bb2o_1 _23392_ (.A1_N(_07445_),
    .A2_N(_07497_),
    .B1(_07445_),
    .B2(_07497_),
    .X(_07498_));
 sky130_fd_sc_hd__o22a_1 _23393_ (.A1(_07388_),
    .A2(_07389_),
    .B1(_07378_),
    .B2(_07390_),
    .X(_07499_));
 sky130_fd_sc_hd__or2_1 _23394_ (.A(_07105_),
    .B(_06339_),
    .X(_07500_));
 sky130_fd_sc_hd__buf_1 _23395_ (.A(\pcpi_mul.rs1[17] ),
    .X(_07501_));
 sky130_fd_sc_hd__and4_1 _23396_ (.A(_06824_),
    .B(_06583_),
    .C(_06825_),
    .D(_07501_),
    .X(_07502_));
 sky130_fd_sc_hd__o22a_1 _23397_ (.A1(_06522_),
    .A2(_06580_),
    .B1(_06523_),
    .B2(_06916_),
    .X(_07503_));
 sky130_fd_sc_hd__or2_1 _23398_ (.A(_07502_),
    .B(_07503_),
    .X(_07504_));
 sky130_fd_sc_hd__a2bb2o_1 _23399_ (.A1_N(_07500_),
    .A2_N(_07504_),
    .B1(_07500_),
    .B2(_07504_),
    .X(_07505_));
 sky130_fd_sc_hd__or2_1 _23400_ (.A(_06967_),
    .B(_06457_),
    .X(_07506_));
 sky130_fd_sc_hd__and4_1 _23401_ (.A(_07234_),
    .B(_07371_),
    .C(_07235_),
    .D(_06342_),
    .X(_07507_));
 sky130_fd_sc_hd__o22a_1 _23402_ (.A1(_07237_),
    .A2(_05836_),
    .B1(_07238_),
    .B2(_06598_),
    .X(_07508_));
 sky130_fd_sc_hd__or2_1 _23403_ (.A(_07507_),
    .B(_07508_),
    .X(_07509_));
 sky130_fd_sc_hd__a2bb2o_1 _23404_ (.A1_N(_07506_),
    .A2_N(_07509_),
    .B1(_07506_),
    .B2(_07509_),
    .X(_07510_));
 sky130_fd_sc_hd__o21ba_1 _23405_ (.A1(_07370_),
    .A2(_07374_),
    .B1_N(_07372_),
    .X(_07511_));
 sky130_fd_sc_hd__a2bb2o_1 _23406_ (.A1_N(_07510_),
    .A2_N(_07511_),
    .B1(_07510_),
    .B2(_07511_),
    .X(_07512_));
 sky130_fd_sc_hd__a2bb2o_2 _23407_ (.A1_N(_07505_),
    .A2_N(_07512_),
    .B1(_07505_),
    .B2(_07512_),
    .X(_07513_));
 sky130_fd_sc_hd__o21ba_1 _23408_ (.A1(_07381_),
    .A2(_07385_),
    .B1_N(_07382_),
    .X(_07514_));
 sky130_fd_sc_hd__o21ba_1 _23409_ (.A1(_07404_),
    .A2(_07409_),
    .B1_N(_07407_),
    .X(_07515_));
 sky130_fd_sc_hd__buf_1 _23410_ (.A(_05998_),
    .X(_07516_));
 sky130_fd_sc_hd__or2_1 _23411_ (.A(_07516_),
    .B(_05928_),
    .X(_07517_));
 sky130_fd_sc_hd__and4_1 _23412_ (.A(_07248_),
    .B(_06974_),
    .C(_07250_),
    .D(_06486_),
    .X(_07518_));
 sky130_fd_sc_hd__o22a_1 _23413_ (.A1(_07383_),
    .A2(_05947_),
    .B1(_07254_),
    .B2(_05817_),
    .X(_07519_));
 sky130_fd_sc_hd__or2_1 _23414_ (.A(_07518_),
    .B(_07519_),
    .X(_07520_));
 sky130_fd_sc_hd__a2bb2o_1 _23415_ (.A1_N(_07517_),
    .A2_N(_07520_),
    .B1(_07517_),
    .B2(_07520_),
    .X(_07521_));
 sky130_fd_sc_hd__a2bb2o_1 _23416_ (.A1_N(_07515_),
    .A2_N(_07521_),
    .B1(_07515_),
    .B2(_07521_),
    .X(_07522_));
 sky130_fd_sc_hd__a2bb2o_1 _23417_ (.A1_N(_07514_),
    .A2_N(_07522_),
    .B1(_07514_),
    .B2(_07522_),
    .X(_07523_));
 sky130_fd_sc_hd__o22a_1 _23418_ (.A1(_07380_),
    .A2(_07386_),
    .B1(_07379_),
    .B2(_07387_),
    .X(_07524_));
 sky130_fd_sc_hd__a2bb2o_1 _23419_ (.A1_N(_07523_),
    .A2_N(_07524_),
    .B1(_07523_),
    .B2(_07524_),
    .X(_07525_));
 sky130_fd_sc_hd__a2bb2o_1 _23420_ (.A1_N(_07513_),
    .A2_N(_07525_),
    .B1(_07513_),
    .B2(_07525_),
    .X(_07526_));
 sky130_fd_sc_hd__a2bb2o_1 _23421_ (.A1_N(_07420_),
    .A2_N(_07526_),
    .B1(_07420_),
    .B2(_07526_),
    .X(_07527_));
 sky130_fd_sc_hd__a2bb2o_1 _23422_ (.A1_N(_07499_),
    .A2_N(_07527_),
    .B1(_07499_),
    .B2(_07527_),
    .X(_07528_));
 sky130_vsdinv _23423_ (.A(\pcpi_mul.rs2[27] ),
    .Y(_07529_));
 sky130_fd_sc_hd__buf_1 _23424_ (.A(_07529_),
    .X(_07530_));
 sky130_fd_sc_hd__clkbuf_2 _23425_ (.A(_07530_),
    .X(_07531_));
 sky130_fd_sc_hd__buf_4 _23426_ (.A(_07531_),
    .X(_07532_));
 sky130_fd_sc_hd__or2_2 _23427_ (.A(_07532_),
    .B(_05152_),
    .X(_07533_));
 sky130_fd_sc_hd__or2_1 _23428_ (.A(_07072_),
    .B(_05339_),
    .X(_07534_));
 sky130_fd_sc_hd__o22a_1 _23429_ (.A1(_07397_),
    .A2(_05296_),
    .B1(_07266_),
    .B2(_06187_),
    .X(_07535_));
 sky130_fd_sc_hd__buf_1 _23430_ (.A(\pcpi_mul.rs2[26] ),
    .X(_07536_));
 sky130_fd_sc_hd__and4_1 _23431_ (.A(_07536_),
    .B(_06695_),
    .C(_07395_),
    .D(_05346_),
    .X(_07537_));
 sky130_fd_sc_hd__or2_1 _23432_ (.A(_07535_),
    .B(_07537_),
    .X(_07538_));
 sky130_fd_sc_hd__a2bb2o_1 _23433_ (.A1_N(_07534_),
    .A2_N(_07538_),
    .B1(_07534_),
    .B2(_07538_),
    .X(_07539_));
 sky130_fd_sc_hd__o21ba_1 _23434_ (.A1(_07394_),
    .A2(_07399_),
    .B1_N(_07396_),
    .X(_07540_));
 sky130_fd_sc_hd__or2_2 _23435_ (.A(_07539_),
    .B(_07540_),
    .X(_07541_));
 sky130_fd_sc_hd__a21bo_1 _23436_ (.A1(_07539_),
    .A2(_07540_),
    .B1_N(_07541_),
    .X(_07542_));
 sky130_fd_sc_hd__or2_2 _23437_ (.A(_07533_),
    .B(_07542_),
    .X(_07543_));
 sky130_fd_sc_hd__a21bo_1 _23438_ (.A1(_07533_),
    .A2(_07542_),
    .B1_N(_07543_),
    .X(_07544_));
 sky130_fd_sc_hd__o22a_1 _23439_ (.A1(_07415_),
    .A2(_07416_),
    .B1(_07410_),
    .B2(_07417_),
    .X(_07545_));
 sky130_fd_sc_hd__buf_1 _23440_ (.A(_06396_),
    .X(_07546_));
 sky130_fd_sc_hd__or2_1 _23441_ (.A(_07546_),
    .B(_05731_),
    .X(_07547_));
 sky130_fd_sc_hd__o22a_1 _23442_ (.A1(_07281_),
    .A2(_07277_),
    .B1(_07282_),
    .B2(_06983_),
    .X(_07548_));
 sky130_fd_sc_hd__buf_1 _23443_ (.A(_06694_),
    .X(_07549_));
 sky130_fd_sc_hd__and4_1 _23444_ (.A(_07549_),
    .B(_06303_),
    .C(_07406_),
    .D(_05846_),
    .X(_07550_));
 sky130_fd_sc_hd__or2_1 _23445_ (.A(_07548_),
    .B(_07550_),
    .X(_07551_));
 sky130_fd_sc_hd__a2bb2o_1 _23446_ (.A1_N(_07547_),
    .A2_N(_07551_),
    .B1(_07547_),
    .B2(_07551_),
    .X(_07552_));
 sky130_fd_sc_hd__or2_1 _23447_ (.A(_06687_),
    .B(_06003_),
    .X(_07553_));
 sky130_fd_sc_hd__and4_1 _23448_ (.A(_13096_),
    .B(_07085_),
    .C(_13101_),
    .D(_13608_),
    .X(_07554_));
 sky130_fd_sc_hd__o22a_1 _23449_ (.A1(_06948_),
    .A2(_05798_),
    .B1(_06805_),
    .B2(_06544_),
    .X(_07555_));
 sky130_fd_sc_hd__or2_1 _23450_ (.A(_07554_),
    .B(_07555_),
    .X(_07556_));
 sky130_fd_sc_hd__a2bb2o_1 _23451_ (.A1_N(_07553_),
    .A2_N(_07556_),
    .B1(_07553_),
    .B2(_07556_),
    .X(_07557_));
 sky130_fd_sc_hd__o21ba_1 _23452_ (.A1(_07411_),
    .A2(_07414_),
    .B1_N(_07412_),
    .X(_07558_));
 sky130_fd_sc_hd__a2bb2o_1 _23453_ (.A1_N(_07557_),
    .A2_N(_07558_),
    .B1(_07557_),
    .B2(_07558_),
    .X(_07559_));
 sky130_fd_sc_hd__a2bb2o_1 _23454_ (.A1_N(_07552_),
    .A2_N(_07559_),
    .B1(_07552_),
    .B2(_07559_),
    .X(_07560_));
 sky130_fd_sc_hd__a2bb2o_1 _23455_ (.A1_N(_07401_),
    .A2_N(_07560_),
    .B1(_07401_),
    .B2(_07560_),
    .X(_07561_));
 sky130_fd_sc_hd__a2bb2o_1 _23456_ (.A1_N(_07545_),
    .A2_N(_07561_),
    .B1(_07545_),
    .B2(_07561_),
    .X(_07562_));
 sky130_fd_sc_hd__or2_1 _23457_ (.A(_07544_),
    .B(_07562_),
    .X(_07563_));
 sky130_fd_sc_hd__a21bo_1 _23458_ (.A1(_07544_),
    .A2(_07562_),
    .B1_N(_07563_),
    .X(_07564_));
 sky130_fd_sc_hd__a2bb2o_1 _23459_ (.A1_N(_07422_),
    .A2_N(_07564_),
    .B1(_07422_),
    .B2(_07564_),
    .X(_07565_));
 sky130_fd_sc_hd__a2bb2o_2 _23460_ (.A1_N(_07528_),
    .A2_N(_07565_),
    .B1(_07528_),
    .B2(_07565_),
    .X(_07566_));
 sky130_fd_sc_hd__o22a_1 _23461_ (.A1(_07296_),
    .A2(_07423_),
    .B1(_07393_),
    .B2(_07424_),
    .X(_07567_));
 sky130_fd_sc_hd__a2bb2o_1 _23462_ (.A1_N(_07566_),
    .A2_N(_07567_),
    .B1(_07566_),
    .B2(_07567_),
    .X(_07568_));
 sky130_fd_sc_hd__a2bb2o_1 _23463_ (.A1_N(_07498_),
    .A2_N(_07568_),
    .B1(_07498_),
    .B2(_07568_),
    .X(_07569_));
 sky130_fd_sc_hd__o22a_1 _23464_ (.A1(_07425_),
    .A2(_07426_),
    .B1(_07360_),
    .B2(_07427_),
    .X(_07570_));
 sky130_fd_sc_hd__a2bb2o_1 _23465_ (.A1_N(_07569_),
    .A2_N(_07570_),
    .B1(_07569_),
    .B2(_07570_),
    .X(_07571_));
 sky130_fd_sc_hd__a2bb2o_1 _23466_ (.A1_N(_07444_),
    .A2_N(_07571_),
    .B1(_07444_),
    .B2(_07571_),
    .X(_07572_));
 sky130_fd_sc_hd__o22a_1 _23467_ (.A1(_07428_),
    .A2(_07429_),
    .B1(_07314_),
    .B2(_07430_),
    .X(_07573_));
 sky130_fd_sc_hd__a2bb2o_1 _23468_ (.A1_N(_07572_),
    .A2_N(_07573_),
    .B1(_07572_),
    .B2(_07573_),
    .X(_07574_));
 sky130_fd_sc_hd__a2bb2o_1 _23469_ (.A1_N(_07313_),
    .A2_N(_07574_),
    .B1(_07313_),
    .B2(_07574_),
    .X(_07575_));
 sky130_fd_sc_hd__and2_1 _23470_ (.A(_07440_),
    .B(_07575_),
    .X(_07576_));
 sky130_fd_sc_hd__or2_1 _23471_ (.A(_07440_),
    .B(_07575_),
    .X(_07577_));
 sky130_fd_sc_hd__or2b_1 _23472_ (.A(_07576_),
    .B_N(_07577_),
    .X(_07578_));
 sky130_fd_sc_hd__o21ai_1 _23473_ (.A1(_07437_),
    .A2(_07439_),
    .B1(_07436_),
    .Y(_07579_));
 sky130_fd_sc_hd__a2bb2o_1 _23474_ (.A1_N(_07578_),
    .A2_N(_07579_),
    .B1(_07578_),
    .B2(_07579_),
    .X(_02646_));
 sky130_fd_sc_hd__o22a_1 _23475_ (.A1(_07446_),
    .A2(_07496_),
    .B1(_07445_),
    .B2(_07497_),
    .X(_07580_));
 sky130_fd_sc_hd__o22a_1 _23476_ (.A1(_07474_),
    .A2(_07475_),
    .B1(_07447_),
    .B2(_07476_),
    .X(_07581_));
 sky130_fd_sc_hd__or2_1 _23477_ (.A(_07580_),
    .B(_07581_),
    .X(_07582_));
 sky130_fd_sc_hd__a21bo_1 _23478_ (.A1(_07580_),
    .A2(_07581_),
    .B1_N(_07582_),
    .X(_07583_));
 sky130_fd_sc_hd__o22a_1 _23479_ (.A1(_07493_),
    .A2(_07494_),
    .B1(_07477_),
    .B2(_07495_),
    .X(_07584_));
 sky130_fd_sc_hd__o22a_2 _23480_ (.A1(_07420_),
    .A2(_07526_),
    .B1(_07499_),
    .B2(_07527_),
    .X(_07585_));
 sky130_fd_sc_hd__o21ba_1 _23481_ (.A1(_07455_),
    .A2(_07460_),
    .B1_N(_07451_),
    .X(_07586_));
 sky130_fd_sc_hd__buf_1 _23482_ (.A(\pcpi_mul.rs1[27] ),
    .X(_07587_));
 sky130_fd_sc_hd__clkbuf_2 _23483_ (.A(_07587_),
    .X(_07588_));
 sky130_fd_sc_hd__and4_1 _23484_ (.A(_05823_),
    .B(_07450_),
    .C(_05824_),
    .D(_07588_),
    .X(_07589_));
 sky130_fd_sc_hd__o22a_1 _23485_ (.A1(_05816_),
    .A2(_07327_),
    .B1(_06753_),
    .B2(_07464_),
    .X(_07590_));
 sky130_fd_sc_hd__or2_1 _23486_ (.A(_07589_),
    .B(_07590_),
    .X(_07591_));
 sky130_fd_sc_hd__or2_1 _23487_ (.A(_07456_),
    .B(_07198_),
    .X(_07592_));
 sky130_fd_sc_hd__a2bb2o_1 _23488_ (.A1_N(_07591_),
    .A2_N(_07592_),
    .B1(_07591_),
    .B2(_07592_),
    .X(_07593_));
 sky130_vsdinv _23489_ (.A(\pcpi_mul.rs1[28] ),
    .Y(_07594_));
 sky130_fd_sc_hd__buf_1 _23490_ (.A(_07594_),
    .X(_07595_));
 sky130_fd_sc_hd__clkbuf_2 _23491_ (.A(_07595_),
    .X(_07596_));
 sky130_fd_sc_hd__or2_1 _23492_ (.A(_07030_),
    .B(_07596_),
    .X(_07597_));
 sky130_fd_sc_hd__clkbuf_2 _23493_ (.A(_13538_),
    .X(_07598_));
 sky130_fd_sc_hd__and4_1 _23494_ (.A(_06897_),
    .B(_07466_),
    .C(_06900_),
    .D(_07598_),
    .X(_07599_));
 sky130_fd_sc_hd__o22a_1 _23495_ (.A1(_06454_),
    .A2(_06891_),
    .B1(_06455_),
    .B2(_07033_),
    .X(_07600_));
 sky130_fd_sc_hd__or2_1 _23496_ (.A(_07599_),
    .B(_07600_),
    .X(_07601_));
 sky130_fd_sc_hd__a2bb2o_1 _23497_ (.A1_N(_07597_),
    .A2_N(_07601_),
    .B1(_07597_),
    .B2(_07601_),
    .X(_07602_));
 sky130_fd_sc_hd__o21ba_1 _23498_ (.A1(_07465_),
    .A2(_07470_),
    .B1_N(_07467_),
    .X(_07603_));
 sky130_fd_sc_hd__a2bb2o_1 _23499_ (.A1_N(_07602_),
    .A2_N(_07603_),
    .B1(_07602_),
    .B2(_07603_),
    .X(_07604_));
 sky130_fd_sc_hd__a2bb2o_1 _23500_ (.A1_N(_07593_),
    .A2_N(_07604_),
    .B1(_07593_),
    .B2(_07604_),
    .X(_07605_));
 sky130_fd_sc_hd__o22a_1 _23501_ (.A1(_07471_),
    .A2(_07472_),
    .B1(_07461_),
    .B2(_07473_),
    .X(_07606_));
 sky130_fd_sc_hd__a2bb2o_1 _23502_ (.A1_N(_07605_),
    .A2_N(_07606_),
    .B1(_07605_),
    .B2(_07606_),
    .X(_07607_));
 sky130_fd_sc_hd__a2bb2o_1 _23503_ (.A1_N(_07586_),
    .A2_N(_07607_),
    .B1(_07586_),
    .B2(_07607_),
    .X(_07608_));
 sky130_fd_sc_hd__o22a_1 _23504_ (.A1(_07481_),
    .A2(_07489_),
    .B1(_07480_),
    .B2(_07490_),
    .X(_07609_));
 sky130_fd_sc_hd__o22a_1 _23505_ (.A1(_07510_),
    .A2(_07511_),
    .B1(_07505_),
    .B2(_07512_),
    .X(_07610_));
 sky130_fd_sc_hd__o21ba_1 _23506_ (.A1(_07483_),
    .A2(_07488_),
    .B1_N(_07486_),
    .X(_07611_));
 sky130_fd_sc_hd__o21ba_1 _23507_ (.A1(_07500_),
    .A2(_07504_),
    .B1_N(_07502_),
    .X(_07612_));
 sky130_fd_sc_hd__clkbuf_2 _23508_ (.A(_06880_),
    .X(_07613_));
 sky130_fd_sc_hd__or2_1 _23509_ (.A(_05424_),
    .B(_07613_),
    .X(_07614_));
 sky130_fd_sc_hd__and4_1 _23510_ (.A(_07057_),
    .B(_13552_),
    .C(_07058_),
    .D(_13549_),
    .X(_07615_));
 sky130_fd_sc_hd__o22a_1 _23511_ (.A1(_07055_),
    .A2(_06574_),
    .B1(_07214_),
    .B2(_06877_),
    .X(_07616_));
 sky130_fd_sc_hd__or2_1 _23512_ (.A(_07615_),
    .B(_07616_),
    .X(_07617_));
 sky130_fd_sc_hd__a2bb2o_1 _23513_ (.A1_N(_07614_),
    .A2_N(_07617_),
    .B1(_07614_),
    .B2(_07617_),
    .X(_07618_));
 sky130_fd_sc_hd__a2bb2o_1 _23514_ (.A1_N(_07612_),
    .A2_N(_07618_),
    .B1(_07612_),
    .B2(_07618_),
    .X(_07619_));
 sky130_fd_sc_hd__a2bb2o_1 _23515_ (.A1_N(_07611_),
    .A2_N(_07619_),
    .B1(_07611_),
    .B2(_07619_),
    .X(_07620_));
 sky130_fd_sc_hd__a2bb2o_1 _23516_ (.A1_N(_07610_),
    .A2_N(_07620_),
    .B1(_07610_),
    .B2(_07620_),
    .X(_07621_));
 sky130_fd_sc_hd__a2bb2o_1 _23517_ (.A1_N(_07609_),
    .A2_N(_07621_),
    .B1(_07609_),
    .B2(_07621_),
    .X(_07622_));
 sky130_fd_sc_hd__o22a_1 _23518_ (.A1(_07479_),
    .A2(_07491_),
    .B1(_07478_),
    .B2(_07492_),
    .X(_07623_));
 sky130_fd_sc_hd__a2bb2o_1 _23519_ (.A1_N(_07622_),
    .A2_N(_07623_),
    .B1(_07622_),
    .B2(_07623_),
    .X(_07624_));
 sky130_fd_sc_hd__a2bb2o_1 _23520_ (.A1_N(_07608_),
    .A2_N(_07624_),
    .B1(_07608_),
    .B2(_07624_),
    .X(_07625_));
 sky130_fd_sc_hd__a2bb2o_1 _23521_ (.A1_N(_07585_),
    .A2_N(_07625_),
    .B1(_07585_),
    .B2(_07625_),
    .X(_07626_));
 sky130_fd_sc_hd__a2bb2o_1 _23522_ (.A1_N(_07584_),
    .A2_N(_07626_),
    .B1(_07584_),
    .B2(_07626_),
    .X(_07627_));
 sky130_fd_sc_hd__o22a_1 _23523_ (.A1(_07523_),
    .A2(_07524_),
    .B1(_07513_),
    .B2(_07525_),
    .X(_07628_));
 sky130_fd_sc_hd__o22a_1 _23524_ (.A1(_07401_),
    .A2(_07560_),
    .B1(_07545_),
    .B2(_07561_),
    .X(_07629_));
 sky130_fd_sc_hd__or2_1 _23525_ (.A(_07105_),
    .B(_07036_),
    .X(_07630_));
 sky130_fd_sc_hd__o22a_1 _23526_ (.A1(_07107_),
    .A2(_06226_),
    .B1(_07108_),
    .B2(_06437_),
    .X(_07631_));
 sky130_fd_sc_hd__and4_1 _23527_ (.A(_06525_),
    .B(_07501_),
    .C(_06527_),
    .D(_06898_),
    .X(_07632_));
 sky130_fd_sc_hd__or2_1 _23528_ (.A(_07631_),
    .B(_07632_),
    .X(_07633_));
 sky130_fd_sc_hd__a2bb2o_1 _23529_ (.A1_N(_07630_),
    .A2_N(_07633_),
    .B1(_07630_),
    .B2(_07633_),
    .X(_07634_));
 sky130_fd_sc_hd__or2_1 _23530_ (.A(_06967_),
    .B(_06581_),
    .X(_07635_));
 sky130_fd_sc_hd__and4_1 _23531_ (.A(_06972_),
    .B(_06342_),
    .C(_06973_),
    .D(_06462_),
    .X(_07636_));
 sky130_fd_sc_hd__o22a_1 _23532_ (.A1(_06830_),
    .A2(_05943_),
    .B1(_07238_),
    .B2(_06668_),
    .X(_07637_));
 sky130_fd_sc_hd__or2_1 _23533_ (.A(_07636_),
    .B(_07637_),
    .X(_07638_));
 sky130_fd_sc_hd__a2bb2o_1 _23534_ (.A1_N(_07635_),
    .A2_N(_07638_),
    .B1(_07635_),
    .B2(_07638_),
    .X(_07639_));
 sky130_fd_sc_hd__o21ba_1 _23535_ (.A1(_07506_),
    .A2(_07509_),
    .B1_N(_07507_),
    .X(_07640_));
 sky130_fd_sc_hd__a2bb2o_1 _23536_ (.A1_N(_07639_),
    .A2_N(_07640_),
    .B1(_07639_),
    .B2(_07640_),
    .X(_07641_));
 sky130_fd_sc_hd__a2bb2o_2 _23537_ (.A1_N(_07634_),
    .A2_N(_07641_),
    .B1(_07634_),
    .B2(_07641_),
    .X(_07642_));
 sky130_fd_sc_hd__o21ba_1 _23538_ (.A1(_07517_),
    .A2(_07520_),
    .B1_N(_07518_),
    .X(_07643_));
 sky130_fd_sc_hd__o21ba_1 _23539_ (.A1(_07547_),
    .A2(_07551_),
    .B1_N(_07550_),
    .X(_07644_));
 sky130_fd_sc_hd__or2_1 _23540_ (.A(_07516_),
    .B(_06479_),
    .X(_07645_));
 sky130_fd_sc_hd__and4_1 _23541_ (.A(_07248_),
    .B(_07117_),
    .C(_07250_),
    .D(_06602_),
    .X(_07646_));
 sky130_fd_sc_hd__o22a_1 _23542_ (.A1(_07253_),
    .A2(_06704_),
    .B1(_07254_),
    .B2(_06356_),
    .X(_07647_));
 sky130_fd_sc_hd__or2_1 _23543_ (.A(_07646_),
    .B(_07647_),
    .X(_07648_));
 sky130_fd_sc_hd__a2bb2o_1 _23544_ (.A1_N(_07645_),
    .A2_N(_07648_),
    .B1(_07645_),
    .B2(_07648_),
    .X(_07649_));
 sky130_fd_sc_hd__a2bb2o_1 _23545_ (.A1_N(_07644_),
    .A2_N(_07649_),
    .B1(_07644_),
    .B2(_07649_),
    .X(_07650_));
 sky130_fd_sc_hd__a2bb2o_1 _23546_ (.A1_N(_07643_),
    .A2_N(_07650_),
    .B1(_07643_),
    .B2(_07650_),
    .X(_07651_));
 sky130_fd_sc_hd__o22a_1 _23547_ (.A1(_07515_),
    .A2(_07521_),
    .B1(_07514_),
    .B2(_07522_),
    .X(_07652_));
 sky130_fd_sc_hd__a2bb2o_1 _23548_ (.A1_N(_07651_),
    .A2_N(_07652_),
    .B1(_07651_),
    .B2(_07652_),
    .X(_07653_));
 sky130_fd_sc_hd__a2bb2o_1 _23549_ (.A1_N(_07642_),
    .A2_N(_07653_),
    .B1(_07642_),
    .B2(_07653_),
    .X(_07654_));
 sky130_fd_sc_hd__a2bb2o_1 _23550_ (.A1_N(_07629_),
    .A2_N(_07654_),
    .B1(_07629_),
    .B2(_07654_),
    .X(_07655_));
 sky130_fd_sc_hd__a2bb2o_1 _23551_ (.A1_N(_07628_),
    .A2_N(_07655_),
    .B1(_07628_),
    .B2(_07655_),
    .X(_07656_));
 sky130_fd_sc_hd__o22a_1 _23552_ (.A1(_07557_),
    .A2(_07558_),
    .B1(_07552_),
    .B2(_07559_),
    .X(_07657_));
 sky130_fd_sc_hd__or2_1 _23553_ (.A(_07078_),
    .B(_06399_),
    .X(_07658_));
 sky130_fd_sc_hd__o22a_1 _23554_ (.A1(_07281_),
    .A2(_05841_),
    .B1(_07282_),
    .B2(_05730_),
    .X(_07659_));
 sky130_fd_sc_hd__and4_1 _23555_ (.A(_07084_),
    .B(_05846_),
    .C(_13111_),
    .D(_05848_),
    .X(_07660_));
 sky130_fd_sc_hd__or2_1 _23556_ (.A(_07659_),
    .B(_07660_),
    .X(_07661_));
 sky130_fd_sc_hd__a2bb2o_1 _23557_ (.A1_N(_07658_),
    .A2_N(_07661_),
    .B1(_07658_),
    .B2(_07661_),
    .X(_07662_));
 sky130_fd_sc_hd__buf_2 _23558_ (.A(_06686_),
    .X(_07663_));
 sky130_fd_sc_hd__or2_1 _23559_ (.A(_07663_),
    .B(_07278_),
    .X(_07664_));
 sky130_fd_sc_hd__buf_1 _23560_ (.A(_06948_),
    .X(_07665_));
 sky130_fd_sc_hd__o22a_1 _23561_ (.A1(_07665_),
    .A2(_06201_),
    .B1(_06801_),
    .B2(_06003_),
    .X(_07666_));
 sky130_fd_sc_hd__buf_1 _23562_ (.A(_07092_),
    .X(_07667_));
 sky130_fd_sc_hd__buf_1 _23563_ (.A(_06950_),
    .X(_07668_));
 sky130_fd_sc_hd__and4_1 _23564_ (.A(_07667_),
    .B(_07086_),
    .C(_07668_),
    .D(_05872_),
    .X(_07669_));
 sky130_fd_sc_hd__or2_1 _23565_ (.A(_07666_),
    .B(_07669_),
    .X(_07670_));
 sky130_fd_sc_hd__a2bb2o_1 _23566_ (.A1_N(_07664_),
    .A2_N(_07670_),
    .B1(_07664_),
    .B2(_07670_),
    .X(_07671_));
 sky130_fd_sc_hd__o21ba_1 _23567_ (.A1(_07553_),
    .A2(_07556_),
    .B1_N(_07554_),
    .X(_07672_));
 sky130_fd_sc_hd__a2bb2o_1 _23568_ (.A1_N(_07671_),
    .A2_N(_07672_),
    .B1(_07671_),
    .B2(_07672_),
    .X(_07673_));
 sky130_fd_sc_hd__a2bb2o_1 _23569_ (.A1_N(_07662_),
    .A2_N(_07673_),
    .B1(_07662_),
    .B2(_07673_),
    .X(_07674_));
 sky130_fd_sc_hd__a2bb2o_1 _23570_ (.A1_N(_07541_),
    .A2_N(_07674_),
    .B1(_07541_),
    .B2(_07674_),
    .X(_07675_));
 sky130_fd_sc_hd__a2bb2o_1 _23571_ (.A1_N(_07657_),
    .A2_N(_07675_),
    .B1(_07657_),
    .B2(_07675_),
    .X(_07676_));
 sky130_vsdinv _23572_ (.A(\pcpi_mul.rs2[28] ),
    .Y(_07677_));
 sky130_fd_sc_hd__buf_1 _23573_ (.A(_07677_),
    .X(_07678_));
 sky130_fd_sc_hd__clkbuf_2 _23574_ (.A(_07678_),
    .X(_07679_));
 sky130_fd_sc_hd__clkbuf_4 _23575_ (.A(_07679_),
    .X(_07680_));
 sky130_fd_sc_hd__clkbuf_2 _23576_ (.A(_07529_),
    .X(_07681_));
 sky130_fd_sc_hd__clkbuf_4 _23577_ (.A(_07681_),
    .X(_07682_));
 sky130_fd_sc_hd__o22a_2 _23578_ (.A1(_07680_),
    .A2(_05151_),
    .B1(_07682_),
    .B2(_05299_),
    .X(_07683_));
 sky130_fd_sc_hd__buf_2 _23579_ (.A(_07678_),
    .X(_07684_));
 sky130_fd_sc_hd__or4_4 _23580_ (.A(_07684_),
    .B(_05459_),
    .C(_07530_),
    .D(_05792_),
    .X(_07685_));
 sky130_fd_sc_hd__or2b_1 _23581_ (.A(_07683_),
    .B_N(_07685_),
    .X(_07686_));
 sky130_fd_sc_hd__o21ba_1 _23582_ (.A1(_07534_),
    .A2(_07538_),
    .B1_N(_07537_),
    .X(_07687_));
 sky130_fd_sc_hd__buf_1 _23583_ (.A(_07072_),
    .X(_07688_));
 sky130_fd_sc_hd__or2_1 _23584_ (.A(_07688_),
    .B(_05799_),
    .X(_07689_));
 sky130_fd_sc_hd__buf_1 _23585_ (.A(_07397_),
    .X(_07690_));
 sky130_fd_sc_hd__buf_1 _23586_ (.A(_07266_),
    .X(_07691_));
 sky130_fd_sc_hd__o22a_1 _23587_ (.A1(_07690_),
    .A2(_06187_),
    .B1(_07691_),
    .B2(_05803_),
    .X(_07692_));
 sky130_fd_sc_hd__and4_2 _23588_ (.A(_07536_),
    .B(_05806_),
    .C(_07395_),
    .D(_06204_),
    .X(_07693_));
 sky130_fd_sc_hd__or2_1 _23589_ (.A(_07692_),
    .B(_07693_),
    .X(_07694_));
 sky130_fd_sc_hd__a2bb2o_1 _23590_ (.A1_N(_07689_),
    .A2_N(_07694_),
    .B1(_07689_),
    .B2(_07694_),
    .X(_07695_));
 sky130_fd_sc_hd__or2_1 _23591_ (.A(_07687_),
    .B(_07695_),
    .X(_07696_));
 sky130_fd_sc_hd__a21bo_1 _23592_ (.A1(_07687_),
    .A2(_07695_),
    .B1_N(_07696_),
    .X(_07697_));
 sky130_fd_sc_hd__or2_1 _23593_ (.A(_07686_),
    .B(_07697_),
    .X(_07698_));
 sky130_fd_sc_hd__a21bo_1 _23594_ (.A1(_07686_),
    .A2(_07697_),
    .B1_N(_07698_),
    .X(_07699_));
 sky130_fd_sc_hd__a2bb2o_1 _23595_ (.A1_N(_07543_),
    .A2_N(_07699_),
    .B1(_07543_),
    .B2(_07699_),
    .X(_07700_));
 sky130_fd_sc_hd__a2bb2o_1 _23596_ (.A1_N(_07676_),
    .A2_N(_07700_),
    .B1(_07676_),
    .B2(_07700_),
    .X(_07701_));
 sky130_fd_sc_hd__a2bb2o_1 _23597_ (.A1_N(_07563_),
    .A2_N(_07701_),
    .B1(_07563_),
    .B2(_07701_),
    .X(_07702_));
 sky130_fd_sc_hd__a2bb2o_2 _23598_ (.A1_N(_07656_),
    .A2_N(_07702_),
    .B1(_07656_),
    .B2(_07702_),
    .X(_07703_));
 sky130_fd_sc_hd__o22a_2 _23599_ (.A1(_07422_),
    .A2(_07564_),
    .B1(_07528_),
    .B2(_07565_),
    .X(_07704_));
 sky130_fd_sc_hd__a2bb2o_1 _23600_ (.A1_N(_07703_),
    .A2_N(_07704_),
    .B1(_07703_),
    .B2(_07704_),
    .X(_07705_));
 sky130_fd_sc_hd__a2bb2o_1 _23601_ (.A1_N(_07627_),
    .A2_N(_07705_),
    .B1(_07627_),
    .B2(_07705_),
    .X(_07706_));
 sky130_fd_sc_hd__o22a_1 _23602_ (.A1(_07566_),
    .A2(_07567_),
    .B1(_07498_),
    .B2(_07568_),
    .X(_07707_));
 sky130_fd_sc_hd__a2bb2o_1 _23603_ (.A1_N(_07706_),
    .A2_N(_07707_),
    .B1(_07706_),
    .B2(_07707_),
    .X(_07708_));
 sky130_fd_sc_hd__a2bb2o_1 _23604_ (.A1_N(_07583_),
    .A2_N(_07708_),
    .B1(_07583_),
    .B2(_07708_),
    .X(_07709_));
 sky130_fd_sc_hd__o22a_1 _23605_ (.A1(_07569_),
    .A2(_07570_),
    .B1(_07444_),
    .B2(_07571_),
    .X(_07710_));
 sky130_fd_sc_hd__a2bb2o_1 _23606_ (.A1_N(_07709_),
    .A2_N(_07710_),
    .B1(_07709_),
    .B2(_07710_),
    .X(_07711_));
 sky130_fd_sc_hd__a2bb2o_1 _23607_ (.A1_N(_07443_),
    .A2_N(_07711_),
    .B1(_07443_),
    .B2(_07711_),
    .X(_07712_));
 sky130_fd_sc_hd__o22a_1 _23608_ (.A1(_07572_),
    .A2(_07573_),
    .B1(_07313_),
    .B2(_07574_),
    .X(_07713_));
 sky130_fd_sc_hd__or2_1 _23609_ (.A(_07712_),
    .B(_07713_),
    .X(_07714_));
 sky130_fd_sc_hd__a21bo_1 _23610_ (.A1(_07712_),
    .A2(_07713_),
    .B1_N(_07714_),
    .X(_07715_));
 sky130_fd_sc_hd__buf_1 _23611_ (.A(_07715_),
    .X(_07716_));
 sky130_fd_sc_hd__or2_1 _23612_ (.A(_07437_),
    .B(_07578_),
    .X(_07717_));
 sky130_fd_sc_hd__or3_1 _23613_ (.A(_07152_),
    .B(_07309_),
    .C(_07717_),
    .X(_07718_));
 sky130_fd_sc_hd__o221a_1 _23614_ (.A1(_07436_),
    .A2(_07576_),
    .B1(_07438_),
    .B2(_07717_),
    .C1(_07577_),
    .X(_07719_));
 sky130_fd_sc_hd__o21ai_1 _23615_ (.A1(_07160_),
    .A2(_07718_),
    .B1(_07719_),
    .Y(_07720_));
 sky130_vsdinv _23616_ (.A(_07720_),
    .Y(_07721_));
 sky130_vsdinv _23617_ (.A(_07716_),
    .Y(_07722_));
 sky130_fd_sc_hd__o22a_1 _23618_ (.A1(_07716_),
    .A2(_07721_),
    .B1(_07722_),
    .B2(_07720_),
    .X(_02647_));
 sky130_fd_sc_hd__o22a_1 _23619_ (.A1(_07709_),
    .A2(_07710_),
    .B1(_07443_),
    .B2(_07711_),
    .X(_07723_));
 sky130_fd_sc_hd__o22a_1 _23620_ (.A1(_07585_),
    .A2(_07625_),
    .B1(_07584_),
    .B2(_07626_),
    .X(_07724_));
 sky130_fd_sc_hd__o22a_1 _23621_ (.A1(_07605_),
    .A2(_07606_),
    .B1(_07586_),
    .B2(_07607_),
    .X(_07725_));
 sky130_fd_sc_hd__or2_1 _23622_ (.A(_07724_),
    .B(_07725_),
    .X(_07726_));
 sky130_fd_sc_hd__a21bo_1 _23623_ (.A1(_07724_),
    .A2(_07725_),
    .B1_N(_07726_),
    .X(_07727_));
 sky130_fd_sc_hd__o22a_1 _23624_ (.A1(_07622_),
    .A2(_07623_),
    .B1(_07608_),
    .B2(_07624_),
    .X(_07728_));
 sky130_fd_sc_hd__o22a_2 _23625_ (.A1(_07629_),
    .A2(_07654_),
    .B1(_07628_),
    .B2(_07655_),
    .X(_07729_));
 sky130_fd_sc_hd__o21ba_1 _23626_ (.A1(_07591_),
    .A2(_07592_),
    .B1_N(_07589_),
    .X(_07730_));
 sky130_fd_sc_hd__and4_1 _23627_ (.A(_05823_),
    .B(_07588_),
    .C(_05824_),
    .D(_13520_),
    .X(_07731_));
 sky130_fd_sc_hd__buf_1 _23628_ (.A(_07462_),
    .X(_07732_));
 sky130_fd_sc_hd__clkbuf_2 _23629_ (.A(_07732_),
    .X(_07733_));
 sky130_fd_sc_hd__o22a_1 _23630_ (.A1(_05816_),
    .A2(_07733_),
    .B1(_06753_),
    .B2(_07596_),
    .X(_07734_));
 sky130_fd_sc_hd__or2_1 _23631_ (.A(_07731_),
    .B(_07734_),
    .X(_07735_));
 sky130_fd_sc_hd__buf_1 _23632_ (.A(_07325_),
    .X(_07736_));
 sky130_fd_sc_hd__buf_2 _23633_ (.A(_07736_),
    .X(_07737_));
 sky130_fd_sc_hd__or2_1 _23634_ (.A(_07456_),
    .B(_07737_),
    .X(_07738_));
 sky130_fd_sc_hd__a2bb2o_1 _23635_ (.A1_N(_07735_),
    .A2_N(_07738_),
    .B1(_07735_),
    .B2(_07738_),
    .X(_07739_));
 sky130_fd_sc_hd__buf_1 _23636_ (.A(_13538_),
    .X(_07740_));
 sky130_fd_sc_hd__buf_1 _23637_ (.A(\pcpi_mul.rs1[25] ),
    .X(_07741_));
 sky130_fd_sc_hd__buf_1 _23638_ (.A(_07741_),
    .X(_07742_));
 sky130_fd_sc_hd__and4_1 _23639_ (.A(_06459_),
    .B(_07740_),
    .C(_06461_),
    .D(_07742_),
    .X(_07743_));
 sky130_fd_sc_hd__clkbuf_2 _23640_ (.A(_07031_),
    .X(_07744_));
 sky130_fd_sc_hd__o22a_1 _23641_ (.A1(_06578_),
    .A2(_07744_),
    .B1(_06579_),
    .B2(_07452_),
    .X(_07745_));
 sky130_fd_sc_hd__or2_1 _23642_ (.A(_07743_),
    .B(_07745_),
    .X(_07746_));
 sky130_vsdinv _23643_ (.A(\pcpi_mul.rs1[29] ),
    .Y(_07747_));
 sky130_fd_sc_hd__buf_1 _23644_ (.A(_07747_),
    .X(_07748_));
 sky130_fd_sc_hd__buf_2 _23645_ (.A(_07748_),
    .X(_07749_));
 sky130_fd_sc_hd__or2_1 _23646_ (.A(_07030_),
    .B(_07749_),
    .X(_07750_));
 sky130_fd_sc_hd__a2bb2o_1 _23647_ (.A1_N(_07746_),
    .A2_N(_07750_),
    .B1(_07746_),
    .B2(_07750_),
    .X(_07751_));
 sky130_fd_sc_hd__o21ba_1 _23648_ (.A1(_07597_),
    .A2(_07601_),
    .B1_N(_07599_),
    .X(_07752_));
 sky130_fd_sc_hd__a2bb2o_1 _23649_ (.A1_N(_07751_),
    .A2_N(_07752_),
    .B1(_07751_),
    .B2(_07752_),
    .X(_07753_));
 sky130_fd_sc_hd__a2bb2o_1 _23650_ (.A1_N(_07739_),
    .A2_N(_07753_),
    .B1(_07739_),
    .B2(_07753_),
    .X(_07754_));
 sky130_fd_sc_hd__o22a_1 _23651_ (.A1(_07602_),
    .A2(_07603_),
    .B1(_07593_),
    .B2(_07604_),
    .X(_07755_));
 sky130_fd_sc_hd__a2bb2o_1 _23652_ (.A1_N(_07754_),
    .A2_N(_07755_),
    .B1(_07754_),
    .B2(_07755_),
    .X(_07756_));
 sky130_fd_sc_hd__a2bb2o_1 _23653_ (.A1_N(_07730_),
    .A2_N(_07756_),
    .B1(_07730_),
    .B2(_07756_),
    .X(_07757_));
 sky130_fd_sc_hd__o22a_1 _23654_ (.A1(_07612_),
    .A2(_07618_),
    .B1(_07611_),
    .B2(_07619_),
    .X(_07758_));
 sky130_fd_sc_hd__o22a_1 _23655_ (.A1(_07639_),
    .A2(_07640_),
    .B1(_07634_),
    .B2(_07641_),
    .X(_07759_));
 sky130_fd_sc_hd__o21ba_1 _23656_ (.A1(_07614_),
    .A2(_07617_),
    .B1_N(_07615_),
    .X(_07760_));
 sky130_fd_sc_hd__o21ba_1 _23657_ (.A1(_07630_),
    .A2(_07633_),
    .B1_N(_07632_),
    .X(_07761_));
 sky130_fd_sc_hd__clkbuf_2 _23658_ (.A(_06648_),
    .X(_07762_));
 sky130_fd_sc_hd__o22a_1 _23659_ (.A1(_06919_),
    .A2(_07762_),
    .B1(_06920_),
    .B2(_06762_),
    .X(_07763_));
 sky130_fd_sc_hd__buf_1 _23660_ (.A(_13545_),
    .X(_07764_));
 sky130_fd_sc_hd__and4_1 _23661_ (.A(_06923_),
    .B(_07191_),
    .C(_06924_),
    .D(_07764_),
    .X(_07765_));
 sky130_fd_sc_hd__nor2_2 _23662_ (.A(_07763_),
    .B(_07765_),
    .Y(_07766_));
 sky130_fd_sc_hd__nor2_2 _23663_ (.A(_06915_),
    .B(_07019_),
    .Y(_07767_));
 sky130_fd_sc_hd__a2bb2o_1 _23664_ (.A1_N(_07766_),
    .A2_N(_07767_),
    .B1(_07766_),
    .B2(_07767_),
    .X(_07768_));
 sky130_fd_sc_hd__a2bb2o_1 _23665_ (.A1_N(_07761_),
    .A2_N(_07768_),
    .B1(_07761_),
    .B2(_07768_),
    .X(_07769_));
 sky130_fd_sc_hd__a2bb2o_1 _23666_ (.A1_N(_07760_),
    .A2_N(_07769_),
    .B1(_07760_),
    .B2(_07769_),
    .X(_07770_));
 sky130_fd_sc_hd__a2bb2o_1 _23667_ (.A1_N(_07759_),
    .A2_N(_07770_),
    .B1(_07759_),
    .B2(_07770_),
    .X(_07771_));
 sky130_fd_sc_hd__a2bb2o_1 _23668_ (.A1_N(_07758_),
    .A2_N(_07771_),
    .B1(_07758_),
    .B2(_07771_),
    .X(_07772_));
 sky130_fd_sc_hd__o22a_1 _23669_ (.A1(_07610_),
    .A2(_07620_),
    .B1(_07609_),
    .B2(_07621_),
    .X(_07773_));
 sky130_fd_sc_hd__a2bb2o_1 _23670_ (.A1_N(_07772_),
    .A2_N(_07773_),
    .B1(_07772_),
    .B2(_07773_),
    .X(_07774_));
 sky130_fd_sc_hd__a2bb2o_1 _23671_ (.A1_N(_07757_),
    .A2_N(_07774_),
    .B1(_07757_),
    .B2(_07774_),
    .X(_07775_));
 sky130_fd_sc_hd__a2bb2o_1 _23672_ (.A1_N(_07729_),
    .A2_N(_07775_),
    .B1(_07729_),
    .B2(_07775_),
    .X(_07776_));
 sky130_fd_sc_hd__a2bb2o_1 _23673_ (.A1_N(_07728_),
    .A2_N(_07776_),
    .B1(_07728_),
    .B2(_07776_),
    .X(_07777_));
 sky130_fd_sc_hd__o22a_1 _23674_ (.A1(_07651_),
    .A2(_07652_),
    .B1(_07642_),
    .B2(_07653_),
    .X(_07778_));
 sky130_fd_sc_hd__o22a_1 _23675_ (.A1(_07541_),
    .A2(_07674_),
    .B1(_07657_),
    .B2(_07675_),
    .X(_07779_));
 sky130_fd_sc_hd__clkbuf_2 _23676_ (.A(_06574_),
    .X(_07780_));
 sky130_fd_sc_hd__or2_1 _23677_ (.A(_06519_),
    .B(_07780_),
    .X(_07781_));
 sky130_fd_sc_hd__o22a_1 _23678_ (.A1(_06522_),
    .A2(_06765_),
    .B1(_07108_),
    .B2(_06565_),
    .X(_07782_));
 sky130_fd_sc_hd__and4_1 _23679_ (.A(_06525_),
    .B(_06898_),
    .C(_06527_),
    .D(_07484_),
    .X(_07783_));
 sky130_fd_sc_hd__or2_1 _23680_ (.A(_07782_),
    .B(_07783_),
    .X(_07784_));
 sky130_fd_sc_hd__a2bb2o_1 _23681_ (.A1_N(_07781_),
    .A2_N(_07784_),
    .B1(_07781_),
    .B2(_07784_),
    .X(_07785_));
 sky130_fd_sc_hd__or2_1 _23682_ (.A(_05791_),
    .B(_06227_),
    .X(_07786_));
 sky130_fd_sc_hd__o22a_1 _23683_ (.A1(_07237_),
    .A2(_06456_),
    .B1(_06970_),
    .B2(_06580_),
    .X(_07787_));
 sky130_fd_sc_hd__and4_1 _23684_ (.A(_07115_),
    .B(_06462_),
    .C(_07116_),
    .D(_06583_),
    .X(_07788_));
 sky130_fd_sc_hd__or2_1 _23685_ (.A(_07787_),
    .B(_07788_),
    .X(_07789_));
 sky130_fd_sc_hd__a2bb2o_1 _23686_ (.A1_N(_07786_),
    .A2_N(_07789_),
    .B1(_07786_),
    .B2(_07789_),
    .X(_07790_));
 sky130_fd_sc_hd__o21ba_1 _23687_ (.A1(_07635_),
    .A2(_07638_),
    .B1_N(_07636_),
    .X(_07791_));
 sky130_fd_sc_hd__a2bb2o_1 _23688_ (.A1_N(_07790_),
    .A2_N(_07791_),
    .B1(_07790_),
    .B2(_07791_),
    .X(_07792_));
 sky130_fd_sc_hd__a2bb2o_2 _23689_ (.A1_N(_07785_),
    .A2_N(_07792_),
    .B1(_07785_),
    .B2(_07792_),
    .X(_07793_));
 sky130_fd_sc_hd__o21ba_1 _23690_ (.A1(_07645_),
    .A2(_07648_),
    .B1_N(_07646_),
    .X(_07794_));
 sky130_fd_sc_hd__o21ba_1 _23691_ (.A1(_07658_),
    .A2(_07661_),
    .B1_N(_07660_),
    .X(_07795_));
 sky130_fd_sc_hd__or2_2 _23692_ (.A(_06096_),
    .B(_06599_),
    .X(_07796_));
 sky130_fd_sc_hd__o22a_1 _23693_ (.A1(_07383_),
    .A2(_05735_),
    .B1(_07254_),
    .B2(_06231_),
    .X(_07797_));
 sky130_fd_sc_hd__buf_2 _23694_ (.A(_06722_),
    .X(_07798_));
 sky130_fd_sc_hd__buf_2 _23695_ (.A(_06723_),
    .X(_07799_));
 sky130_fd_sc_hd__and4_1 _23696_ (.A(_07798_),
    .B(_06234_),
    .C(_07799_),
    .D(_06236_),
    .X(_07800_));
 sky130_fd_sc_hd__or2_1 _23697_ (.A(_07797_),
    .B(_07800_),
    .X(_07801_));
 sky130_fd_sc_hd__a2bb2o_1 _23698_ (.A1_N(_07796_),
    .A2_N(_07801_),
    .B1(_07796_),
    .B2(_07801_),
    .X(_07802_));
 sky130_fd_sc_hd__a2bb2o_1 _23699_ (.A1_N(_07795_),
    .A2_N(_07802_),
    .B1(_07795_),
    .B2(_07802_),
    .X(_07803_));
 sky130_fd_sc_hd__a2bb2o_1 _23700_ (.A1_N(_07794_),
    .A2_N(_07803_),
    .B1(_07794_),
    .B2(_07803_),
    .X(_07804_));
 sky130_fd_sc_hd__o22a_1 _23701_ (.A1(_07644_),
    .A2(_07649_),
    .B1(_07643_),
    .B2(_07650_),
    .X(_07805_));
 sky130_fd_sc_hd__a2bb2o_1 _23702_ (.A1_N(_07804_),
    .A2_N(_07805_),
    .B1(_07804_),
    .B2(_07805_),
    .X(_07806_));
 sky130_fd_sc_hd__a2bb2o_1 _23703_ (.A1_N(_07793_),
    .A2_N(_07806_),
    .B1(_07793_),
    .B2(_07806_),
    .X(_07807_));
 sky130_fd_sc_hd__a2bb2o_1 _23704_ (.A1_N(_07779_),
    .A2_N(_07807_),
    .B1(_07779_),
    .B2(_07807_),
    .X(_07808_));
 sky130_fd_sc_hd__a2bb2o_1 _23705_ (.A1_N(_07778_),
    .A2_N(_07808_),
    .B1(_07778_),
    .B2(_07808_),
    .X(_07809_));
 sky130_fd_sc_hd__o22a_1 _23706_ (.A1(_07671_),
    .A2(_07672_),
    .B1(_07662_),
    .B2(_07673_),
    .X(_07810_));
 sky130_fd_sc_hd__or2_1 _23707_ (.A(_07546_),
    .B(_06520_),
    .X(_07811_));
 sky130_fd_sc_hd__clkbuf_2 _23708_ (.A(_06810_),
    .X(_07812_));
 sky130_fd_sc_hd__o22a_1 _23709_ (.A1(_07812_),
    .A2(_05843_),
    .B1(_06395_),
    .B2(_05830_),
    .X(_07813_));
 sky130_fd_sc_hd__and4_1 _23710_ (.A(_07549_),
    .B(_06526_),
    .C(_07406_),
    .D(_06528_),
    .X(_07814_));
 sky130_fd_sc_hd__or2_1 _23711_ (.A(_07813_),
    .B(_07814_),
    .X(_07815_));
 sky130_fd_sc_hd__a2bb2o_1 _23712_ (.A1_N(_07811_),
    .A2_N(_07815_),
    .B1(_07811_),
    .B2(_07815_),
    .X(_07816_));
 sky130_fd_sc_hd__or2_1 _23713_ (.A(_06803_),
    .B(_07403_),
    .X(_07817_));
 sky130_fd_sc_hd__clkbuf_2 _23714_ (.A(_06805_),
    .X(_07818_));
 sky130_fd_sc_hd__o22a_1 _23715_ (.A1(_07665_),
    .A2(_06003_),
    .B1(_07818_),
    .B2(_06099_),
    .X(_07819_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _23716_ (.A(_05741_),
    .X(_07820_));
 sky130_fd_sc_hd__and4_1 _23717_ (.A(_07667_),
    .B(_07405_),
    .C(_07668_),
    .D(_07820_),
    .X(_07821_));
 sky130_fd_sc_hd__or2_1 _23718_ (.A(_07819_),
    .B(_07821_),
    .X(_07822_));
 sky130_fd_sc_hd__a2bb2o_1 _23719_ (.A1_N(_07817_),
    .A2_N(_07822_),
    .B1(_07817_),
    .B2(_07822_),
    .X(_07823_));
 sky130_fd_sc_hd__o21ba_1 _23720_ (.A1(_07664_),
    .A2(_07670_),
    .B1_N(_07669_),
    .X(_07824_));
 sky130_fd_sc_hd__a2bb2o_1 _23721_ (.A1_N(_07823_),
    .A2_N(_07824_),
    .B1(_07823_),
    .B2(_07824_),
    .X(_07825_));
 sky130_fd_sc_hd__a2bb2o_1 _23722_ (.A1_N(_07816_),
    .A2_N(_07825_),
    .B1(_07816_),
    .B2(_07825_),
    .X(_07826_));
 sky130_fd_sc_hd__a2bb2o_1 _23723_ (.A1_N(_07696_),
    .A2_N(_07826_),
    .B1(_07696_),
    .B2(_07826_),
    .X(_07827_));
 sky130_fd_sc_hd__a2bb2o_1 _23724_ (.A1_N(_07810_),
    .A2_N(_07827_),
    .B1(_07810_),
    .B2(_07827_),
    .X(_07828_));
 sky130_fd_sc_hd__or2_1 _23725_ (.A(_07529_),
    .B(_05316_),
    .X(_07829_));
 sky130_fd_sc_hd__buf_1 _23726_ (.A(\pcpi_mul.rs2[28] ),
    .X(_07830_));
 sky130_fd_sc_hd__and4_1 _23727_ (.A(_07830_),
    .B(_05915_),
    .C(\pcpi_mul.rs2[29] ),
    .D(_13626_),
    .X(_07831_));
 sky130_vsdinv _23728_ (.A(\pcpi_mul.rs2[29] ),
    .Y(_07832_));
 sky130_fd_sc_hd__o22a_1 _23729_ (.A1(_07677_),
    .A2(_05910_),
    .B1(_07832_),
    .B2(_05324_),
    .X(_07833_));
 sky130_fd_sc_hd__or2_1 _23730_ (.A(_07831_),
    .B(_07833_),
    .X(_07834_));
 sky130_fd_sc_hd__a2bb2o_1 _23731_ (.A1_N(_07829_),
    .A2_N(_07834_),
    .B1(_07829_),
    .B2(_07834_),
    .X(_07835_));
 sky130_fd_sc_hd__o21ba_1 _23732_ (.A1(_07689_),
    .A2(_07694_),
    .B1_N(_07693_),
    .X(_07836_));
 sky130_fd_sc_hd__or2_1 _23733_ (.A(_07688_),
    .B(_05900_),
    .X(_07837_));
 sky130_fd_sc_hd__o22a_1 _23734_ (.A1(_07690_),
    .A2(_06112_),
    .B1(_07691_),
    .B2(_06939_),
    .X(_07838_));
 sky130_fd_sc_hd__and4_1 _23735_ (.A(_07536_),
    .B(_06116_),
    .C(_13091_),
    .D(_07085_),
    .X(_07839_));
 sky130_fd_sc_hd__or2_1 _23736_ (.A(_07838_),
    .B(_07839_),
    .X(_07840_));
 sky130_fd_sc_hd__a2bb2o_1 _23737_ (.A1_N(_07837_),
    .A2_N(_07840_),
    .B1(_07837_),
    .B2(_07840_),
    .X(_07841_));
 sky130_fd_sc_hd__a2bb2o_1 _23738_ (.A1_N(_07685_),
    .A2_N(_07841_),
    .B1(_07685_),
    .B2(_07841_),
    .X(_07842_));
 sky130_fd_sc_hd__a2bb2o_1 _23739_ (.A1_N(_07836_),
    .A2_N(_07842_),
    .B1(_07836_),
    .B2(_07842_),
    .X(_07843_));
 sky130_fd_sc_hd__or2_1 _23740_ (.A(_07835_),
    .B(_07843_),
    .X(_07844_));
 sky130_fd_sc_hd__a21bo_1 _23741_ (.A1(_07835_),
    .A2(_07843_),
    .B1_N(_07844_),
    .X(_07845_));
 sky130_fd_sc_hd__a2bb2o_1 _23742_ (.A1_N(_07698_),
    .A2_N(_07845_),
    .B1(_07698_),
    .B2(_07845_),
    .X(_07846_));
 sky130_fd_sc_hd__a2bb2o_1 _23743_ (.A1_N(_07828_),
    .A2_N(_07846_),
    .B1(_07828_),
    .B2(_07846_),
    .X(_07847_));
 sky130_fd_sc_hd__o22a_1 _23744_ (.A1(_07543_),
    .A2(_07699_),
    .B1(_07676_),
    .B2(_07700_),
    .X(_07848_));
 sky130_fd_sc_hd__a2bb2o_1 _23745_ (.A1_N(_07847_),
    .A2_N(_07848_),
    .B1(_07847_),
    .B2(_07848_),
    .X(_07849_));
 sky130_fd_sc_hd__a2bb2o_2 _23746_ (.A1_N(_07809_),
    .A2_N(_07849_),
    .B1(_07809_),
    .B2(_07849_),
    .X(_07850_));
 sky130_fd_sc_hd__o22a_2 _23747_ (.A1(_07563_),
    .A2(_07701_),
    .B1(_07656_),
    .B2(_07702_),
    .X(_07851_));
 sky130_fd_sc_hd__a2bb2o_1 _23748_ (.A1_N(_07850_),
    .A2_N(_07851_),
    .B1(_07850_),
    .B2(_07851_),
    .X(_07852_));
 sky130_fd_sc_hd__a2bb2o_1 _23749_ (.A1_N(_07777_),
    .A2_N(_07852_),
    .B1(_07777_),
    .B2(_07852_),
    .X(_07853_));
 sky130_fd_sc_hd__o22a_1 _23750_ (.A1(_07703_),
    .A2(_07704_),
    .B1(_07627_),
    .B2(_07705_),
    .X(_07854_));
 sky130_fd_sc_hd__a2bb2o_1 _23751_ (.A1_N(_07853_),
    .A2_N(_07854_),
    .B1(_07853_),
    .B2(_07854_),
    .X(_07855_));
 sky130_fd_sc_hd__a2bb2o_1 _23752_ (.A1_N(_07727_),
    .A2_N(_07855_),
    .B1(_07727_),
    .B2(_07855_),
    .X(_07856_));
 sky130_fd_sc_hd__o22a_1 _23753_ (.A1(_07706_),
    .A2(_07707_),
    .B1(_07583_),
    .B2(_07708_),
    .X(_07857_));
 sky130_fd_sc_hd__a2bb2o_1 _23754_ (.A1_N(_07856_),
    .A2_N(_07857_),
    .B1(_07856_),
    .B2(_07857_),
    .X(_07858_));
 sky130_fd_sc_hd__a2bb2o_1 _23755_ (.A1_N(_07582_),
    .A2_N(_07858_),
    .B1(_07582_),
    .B2(_07858_),
    .X(_07859_));
 sky130_fd_sc_hd__or2_1 _23756_ (.A(_07723_),
    .B(_07859_),
    .X(_07860_));
 sky130_fd_sc_hd__a21bo_1 _23757_ (.A1(_07723_),
    .A2(_07859_),
    .B1_N(_07860_),
    .X(_07861_));
 sky130_fd_sc_hd__o21ai_1 _23758_ (.A1(_07716_),
    .A2(_07721_),
    .B1(_07714_),
    .Y(_07862_));
 sky130_fd_sc_hd__a2bb2o_1 _23759_ (.A1_N(_07861_),
    .A2_N(_07862_),
    .B1(_07861_),
    .B2(_07862_),
    .X(_02648_));
 sky130_fd_sc_hd__o22a_1 _23760_ (.A1(_07729_),
    .A2(_07775_),
    .B1(_07728_),
    .B2(_07776_),
    .X(_07863_));
 sky130_fd_sc_hd__o22a_1 _23761_ (.A1(_07754_),
    .A2(_07755_),
    .B1(_07730_),
    .B2(_07756_),
    .X(_07864_));
 sky130_fd_sc_hd__or2_2 _23762_ (.A(_07863_),
    .B(_07864_),
    .X(_07865_));
 sky130_fd_sc_hd__a21bo_1 _23763_ (.A1(_07863_),
    .A2(_07864_),
    .B1_N(_07865_),
    .X(_07866_));
 sky130_fd_sc_hd__o22a_4 _23764_ (.A1(_07772_),
    .A2(_07773_),
    .B1(_07757_),
    .B2(_07774_),
    .X(_07867_));
 sky130_fd_sc_hd__o22a_1 _23765_ (.A1(_07779_),
    .A2(_07807_),
    .B1(_07778_),
    .B2(_07808_),
    .X(_07868_));
 sky130_fd_sc_hd__o21ba_1 _23766_ (.A1(_07735_),
    .A2(_07738_),
    .B1_N(_07731_),
    .X(_07869_));
 sky130_fd_sc_hd__buf_1 _23767_ (.A(_07594_),
    .X(_07870_));
 sky130_fd_sc_hd__clkbuf_4 _23768_ (.A(_07870_),
    .X(_07871_));
 sky130_fd_sc_hd__buf_1 _23769_ (.A(_07747_),
    .X(_07872_));
 sky130_fd_sc_hd__buf_1 _23770_ (.A(_07872_),
    .X(_07873_));
 sky130_fd_sc_hd__buf_2 _23771_ (.A(_07873_),
    .X(_07874_));
 sky130_fd_sc_hd__o22a_1 _23772_ (.A1(_06433_),
    .A2(_07871_),
    .B1(_06436_),
    .B2(_07874_),
    .X(_07875_));
 sky130_fd_sc_hd__buf_1 _23773_ (.A(\pcpi_mul.rs1[28] ),
    .X(_07876_));
 sky130_fd_sc_hd__buf_1 _23774_ (.A(_07876_),
    .X(_07877_));
 sky130_fd_sc_hd__buf_1 _23775_ (.A(_07877_),
    .X(_07878_));
 sky130_fd_sc_hd__and4_1 _23776_ (.A(_07022_),
    .B(_07878_),
    .C(_07023_),
    .D(_13516_),
    .X(_07879_));
 sky130_fd_sc_hd__nor2_1 _23777_ (.A(_07875_),
    .B(_07879_),
    .Y(_07880_));
 sky130_fd_sc_hd__buf_2 _23778_ (.A(_07733_),
    .X(_07881_));
 sky130_fd_sc_hd__nor2_2 _23779_ (.A(_07027_),
    .B(_07881_),
    .Y(_07882_));
 sky130_fd_sc_hd__a2bb2o_1 _23780_ (.A1_N(_07880_),
    .A2_N(_07882_),
    .B1(_07880_),
    .B2(_07882_),
    .X(_07883_));
 sky130_fd_sc_hd__buf_2 _23781_ (.A(_07325_),
    .X(_07884_));
 sky130_fd_sc_hd__o22a_1 _23782_ (.A1(_06894_),
    .A2(_07197_),
    .B1(_06895_),
    .B2(_07884_),
    .X(_07885_));
 sky130_fd_sc_hd__buf_1 _23783_ (.A(_07741_),
    .X(_07886_));
 sky130_fd_sc_hd__and4_1 _23784_ (.A(_07186_),
    .B(_07886_),
    .C(_07189_),
    .D(_07449_),
    .X(_07887_));
 sky130_fd_sc_hd__nor2_2 _23785_ (.A(_07885_),
    .B(_07887_),
    .Y(_07888_));
 sky130_vsdinv _23786_ (.A(\pcpi_mul.rs1[30] ),
    .Y(_07889_));
 sky130_fd_sc_hd__buf_1 _23787_ (.A(_07889_),
    .X(_07890_));
 sky130_fd_sc_hd__buf_1 _23788_ (.A(_07890_),
    .X(_07891_));
 sky130_fd_sc_hd__buf_2 _23789_ (.A(_07891_),
    .X(_07892_));
 sky130_fd_sc_hd__nor2_2 _23790_ (.A(_05311_),
    .B(_07892_),
    .Y(_07893_));
 sky130_fd_sc_hd__a2bb2o_1 _23791_ (.A1_N(_07888_),
    .A2_N(_07893_),
    .B1(_07888_),
    .B2(_07893_),
    .X(_07894_));
 sky130_fd_sc_hd__o21ba_1 _23792_ (.A1(_07746_),
    .A2(_07750_),
    .B1_N(_07743_),
    .X(_07895_));
 sky130_fd_sc_hd__a2bb2o_1 _23793_ (.A1_N(_07894_),
    .A2_N(_07895_),
    .B1(_07894_),
    .B2(_07895_),
    .X(_07896_));
 sky130_fd_sc_hd__a2bb2o_1 _23794_ (.A1_N(_07883_),
    .A2_N(_07896_),
    .B1(_07883_),
    .B2(_07896_),
    .X(_07897_));
 sky130_fd_sc_hd__o22a_1 _23795_ (.A1(_07751_),
    .A2(_07752_),
    .B1(_07739_),
    .B2(_07753_),
    .X(_07898_));
 sky130_fd_sc_hd__a2bb2o_1 _23796_ (.A1_N(_07897_),
    .A2_N(_07898_),
    .B1(_07897_),
    .B2(_07898_),
    .X(_07899_));
 sky130_fd_sc_hd__a2bb2o_1 _23797_ (.A1_N(_07869_),
    .A2_N(_07899_),
    .B1(_07869_),
    .B2(_07899_),
    .X(_07900_));
 sky130_fd_sc_hd__o22a_1 _23798_ (.A1(_07761_),
    .A2(_07768_),
    .B1(_07760_),
    .B2(_07769_),
    .X(_07901_));
 sky130_fd_sc_hd__o22a_1 _23799_ (.A1(_07790_),
    .A2(_07791_),
    .B1(_07785_),
    .B2(_07792_),
    .X(_07902_));
 sky130_fd_sc_hd__a21oi_2 _23800_ (.A1(_07766_),
    .A2(_07767_),
    .B1(_07765_),
    .Y(_07903_));
 sky130_fd_sc_hd__o21ba_1 _23801_ (.A1(_07781_),
    .A2(_07784_),
    .B1_N(_07783_),
    .X(_07904_));
 sky130_fd_sc_hd__buf_1 _23802_ (.A(_06761_),
    .X(_07905_));
 sky130_fd_sc_hd__o22a_1 _23803_ (.A1(_06919_),
    .A2(_07905_),
    .B1(_06920_),
    .B2(_06891_),
    .X(_07906_));
 sky130_fd_sc_hd__buf_1 _23804_ (.A(\pcpi_mul.rs1[22] ),
    .X(_07907_));
 sky130_fd_sc_hd__buf_1 _23805_ (.A(\pcpi_mul.rs1[23] ),
    .X(_07908_));
 sky130_fd_sc_hd__and4_1 _23806_ (.A(_06923_),
    .B(_07907_),
    .C(_06924_),
    .D(_07908_),
    .X(_07909_));
 sky130_fd_sc_hd__nor2_2 _23807_ (.A(_07906_),
    .B(_07909_),
    .Y(_07910_));
 sky130_fd_sc_hd__nor2_2 _23808_ (.A(_06915_),
    .B(_07458_),
    .Y(_07911_));
 sky130_fd_sc_hd__a2bb2o_1 _23809_ (.A1_N(_07910_),
    .A2_N(_07911_),
    .B1(_07910_),
    .B2(_07911_),
    .X(_07912_));
 sky130_fd_sc_hd__a2bb2o_1 _23810_ (.A1_N(_07904_),
    .A2_N(_07912_),
    .B1(_07904_),
    .B2(_07912_),
    .X(_07913_));
 sky130_fd_sc_hd__a2bb2o_1 _23811_ (.A1_N(_07903_),
    .A2_N(_07913_),
    .B1(_07903_),
    .B2(_07913_),
    .X(_07914_));
 sky130_fd_sc_hd__a2bb2o_1 _23812_ (.A1_N(_07902_),
    .A2_N(_07914_),
    .B1(_07902_),
    .B2(_07914_),
    .X(_07915_));
 sky130_fd_sc_hd__a2bb2o_1 _23813_ (.A1_N(_07901_),
    .A2_N(_07915_),
    .B1(_07901_),
    .B2(_07915_),
    .X(_07916_));
 sky130_fd_sc_hd__o22a_1 _23814_ (.A1(_07759_),
    .A2(_07770_),
    .B1(_07758_),
    .B2(_07771_),
    .X(_07917_));
 sky130_fd_sc_hd__a2bb2o_1 _23815_ (.A1_N(_07916_),
    .A2_N(_07917_),
    .B1(_07916_),
    .B2(_07917_),
    .X(_07918_));
 sky130_fd_sc_hd__a2bb2o_2 _23816_ (.A1_N(_07900_),
    .A2_N(_07918_),
    .B1(_07900_),
    .B2(_07918_),
    .X(_07919_));
 sky130_fd_sc_hd__a2bb2o_1 _23817_ (.A1_N(_07868_),
    .A2_N(_07919_),
    .B1(_07868_),
    .B2(_07919_),
    .X(_07920_));
 sky130_fd_sc_hd__a2bb2o_2 _23818_ (.A1_N(_07867_),
    .A2_N(_07920_),
    .B1(_07867_),
    .B2(_07920_),
    .X(_07921_));
 sky130_fd_sc_hd__o22a_1 _23819_ (.A1(_07804_),
    .A2(_07805_),
    .B1(_07793_),
    .B2(_07806_),
    .X(_07922_));
 sky130_fd_sc_hd__o22a_1 _23820_ (.A1(_07696_),
    .A2(_07826_),
    .B1(_07810_),
    .B2(_07827_),
    .X(_07923_));
 sky130_fd_sc_hd__or2_1 _23821_ (.A(_06820_),
    .B(_06754_),
    .X(_07924_));
 sky130_fd_sc_hd__o22a_1 _23822_ (.A1(_06822_),
    .A2(_06450_),
    .B1(_06960_),
    .B2(_06640_),
    .X(_07925_));
 sky130_fd_sc_hd__and4_1 _23823_ (.A(_06824_),
    .B(_13555_),
    .C(_06825_),
    .D(_07039_),
    .X(_07926_));
 sky130_fd_sc_hd__or2_1 _23824_ (.A(_07925_),
    .B(_07926_),
    .X(_07927_));
 sky130_fd_sc_hd__a2bb2o_1 _23825_ (.A1_N(_07924_),
    .A2_N(_07927_),
    .B1(_07924_),
    .B2(_07927_),
    .X(_07928_));
 sky130_fd_sc_hd__or2_1 _23826_ (.A(_07369_),
    .B(_06766_),
    .X(_07929_));
 sky130_fd_sc_hd__clkbuf_2 _23827_ (.A(_06111_),
    .X(_07930_));
 sky130_fd_sc_hd__o22a_1 _23828_ (.A1(_06969_),
    .A2(_06580_),
    .B1(_07930_),
    .B2(_06226_),
    .X(_07931_));
 sky130_fd_sc_hd__and4_1 _23829_ (.A(_06972_),
    .B(_06583_),
    .C(_06973_),
    .D(_07501_),
    .X(_07932_));
 sky130_fd_sc_hd__or2_1 _23830_ (.A(_07931_),
    .B(_07932_),
    .X(_07933_));
 sky130_fd_sc_hd__a2bb2o_1 _23831_ (.A1_N(_07929_),
    .A2_N(_07933_),
    .B1(_07929_),
    .B2(_07933_),
    .X(_07934_));
 sky130_fd_sc_hd__o21ba_1 _23832_ (.A1(_07786_),
    .A2(_07789_),
    .B1_N(_07788_),
    .X(_07935_));
 sky130_fd_sc_hd__a2bb2o_1 _23833_ (.A1_N(_07934_),
    .A2_N(_07935_),
    .B1(_07934_),
    .B2(_07935_),
    .X(_07936_));
 sky130_fd_sc_hd__a2bb2o_2 _23834_ (.A1_N(_07928_),
    .A2_N(_07936_),
    .B1(_07928_),
    .B2(_07936_),
    .X(_07937_));
 sky130_fd_sc_hd__o21ba_1 _23835_ (.A1(_07796_),
    .A2(_07801_),
    .B1_N(_07800_),
    .X(_07938_));
 sky130_fd_sc_hd__o21ba_1 _23836_ (.A1(_07811_),
    .A2(_07815_),
    .B1_N(_07814_),
    .X(_07939_));
 sky130_fd_sc_hd__or2_1 _23837_ (.A(_07516_),
    .B(_06669_),
    .X(_07940_));
 sky130_fd_sc_hd__buf_2 _23838_ (.A(_07128_),
    .X(_07941_));
 sky130_fd_sc_hd__o22a_1 _23839_ (.A1(_07941_),
    .A2(_06478_),
    .B1(_06089_),
    .B2(_06031_),
    .X(_07942_));
 sky130_fd_sc_hd__and4_1 _23840_ (.A(_07248_),
    .B(_06603_),
    .C(_07250_),
    .D(_13575_),
    .X(_07943_));
 sky130_fd_sc_hd__or2_1 _23841_ (.A(_07942_),
    .B(_07943_),
    .X(_07944_));
 sky130_fd_sc_hd__a2bb2o_1 _23842_ (.A1_N(_07940_),
    .A2_N(_07944_),
    .B1(_07940_),
    .B2(_07944_),
    .X(_07945_));
 sky130_fd_sc_hd__a2bb2o_1 _23843_ (.A1_N(_07939_),
    .A2_N(_07945_),
    .B1(_07939_),
    .B2(_07945_),
    .X(_07946_));
 sky130_fd_sc_hd__a2bb2o_1 _23844_ (.A1_N(_07938_),
    .A2_N(_07946_),
    .B1(_07938_),
    .B2(_07946_),
    .X(_07947_));
 sky130_fd_sc_hd__o22a_1 _23845_ (.A1(_07795_),
    .A2(_07802_),
    .B1(_07794_),
    .B2(_07803_),
    .X(_07948_));
 sky130_fd_sc_hd__a2bb2o_1 _23846_ (.A1_N(_07947_),
    .A2_N(_07948_),
    .B1(_07947_),
    .B2(_07948_),
    .X(_07949_));
 sky130_fd_sc_hd__a2bb2o_1 _23847_ (.A1_N(_07937_),
    .A2_N(_07949_),
    .B1(_07937_),
    .B2(_07949_),
    .X(_07950_));
 sky130_fd_sc_hd__a2bb2o_1 _23848_ (.A1_N(_07923_),
    .A2_N(_07950_),
    .B1(_07923_),
    .B2(_07950_),
    .X(_07951_));
 sky130_fd_sc_hd__a2bb2o_1 _23849_ (.A1_N(_07922_),
    .A2_N(_07951_),
    .B1(_07922_),
    .B2(_07951_),
    .X(_07952_));
 sky130_fd_sc_hd__o22a_1 _23850_ (.A1(_07823_),
    .A2(_07824_),
    .B1(_07816_),
    .B2(_07825_),
    .X(_07953_));
 sky130_fd_sc_hd__o22a_1 _23851_ (.A1(_07685_),
    .A2(_07841_),
    .B1(_07836_),
    .B2(_07842_),
    .X(_07954_));
 sky130_fd_sc_hd__or2_1 _23852_ (.A(_07546_),
    .B(_06702_),
    .X(_07955_));
 sky130_fd_sc_hd__o22a_1 _23853_ (.A1(_07812_),
    .A2(_06042_),
    .B1(_06395_),
    .B2(_06704_),
    .X(_07956_));
 sky130_fd_sc_hd__and4_1 _23854_ (.A(_07549_),
    .B(_06528_),
    .C(_07406_),
    .D(_06144_),
    .X(_07957_));
 sky130_fd_sc_hd__or2_1 _23855_ (.A(_07956_),
    .B(_07957_),
    .X(_07958_));
 sky130_fd_sc_hd__a2bb2o_1 _23856_ (.A1_N(_07955_),
    .A2_N(_07958_),
    .B1(_07955_),
    .B2(_07958_),
    .X(_07959_));
 sky130_fd_sc_hd__or2_1 _23857_ (.A(_07663_),
    .B(_06298_),
    .X(_07960_));
 sky130_fd_sc_hd__o22a_1 _23858_ (.A1(_07665_),
    .A2(_07277_),
    .B1(_06801_),
    .B2(_06983_),
    .X(_07961_));
 sky130_fd_sc_hd__and4_1 _23859_ (.A(_07667_),
    .B(_07820_),
    .C(_07668_),
    .D(_07249_),
    .X(_07962_));
 sky130_fd_sc_hd__or2_1 _23860_ (.A(_07961_),
    .B(_07962_),
    .X(_07963_));
 sky130_fd_sc_hd__a2bb2o_1 _23861_ (.A1_N(_07960_),
    .A2_N(_07963_),
    .B1(_07960_),
    .B2(_07963_),
    .X(_07964_));
 sky130_fd_sc_hd__o21ba_1 _23862_ (.A1(_07817_),
    .A2(_07822_),
    .B1_N(_07821_),
    .X(_07965_));
 sky130_fd_sc_hd__a2bb2o_1 _23863_ (.A1_N(_07964_),
    .A2_N(_07965_),
    .B1(_07964_),
    .B2(_07965_),
    .X(_07966_));
 sky130_fd_sc_hd__a2bb2o_1 _23864_ (.A1_N(_07959_),
    .A2_N(_07966_),
    .B1(_07959_),
    .B2(_07966_),
    .X(_07967_));
 sky130_fd_sc_hd__a2bb2o_1 _23865_ (.A1_N(_07954_),
    .A2_N(_07967_),
    .B1(_07954_),
    .B2(_07967_),
    .X(_07968_));
 sky130_fd_sc_hd__a2bb2o_1 _23866_ (.A1_N(_07953_),
    .A2_N(_07968_),
    .B1(_07953_),
    .B2(_07968_),
    .X(_07969_));
 sky130_vsdinv _23867_ (.A(\pcpi_mul.rs2[30] ),
    .Y(_07970_));
 sky130_fd_sc_hd__clkbuf_2 _23868_ (.A(_07970_),
    .X(_07971_));
 sky130_fd_sc_hd__clkbuf_4 _23869_ (.A(_07971_),
    .X(_07972_));
 sky130_fd_sc_hd__or2_2 _23870_ (.A(_07972_),
    .B(_05150_),
    .X(_07973_));
 sky130_fd_sc_hd__or2_1 _23871_ (.A(_07529_),
    .B(_06011_),
    .X(_07974_));
 sky130_fd_sc_hd__and4_1 _23872_ (.A(\pcpi_mul.rs2[29] ),
    .B(_05915_),
    .C(_07830_),
    .D(_06115_),
    .X(_07975_));
 sky130_fd_sc_hd__o22a_1 _23873_ (.A1(_07832_),
    .A2(_05910_),
    .B1(_07677_),
    .B2(_06015_),
    .X(_07976_));
 sky130_fd_sc_hd__or2_1 _23874_ (.A(_07975_),
    .B(_07976_),
    .X(_07977_));
 sky130_fd_sc_hd__a2bb2o_1 _23875_ (.A1_N(_07974_),
    .A2_N(_07977_),
    .B1(_07974_),
    .B2(_07977_),
    .X(_07978_));
 sky130_fd_sc_hd__or2_1 _23876_ (.A(_07973_),
    .B(_07978_),
    .X(_07979_));
 sky130_fd_sc_hd__a21bo_1 _23877_ (.A1(_07973_),
    .A2(_07978_),
    .B1_N(_07979_),
    .X(_07980_));
 sky130_fd_sc_hd__o21ba_1 _23878_ (.A1(_07837_),
    .A2(_07840_),
    .B1_N(_07839_),
    .X(_07981_));
 sky130_fd_sc_hd__o21ba_1 _23879_ (.A1(_07829_),
    .A2(_07834_),
    .B1_N(_07831_),
    .X(_07982_));
 sky130_fd_sc_hd__clkbuf_2 _23880_ (.A(_06101_),
    .X(_07983_));
 sky130_fd_sc_hd__or2_1 _23881_ (.A(_07688_),
    .B(_07983_),
    .X(_07984_));
 sky130_fd_sc_hd__o22a_1 _23882_ (.A1(_07690_),
    .A2(_06939_),
    .B1(_07691_),
    .B2(_06544_),
    .X(_07985_));
 sky130_fd_sc_hd__and4_2 _23883_ (.A(_07536_),
    .B(_13612_),
    .C(_13091_),
    .D(_06007_),
    .X(_07986_));
 sky130_fd_sc_hd__or2_1 _23884_ (.A(_07985_),
    .B(_07986_),
    .X(_07987_));
 sky130_fd_sc_hd__a2bb2o_1 _23885_ (.A1_N(_07984_),
    .A2_N(_07987_),
    .B1(_07984_),
    .B2(_07987_),
    .X(_07988_));
 sky130_fd_sc_hd__a2bb2o_1 _23886_ (.A1_N(_07982_),
    .A2_N(_07988_),
    .B1(_07982_),
    .B2(_07988_),
    .X(_07989_));
 sky130_fd_sc_hd__a2bb2o_1 _23887_ (.A1_N(_07981_),
    .A2_N(_07989_),
    .B1(_07981_),
    .B2(_07989_),
    .X(_07990_));
 sky130_fd_sc_hd__or2_1 _23888_ (.A(_07980_),
    .B(_07990_),
    .X(_07991_));
 sky130_fd_sc_hd__a21bo_1 _23889_ (.A1(_07980_),
    .A2(_07990_),
    .B1_N(_07991_),
    .X(_07992_));
 sky130_fd_sc_hd__a2bb2o_1 _23890_ (.A1_N(_07844_),
    .A2_N(_07992_),
    .B1(_07844_),
    .B2(_07992_),
    .X(_07993_));
 sky130_fd_sc_hd__a2bb2o_1 _23891_ (.A1_N(_07969_),
    .A2_N(_07993_),
    .B1(_07969_),
    .B2(_07993_),
    .X(_07994_));
 sky130_fd_sc_hd__o22a_1 _23892_ (.A1(_07698_),
    .A2(_07845_),
    .B1(_07828_),
    .B2(_07846_),
    .X(_07995_));
 sky130_fd_sc_hd__a2bb2o_1 _23893_ (.A1_N(_07994_),
    .A2_N(_07995_),
    .B1(_07994_),
    .B2(_07995_),
    .X(_07996_));
 sky130_fd_sc_hd__a2bb2o_1 _23894_ (.A1_N(_07952_),
    .A2_N(_07996_),
    .B1(_07952_),
    .B2(_07996_),
    .X(_07997_));
 sky130_fd_sc_hd__o22a_1 _23895_ (.A1(_07847_),
    .A2(_07848_),
    .B1(_07809_),
    .B2(_07849_),
    .X(_07998_));
 sky130_fd_sc_hd__a2bb2o_1 _23896_ (.A1_N(_07997_),
    .A2_N(_07998_),
    .B1(_07997_),
    .B2(_07998_),
    .X(_07999_));
 sky130_fd_sc_hd__a2bb2o_4 _23897_ (.A1_N(_07921_),
    .A2_N(_07999_),
    .B1(_07921_),
    .B2(_07999_),
    .X(_08000_));
 sky130_fd_sc_hd__o22a_1 _23898_ (.A1(_07850_),
    .A2(_07851_),
    .B1(_07777_),
    .B2(_07852_),
    .X(_08001_));
 sky130_fd_sc_hd__a2bb2o_1 _23899_ (.A1_N(_08000_),
    .A2_N(_08001_),
    .B1(_08000_),
    .B2(_08001_),
    .X(_08002_));
 sky130_fd_sc_hd__a2bb2o_1 _23900_ (.A1_N(_07866_),
    .A2_N(_08002_),
    .B1(_07866_),
    .B2(_08002_),
    .X(_08003_));
 sky130_fd_sc_hd__o22a_1 _23901_ (.A1(_07853_),
    .A2(_07854_),
    .B1(_07727_),
    .B2(_07855_),
    .X(_08004_));
 sky130_fd_sc_hd__a2bb2o_1 _23902_ (.A1_N(_08003_),
    .A2_N(_08004_),
    .B1(_08003_),
    .B2(_08004_),
    .X(_08005_));
 sky130_fd_sc_hd__a2bb2o_1 _23903_ (.A1_N(_07726_),
    .A2_N(_08005_),
    .B1(_07726_),
    .B2(_08005_),
    .X(_08006_));
 sky130_fd_sc_hd__o22a_1 _23904_ (.A1(_07856_),
    .A2(_07857_),
    .B1(_07582_),
    .B2(_07858_),
    .X(_08007_));
 sky130_fd_sc_hd__or2_1 _23905_ (.A(_08006_),
    .B(_08007_),
    .X(_08008_));
 sky130_fd_sc_hd__a21bo_1 _23906_ (.A1(_08006_),
    .A2(_08007_),
    .B1_N(_08008_),
    .X(_08009_));
 sky130_fd_sc_hd__a22o_1 _23907_ (.A1(_07723_),
    .A2(_07859_),
    .B1(_07714_),
    .B2(_07860_),
    .X(_08010_));
 sky130_fd_sc_hd__o31a_1 _23908_ (.A1(_07716_),
    .A2(_07861_),
    .A3(_07721_),
    .B1(_08010_),
    .X(_08011_));
 sky130_fd_sc_hd__a2bb2oi_2 _23909_ (.A1_N(_08009_),
    .A2_N(_08011_),
    .B1(_08009_),
    .B2(_08011_),
    .Y(_02649_));
 sky130_fd_sc_hd__o22a_1 _23910_ (.A1(_08003_),
    .A2(_08004_),
    .B1(_07726_),
    .B2(_08005_),
    .X(_08012_));
 sky130_fd_sc_hd__o22a_1 _23911_ (.A1(_07868_),
    .A2(_07919_),
    .B1(_07867_),
    .B2(_07920_),
    .X(_08013_));
 sky130_fd_sc_hd__o22a_4 _23912_ (.A1(_07897_),
    .A2(_07898_),
    .B1(_07869_),
    .B2(_07899_),
    .X(_08014_));
 sky130_fd_sc_hd__or2_2 _23913_ (.A(_08013_),
    .B(_08014_),
    .X(_08015_));
 sky130_fd_sc_hd__a21bo_1 _23914_ (.A1(_08013_),
    .A2(_08014_),
    .B1_N(_08015_),
    .X(_08016_));
 sky130_fd_sc_hd__o22a_1 _23915_ (.A1(_07916_),
    .A2(_07917_),
    .B1(_07900_),
    .B2(_07918_),
    .X(_08017_));
 sky130_fd_sc_hd__o22a_4 _23916_ (.A1(_07923_),
    .A2(_07950_),
    .B1(_07922_),
    .B2(_07951_),
    .X(_08018_));
 sky130_fd_sc_hd__a21oi_2 _23917_ (.A1(_07880_),
    .A2(_07882_),
    .B1(_07879_),
    .Y(_08019_));
 sky130_fd_sc_hd__clkbuf_2 _23918_ (.A(_07891_),
    .X(_08020_));
 sky130_fd_sc_hd__o22a_1 _23919_ (.A1(_06876_),
    .A2(_07874_),
    .B1(_05308_),
    .B2(_08020_),
    .X(_08021_));
 sky130_fd_sc_hd__buf_1 _23920_ (.A(\pcpi_mul.rs1[29] ),
    .X(_08022_));
 sky130_fd_sc_hd__buf_1 _23921_ (.A(_08022_),
    .X(_08023_));
 sky130_fd_sc_hd__buf_1 _23922_ (.A(_08023_),
    .X(_08024_));
 sky130_fd_sc_hd__and4_1 _23923_ (.A(_13175_),
    .B(_08024_),
    .C(_13180_),
    .D(_13511_),
    .X(_08025_));
 sky130_fd_sc_hd__nor2_2 _23924_ (.A(_08021_),
    .B(_08025_),
    .Y(_08026_));
 sky130_fd_sc_hd__buf_2 _23925_ (.A(_07596_),
    .X(_08027_));
 sky130_fd_sc_hd__nor2_2 _23926_ (.A(_06887_),
    .B(_08027_),
    .Y(_08028_));
 sky130_fd_sc_hd__a2bb2o_1 _23927_ (.A1_N(_08026_),
    .A2_N(_08028_),
    .B1(_08026_),
    .B2(_08028_),
    .X(_08029_));
 sky130_fd_sc_hd__o22a_1 _23928_ (.A1(_07182_),
    .A2(_07736_),
    .B1(_07184_),
    .B2(_07733_),
    .X(_08030_));
 sky130_fd_sc_hd__and4_2 _23929_ (.A(_13162_),
    .B(_13529_),
    .C(_13168_),
    .D(_13524_),
    .X(_08031_));
 sky130_fd_sc_hd__nor2_2 _23930_ (.A(_08030_),
    .B(_08031_),
    .Y(_08032_));
 sky130_vsdinv _23931_ (.A(\pcpi_mul.rs1[31] ),
    .Y(_08033_));
 sky130_fd_sc_hd__clkbuf_2 _23932_ (.A(_08033_),
    .X(_08034_));
 sky130_fd_sc_hd__clkbuf_2 _23933_ (.A(_08034_),
    .X(_08035_));
 sky130_fd_sc_hd__buf_2 _23934_ (.A(_08035_),
    .X(_08036_));
 sky130_fd_sc_hd__nor2_2 _23935_ (.A(_05143_),
    .B(_08036_),
    .Y(_08037_));
 sky130_fd_sc_hd__a2bb2o_1 _23936_ (.A1_N(_08032_),
    .A2_N(_08037_),
    .B1(_08032_),
    .B2(_08037_),
    .X(_08038_));
 sky130_fd_sc_hd__a21oi_2 _23937_ (.A1(_07888_),
    .A2(_07893_),
    .B1(_07887_),
    .Y(_08039_));
 sky130_fd_sc_hd__a2bb2o_1 _23938_ (.A1_N(_08038_),
    .A2_N(_08039_),
    .B1(_08038_),
    .B2(_08039_),
    .X(_08040_));
 sky130_fd_sc_hd__a2bb2o_1 _23939_ (.A1_N(_08029_),
    .A2_N(_08040_),
    .B1(_08029_),
    .B2(_08040_),
    .X(_08041_));
 sky130_fd_sc_hd__o22a_1 _23940_ (.A1(_07894_),
    .A2(_07895_),
    .B1(_07883_),
    .B2(_07896_),
    .X(_08042_));
 sky130_fd_sc_hd__a2bb2o_1 _23941_ (.A1_N(_08041_),
    .A2_N(_08042_),
    .B1(_08041_),
    .B2(_08042_),
    .X(_08043_));
 sky130_fd_sc_hd__a2bb2o_2 _23942_ (.A1_N(_08019_),
    .A2_N(_08043_),
    .B1(_08019_),
    .B2(_08043_),
    .X(_08044_));
 sky130_fd_sc_hd__o22a_1 _23943_ (.A1(_07904_),
    .A2(_07912_),
    .B1(_07903_),
    .B2(_07913_),
    .X(_08045_));
 sky130_fd_sc_hd__o22a_1 _23944_ (.A1(_07934_),
    .A2(_07935_),
    .B1(_07928_),
    .B2(_07936_),
    .X(_08046_));
 sky130_fd_sc_hd__a21oi_2 _23945_ (.A1(_07910_),
    .A2(_07911_),
    .B1(_07909_),
    .Y(_08047_));
 sky130_fd_sc_hd__o21ba_1 _23946_ (.A1(_07924_),
    .A2(_07927_),
    .B1_N(_07926_),
    .X(_08048_));
 sky130_fd_sc_hd__buf_1 _23947_ (.A(_06671_),
    .X(_08049_));
 sky130_fd_sc_hd__buf_1 _23948_ (.A(_06890_),
    .X(_08050_));
 sky130_fd_sc_hd__o22a_1 _23949_ (.A1(_08049_),
    .A2(_08050_),
    .B1(_05458_),
    .B2(_07744_),
    .X(_08051_));
 sky130_fd_sc_hd__buf_1 _23950_ (.A(_05870_),
    .X(_08052_));
 sky130_fd_sc_hd__buf_1 _23951_ (.A(_13541_),
    .X(_08053_));
 sky130_fd_sc_hd__buf_1 _23952_ (.A(_05871_),
    .X(_08054_));
 sky130_fd_sc_hd__and4_1 _23953_ (.A(_08052_),
    .B(_08053_),
    .C(_08054_),
    .D(_07740_),
    .X(_08055_));
 sky130_fd_sc_hd__nor2_2 _23954_ (.A(_08051_),
    .B(_08055_),
    .Y(_08056_));
 sky130_fd_sc_hd__buf_2 _23955_ (.A(_05460_),
    .X(_08057_));
 sky130_fd_sc_hd__nor2_2 _23956_ (.A(_08057_),
    .B(_07453_),
    .Y(_08058_));
 sky130_fd_sc_hd__a2bb2o_1 _23957_ (.A1_N(_08056_),
    .A2_N(_08058_),
    .B1(_08056_),
    .B2(_08058_),
    .X(_08059_));
 sky130_fd_sc_hd__a2bb2o_1 _23958_ (.A1_N(_08048_),
    .A2_N(_08059_),
    .B1(_08048_),
    .B2(_08059_),
    .X(_08060_));
 sky130_fd_sc_hd__a2bb2o_1 _23959_ (.A1_N(_08047_),
    .A2_N(_08060_),
    .B1(_08047_),
    .B2(_08060_),
    .X(_08061_));
 sky130_fd_sc_hd__a2bb2o_1 _23960_ (.A1_N(_08046_),
    .A2_N(_08061_),
    .B1(_08046_),
    .B2(_08061_),
    .X(_08062_));
 sky130_fd_sc_hd__a2bb2o_1 _23961_ (.A1_N(_08045_),
    .A2_N(_08062_),
    .B1(_08045_),
    .B2(_08062_),
    .X(_08063_));
 sky130_fd_sc_hd__o22a_1 _23962_ (.A1(_07902_),
    .A2(_07914_),
    .B1(_07901_),
    .B2(_07915_),
    .X(_08064_));
 sky130_fd_sc_hd__a2bb2o_1 _23963_ (.A1_N(_08063_),
    .A2_N(_08064_),
    .B1(_08063_),
    .B2(_08064_),
    .X(_08065_));
 sky130_fd_sc_hd__a2bb2o_1 _23964_ (.A1_N(_08044_),
    .A2_N(_08065_),
    .B1(_08044_),
    .B2(_08065_),
    .X(_08066_));
 sky130_fd_sc_hd__a2bb2o_1 _23965_ (.A1_N(_08018_),
    .A2_N(_08066_),
    .B1(_08018_),
    .B2(_08066_),
    .X(_08067_));
 sky130_fd_sc_hd__a2bb2o_2 _23966_ (.A1_N(_08017_),
    .A2_N(_08067_),
    .B1(_08017_),
    .B2(_08067_),
    .X(_08068_));
 sky130_fd_sc_hd__o22a_1 _23967_ (.A1(_07947_),
    .A2(_07948_),
    .B1(_07937_),
    .B2(_07949_),
    .X(_08069_));
 sky130_fd_sc_hd__o22a_1 _23968_ (.A1(_07954_),
    .A2(_07967_),
    .B1(_07953_),
    .B2(_07968_),
    .X(_08070_));
 sky130_fd_sc_hd__or2_1 _23969_ (.A(_07105_),
    .B(_07613_),
    .X(_08071_));
 sky130_fd_sc_hd__o22a_1 _23970_ (.A1(_06822_),
    .A2(_06574_),
    .B1(_06960_),
    .B2(_06649_),
    .X(_08072_));
 sky130_fd_sc_hd__and4_1 _23971_ (.A(_06962_),
    .B(_07039_),
    .C(_06963_),
    .D(_07190_),
    .X(_08073_));
 sky130_fd_sc_hd__or2_1 _23972_ (.A(_08072_),
    .B(_08073_),
    .X(_08074_));
 sky130_fd_sc_hd__a2bb2o_1 _23973_ (.A1_N(_08071_),
    .A2_N(_08074_),
    .B1(_08071_),
    .B2(_08074_),
    .X(_08075_));
 sky130_fd_sc_hd__or2_1 _23974_ (.A(_07369_),
    .B(_07036_),
    .X(_08076_));
 sky130_fd_sc_hd__o22a_1 _23975_ (.A1(_06969_),
    .A2(_06328_),
    .B1(_07930_),
    .B2(_06338_),
    .X(_08077_));
 sky130_fd_sc_hd__and4_1 _23976_ (.A(_06972_),
    .B(_07501_),
    .C(_06973_),
    .D(_13559_),
    .X(_08078_));
 sky130_fd_sc_hd__or2_1 _23977_ (.A(_08077_),
    .B(_08078_),
    .X(_08079_));
 sky130_fd_sc_hd__a2bb2o_1 _23978_ (.A1_N(_08076_),
    .A2_N(_08079_),
    .B1(_08076_),
    .B2(_08079_),
    .X(_08080_));
 sky130_fd_sc_hd__o21ba_1 _23979_ (.A1(_07929_),
    .A2(_07933_),
    .B1_N(_07932_),
    .X(_08081_));
 sky130_fd_sc_hd__a2bb2o_1 _23980_ (.A1_N(_08080_),
    .A2_N(_08081_),
    .B1(_08080_),
    .B2(_08081_),
    .X(_08082_));
 sky130_fd_sc_hd__a2bb2o_2 _23981_ (.A1_N(_08075_),
    .A2_N(_08082_),
    .B1(_08075_),
    .B2(_08082_),
    .X(_08083_));
 sky130_fd_sc_hd__o21ba_1 _23982_ (.A1(_07940_),
    .A2(_07944_),
    .B1_N(_07943_),
    .X(_08084_));
 sky130_fd_sc_hd__o21ba_1 _23983_ (.A1(_07955_),
    .A2(_07958_),
    .B1_N(_07957_),
    .X(_08085_));
 sky130_fd_sc_hd__or2_1 _23984_ (.A(_07516_),
    .B(_06783_),
    .X(_08086_));
 sky130_fd_sc_hd__o22a_1 _23985_ (.A1(_07941_),
    .A2(_06598_),
    .B1(_06089_),
    .B2(_06131_),
    .X(_08087_));
 sky130_fd_sc_hd__and4_1 _23986_ (.A(_07798_),
    .B(_13575_),
    .C(_07799_),
    .D(_06786_),
    .X(_08088_));
 sky130_fd_sc_hd__or2_1 _23987_ (.A(_08087_),
    .B(_08088_),
    .X(_08089_));
 sky130_fd_sc_hd__a2bb2o_1 _23988_ (.A1_N(_08086_),
    .A2_N(_08089_),
    .B1(_08086_),
    .B2(_08089_),
    .X(_08090_));
 sky130_fd_sc_hd__a2bb2o_1 _23989_ (.A1_N(_08085_),
    .A2_N(_08090_),
    .B1(_08085_),
    .B2(_08090_),
    .X(_08091_));
 sky130_fd_sc_hd__a2bb2o_1 _23990_ (.A1_N(_08084_),
    .A2_N(_08091_),
    .B1(_08084_),
    .B2(_08091_),
    .X(_08092_));
 sky130_fd_sc_hd__o22a_1 _23991_ (.A1(_07939_),
    .A2(_07945_),
    .B1(_07938_),
    .B2(_07946_),
    .X(_08093_));
 sky130_fd_sc_hd__a2bb2o_1 _23992_ (.A1_N(_08092_),
    .A2_N(_08093_),
    .B1(_08092_),
    .B2(_08093_),
    .X(_08094_));
 sky130_fd_sc_hd__a2bb2o_1 _23993_ (.A1_N(_08083_),
    .A2_N(_08094_),
    .B1(_08083_),
    .B2(_08094_),
    .X(_08095_));
 sky130_fd_sc_hd__a2bb2o_1 _23994_ (.A1_N(_08070_),
    .A2_N(_08095_),
    .B1(_08070_),
    .B2(_08095_),
    .X(_08096_));
 sky130_fd_sc_hd__a2bb2o_1 _23995_ (.A1_N(_08069_),
    .A2_N(_08096_),
    .B1(_08069_),
    .B2(_08096_),
    .X(_08097_));
 sky130_fd_sc_hd__o22a_1 _23996_ (.A1(_07964_),
    .A2(_07965_),
    .B1(_07959_),
    .B2(_07966_),
    .X(_08098_));
 sky130_fd_sc_hd__o22a_1 _23997_ (.A1(_07982_),
    .A2(_07988_),
    .B1(_07981_),
    .B2(_07989_),
    .X(_08099_));
 sky130_fd_sc_hd__or2_1 _23998_ (.A(_07546_),
    .B(_06479_),
    .X(_08100_));
 sky130_fd_sc_hd__o22a_1 _23999_ (.A1(_07812_),
    .A2(_06704_),
    .B1(_06395_),
    .B2(_06356_),
    .X(_08101_));
 sky130_fd_sc_hd__buf_1 _24000_ (.A(_06941_),
    .X(_08102_));
 sky130_fd_sc_hd__and4_1 _24001_ (.A(_07549_),
    .B(_07117_),
    .C(_08102_),
    .D(_06234_),
    .X(_08103_));
 sky130_fd_sc_hd__or2_1 _24002_ (.A(_08101_),
    .B(_08103_),
    .X(_08104_));
 sky130_fd_sc_hd__a2bb2o_1 _24003_ (.A1_N(_08100_),
    .A2_N(_08104_),
    .B1(_08100_),
    .B2(_08104_),
    .X(_08105_));
 sky130_fd_sc_hd__or2_1 _24004_ (.A(_06803_),
    .B(_06399_),
    .X(_08106_));
 sky130_fd_sc_hd__o22a_1 _24005_ (.A1(_07665_),
    .A2(_06983_),
    .B1(_07818_),
    .B2(_07255_),
    .X(_08107_));
 sky130_fd_sc_hd__and4_1 _24006_ (.A(_13097_),
    .B(_07249_),
    .C(_13102_),
    .D(_06526_),
    .X(_08108_));
 sky130_fd_sc_hd__or2_1 _24007_ (.A(_08107_),
    .B(_08108_),
    .X(_08109_));
 sky130_fd_sc_hd__a2bb2o_1 _24008_ (.A1_N(_08106_),
    .A2_N(_08109_),
    .B1(_08106_),
    .B2(_08109_),
    .X(_08110_));
 sky130_fd_sc_hd__o21ba_1 _24009_ (.A1(_07960_),
    .A2(_07963_),
    .B1_N(_07962_),
    .X(_08111_));
 sky130_fd_sc_hd__a2bb2o_1 _24010_ (.A1_N(_08110_),
    .A2_N(_08111_),
    .B1(_08110_),
    .B2(_08111_),
    .X(_08112_));
 sky130_fd_sc_hd__a2bb2o_1 _24011_ (.A1_N(_08105_),
    .A2_N(_08112_),
    .B1(_08105_),
    .B2(_08112_),
    .X(_08113_));
 sky130_fd_sc_hd__a2bb2o_1 _24012_ (.A1_N(_08099_),
    .A2_N(_08113_),
    .B1(_08099_),
    .B2(_08113_),
    .X(_08114_));
 sky130_fd_sc_hd__a2bb2o_1 _24013_ (.A1_N(_08098_),
    .A2_N(_08114_),
    .B1(_08098_),
    .B2(_08114_),
    .X(_08115_));
 sky130_fd_sc_hd__o21ba_1 _24014_ (.A1(_07984_),
    .A2(_07987_),
    .B1_N(_07986_),
    .X(_08116_));
 sky130_fd_sc_hd__o21ba_1 _24015_ (.A1(_07974_),
    .A2(_07977_),
    .B1_N(_07975_),
    .X(_08117_));
 sky130_fd_sc_hd__clkbuf_2 _24016_ (.A(_07688_),
    .X(_08118_));
 sky130_fd_sc_hd__or2_1 _24017_ (.A(_08118_),
    .B(_07278_),
    .X(_08119_));
 sky130_fd_sc_hd__clkbuf_2 _24018_ (.A(_07690_),
    .X(_08120_));
 sky130_fd_sc_hd__clkbuf_2 _24019_ (.A(_07691_),
    .X(_08121_));
 sky130_fd_sc_hd__o22a_1 _24020_ (.A1(_08120_),
    .A2(_05900_),
    .B1(_08121_),
    .B2(_07983_),
    .X(_08122_));
 sky130_fd_sc_hd__clkbuf_2 _24021_ (.A(_13087_),
    .X(_08123_));
 sky130_fd_sc_hd__clkbuf_2 _24022_ (.A(_07395_),
    .X(_08124_));
 sky130_fd_sc_hd__and4_1 _24023_ (.A(_08123_),
    .B(_13609_),
    .C(_08124_),
    .D(_07405_),
    .X(_08125_));
 sky130_fd_sc_hd__or2_1 _24024_ (.A(_08122_),
    .B(_08125_),
    .X(_08126_));
 sky130_fd_sc_hd__a2bb2o_1 _24025_ (.A1_N(_08119_),
    .A2_N(_08126_),
    .B1(_08119_),
    .B2(_08126_),
    .X(_08127_));
 sky130_fd_sc_hd__a2bb2o_1 _24026_ (.A1_N(_08117_),
    .A2_N(_08127_),
    .B1(_08117_),
    .B2(_08127_),
    .X(_08128_));
 sky130_fd_sc_hd__a2bb2o_1 _24027_ (.A1_N(_08116_),
    .A2_N(_08128_),
    .B1(_08116_),
    .B2(_08128_),
    .X(_08129_));
 sky130_vsdinv _24028_ (.A(\pcpi_mul.rs2[31] ),
    .Y(_08130_));
 sky130_fd_sc_hd__buf_1 _24029_ (.A(_08130_),
    .X(_08131_));
 sky130_fd_sc_hd__clkbuf_2 _24030_ (.A(_08131_),
    .X(_08132_));
 sky130_fd_sc_hd__o22a_1 _24031_ (.A1(_08132_),
    .A2(_05325_),
    .B1(_07971_),
    .B2(_05319_),
    .X(_08133_));
 sky130_fd_sc_hd__or4_4 _24032_ (.A(_08132_),
    .B(_05149_),
    .C(_07971_),
    .D(_05297_),
    .X(_08134_));
 sky130_fd_sc_hd__or2b_1 _24033_ (.A(_08133_),
    .B_N(_08134_),
    .X(_08135_));
 sky130_fd_sc_hd__buf_1 _24034_ (.A(_06939_),
    .X(_08136_));
 sky130_fd_sc_hd__or2_1 _24035_ (.A(_07530_),
    .B(_08136_),
    .X(_08137_));
 sky130_fd_sc_hd__and4_1 _24036_ (.A(_13072_),
    .B(_06115_),
    .C(_07830_),
    .D(_06116_),
    .X(_08138_));
 sky130_fd_sc_hd__o22a_1 _24037_ (.A1(_07832_),
    .A2(_05315_),
    .B1(_07677_),
    .B2(_06112_),
    .X(_08139_));
 sky130_fd_sc_hd__or2_1 _24038_ (.A(_08138_),
    .B(_08139_),
    .X(_08140_));
 sky130_fd_sc_hd__a2bb2o_1 _24039_ (.A1_N(_08137_),
    .A2_N(_08140_),
    .B1(_08137_),
    .B2(_08140_),
    .X(_08141_));
 sky130_fd_sc_hd__or2_1 _24040_ (.A(_08135_),
    .B(_08141_),
    .X(_08142_));
 sky130_fd_sc_hd__a21bo_1 _24041_ (.A1(_08135_),
    .A2(_08141_),
    .B1_N(_08142_),
    .X(_08143_));
 sky130_fd_sc_hd__a2bb2o_1 _24042_ (.A1_N(_07979_),
    .A2_N(_08143_),
    .B1(_07979_),
    .B2(_08143_),
    .X(_08144_));
 sky130_fd_sc_hd__a2bb2o_1 _24043_ (.A1_N(_08129_),
    .A2_N(_08144_),
    .B1(_08129_),
    .B2(_08144_),
    .X(_08145_));
 sky130_fd_sc_hd__a2bb2o_1 _24044_ (.A1_N(_07991_),
    .A2_N(_08145_),
    .B1(_07991_),
    .B2(_08145_),
    .X(_08146_));
 sky130_fd_sc_hd__a2bb2o_1 _24045_ (.A1_N(_08115_),
    .A2_N(_08146_),
    .B1(_08115_),
    .B2(_08146_),
    .X(_08147_));
 sky130_fd_sc_hd__o22a_1 _24046_ (.A1(_07844_),
    .A2(_07992_),
    .B1(_07969_),
    .B2(_07993_),
    .X(_08148_));
 sky130_fd_sc_hd__a2bb2o_1 _24047_ (.A1_N(_08147_),
    .A2_N(_08148_),
    .B1(_08147_),
    .B2(_08148_),
    .X(_08149_));
 sky130_fd_sc_hd__a2bb2o_1 _24048_ (.A1_N(_08097_),
    .A2_N(_08149_),
    .B1(_08097_),
    .B2(_08149_),
    .X(_08150_));
 sky130_fd_sc_hd__o22a_1 _24049_ (.A1(_07994_),
    .A2(_07995_),
    .B1(_07952_),
    .B2(_07996_),
    .X(_08151_));
 sky130_fd_sc_hd__a2bb2o_1 _24050_ (.A1_N(_08150_),
    .A2_N(_08151_),
    .B1(_08150_),
    .B2(_08151_),
    .X(_08152_));
 sky130_fd_sc_hd__a2bb2o_1 _24051_ (.A1_N(_08068_),
    .A2_N(_08152_),
    .B1(_08068_),
    .B2(_08152_),
    .X(_08153_));
 sky130_fd_sc_hd__o22a_1 _24052_ (.A1(_07997_),
    .A2(_07998_),
    .B1(_07921_),
    .B2(_07999_),
    .X(_08154_));
 sky130_fd_sc_hd__a2bb2o_1 _24053_ (.A1_N(_08153_),
    .A2_N(_08154_),
    .B1(_08153_),
    .B2(_08154_),
    .X(_08155_));
 sky130_fd_sc_hd__a2bb2o_4 _24054_ (.A1_N(_08016_),
    .A2_N(_08155_),
    .B1(_08016_),
    .B2(_08155_),
    .X(_08156_));
 sky130_fd_sc_hd__o22a_1 _24055_ (.A1(_08000_),
    .A2(_08001_),
    .B1(_07866_),
    .B2(_08002_),
    .X(_08157_));
 sky130_fd_sc_hd__a2bb2o_1 _24056_ (.A1_N(_08156_),
    .A2_N(_08157_),
    .B1(_08156_),
    .B2(_08157_),
    .X(_08158_));
 sky130_fd_sc_hd__a2bb2o_1 _24057_ (.A1_N(_07865_),
    .A2_N(_08158_),
    .B1(_07865_),
    .B2(_08158_),
    .X(_08159_));
 sky130_fd_sc_hd__and2_1 _24058_ (.A(_08012_),
    .B(_08159_),
    .X(_08160_));
 sky130_fd_sc_hd__or2_1 _24059_ (.A(_08012_),
    .B(_08159_),
    .X(_08161_));
 sky130_fd_sc_hd__or2b_1 _24060_ (.A(_08160_),
    .B_N(_08161_),
    .X(_08162_));
 sky130_fd_sc_hd__o21ai_1 _24061_ (.A1(_08009_),
    .A2(_08011_),
    .B1(_08008_),
    .Y(_08163_));
 sky130_fd_sc_hd__a2bb2o_1 _24062_ (.A1_N(_08162_),
    .A2_N(_08163_),
    .B1(_08162_),
    .B2(_08163_),
    .X(_02650_));
 sky130_fd_sc_hd__o22a_2 _24063_ (.A1(_08018_),
    .A2(_08066_),
    .B1(_08017_),
    .B2(_08067_),
    .X(_08164_));
 sky130_fd_sc_hd__o22a_1 _24064_ (.A1(_08041_),
    .A2(_08042_),
    .B1(_08019_),
    .B2(_08043_),
    .X(_08165_));
 sky130_fd_sc_hd__a2bb2o_2 _24065_ (.A1_N(_08164_),
    .A2_N(_08165_),
    .B1(_08164_),
    .B2(_08165_),
    .X(_08166_));
 sky130_fd_sc_hd__a2bb2o_4 _24066_ (.A1_N(_11723_),
    .A2_N(_08166_),
    .B1(_11722_),
    .B2(_08166_),
    .X(_08167_));
 sky130_fd_sc_hd__o22a_4 _24067_ (.A1(_08063_),
    .A2(_08064_),
    .B1(_08044_),
    .B2(_08065_),
    .X(_08168_));
 sky130_fd_sc_hd__o22a_1 _24068_ (.A1(_08070_),
    .A2(_08095_),
    .B1(_08069_),
    .B2(_08096_),
    .X(_08169_));
 sky130_fd_sc_hd__a21oi_4 _24069_ (.A1(_08026_),
    .A2(_08028_),
    .B1(_08025_),
    .Y(_08170_));
 sky130_fd_sc_hd__o22a_1 _24070_ (.A1(_06876_),
    .A2(_08020_),
    .B1(_07017_),
    .B2(_08036_),
    .X(_08171_));
 sky130_fd_sc_hd__buf_1 _24071_ (.A(_13509_),
    .X(_08172_));
 sky130_fd_sc_hd__and4_1 _24072_ (.A(_13175_),
    .B(_08172_),
    .C(_13180_),
    .D(_13506_),
    .X(_08173_));
 sky130_fd_sc_hd__nor2_2 _24073_ (.A(_08171_),
    .B(_08173_),
    .Y(_08174_));
 sky130_fd_sc_hd__clkbuf_2 _24074_ (.A(_07749_),
    .X(_08175_));
 sky130_fd_sc_hd__nor2_2 _24075_ (.A(_06887_),
    .B(_08175_),
    .Y(_08176_));
 sky130_fd_sc_hd__a2bb2o_1 _24076_ (.A1_N(_08174_),
    .A2_N(_08176_),
    .B1(_08174_),
    .B2(_08176_),
    .X(_08177_));
 sky130_fd_sc_hd__clkbuf_2 _24077_ (.A(_07732_),
    .X(_08178_));
 sky130_fd_sc_hd__buf_1 _24078_ (.A(_07594_),
    .X(_08179_));
 sky130_fd_sc_hd__buf_1 _24079_ (.A(_08179_),
    .X(_08180_));
 sky130_fd_sc_hd__o22a_1 _24080_ (.A1(_07182_),
    .A2(_08178_),
    .B1(_07184_),
    .B2(_08180_),
    .X(_08181_));
 sky130_fd_sc_hd__and4_2 _24081_ (.A(_13162_),
    .B(_13524_),
    .C(_13168_),
    .D(_13520_),
    .X(_08182_));
 sky130_fd_sc_hd__nor2_2 _24082_ (.A(_08181_),
    .B(_08182_),
    .Y(_08183_));
 sky130_fd_sc_hd__or2_4 _24083_ (.A(_11702_),
    .B(_05941_),
    .X(_08184_));
 sky130_vsdinv _24084_ (.A(_08184_),
    .Y(_08185_));
 sky130_fd_sc_hd__buf_1 _24085_ (.A(_08185_),
    .X(_08186_));
 sky130_fd_sc_hd__a2bb2o_1 _24086_ (.A1_N(_08183_),
    .A2_N(_08186_),
    .B1(_08183_),
    .B2(_08186_),
    .X(_08187_));
 sky130_fd_sc_hd__a21oi_4 _24087_ (.A1(_08032_),
    .A2(_08037_),
    .B1(_08031_),
    .Y(_08188_));
 sky130_fd_sc_hd__a2bb2o_1 _24088_ (.A1_N(_08187_),
    .A2_N(_08188_),
    .B1(_08187_),
    .B2(_08188_),
    .X(_08189_));
 sky130_fd_sc_hd__a2bb2o_1 _24089_ (.A1_N(_08177_),
    .A2_N(_08189_),
    .B1(_08177_),
    .B2(_08189_),
    .X(_08190_));
 sky130_fd_sc_hd__o22a_2 _24090_ (.A1(_08038_),
    .A2(_08039_),
    .B1(_08029_),
    .B2(_08040_),
    .X(_08191_));
 sky130_fd_sc_hd__a2bb2o_1 _24091_ (.A1_N(_08190_),
    .A2_N(_08191_),
    .B1(_08190_),
    .B2(_08191_),
    .X(_08192_));
 sky130_fd_sc_hd__a2bb2o_2 _24092_ (.A1_N(_08170_),
    .A2_N(_08192_),
    .B1(_08170_),
    .B2(_08192_),
    .X(_08193_));
 sky130_fd_sc_hd__o22a_1 _24093_ (.A1(_08048_),
    .A2(_08059_),
    .B1(_08047_),
    .B2(_08060_),
    .X(_08194_));
 sky130_fd_sc_hd__o22a_1 _24094_ (.A1(_08080_),
    .A2(_08081_),
    .B1(_08075_),
    .B2(_08082_),
    .X(_08195_));
 sky130_fd_sc_hd__a21oi_2 _24095_ (.A1(_08056_),
    .A2(_08058_),
    .B1(_08055_),
    .Y(_08196_));
 sky130_fd_sc_hd__o21ba_1 _24096_ (.A1(_08071_),
    .A2(_08074_),
    .B1_N(_08073_),
    .X(_08197_));
 sky130_fd_sc_hd__buf_1 _24097_ (.A(_07195_),
    .X(_08198_));
 sky130_fd_sc_hd__o22a_1 _24098_ (.A1(_06919_),
    .A2(_07457_),
    .B1(_05458_),
    .B2(_08198_),
    .X(_08199_));
 sky130_fd_sc_hd__buf_1 _24099_ (.A(\pcpi_mul.rs1[24] ),
    .X(_08200_));
 sky130_fd_sc_hd__and4_1 _24100_ (.A(_08052_),
    .B(_08200_),
    .C(_08054_),
    .D(_13534_),
    .X(_08201_));
 sky130_fd_sc_hd__nor2_1 _24101_ (.A(_08199_),
    .B(_08201_),
    .Y(_08202_));
 sky130_fd_sc_hd__nor2_2 _24102_ (.A(_08057_),
    .B(_07884_),
    .Y(_08203_));
 sky130_fd_sc_hd__a2bb2o_1 _24103_ (.A1_N(_08202_),
    .A2_N(_08203_),
    .B1(_08202_),
    .B2(_08203_),
    .X(_08204_));
 sky130_fd_sc_hd__a2bb2o_1 _24104_ (.A1_N(_08197_),
    .A2_N(_08204_),
    .B1(_08197_),
    .B2(_08204_),
    .X(_08205_));
 sky130_fd_sc_hd__a2bb2o_1 _24105_ (.A1_N(_08196_),
    .A2_N(_08205_),
    .B1(_08196_),
    .B2(_08205_),
    .X(_08206_));
 sky130_fd_sc_hd__a2bb2o_1 _24106_ (.A1_N(_08195_),
    .A2_N(_08206_),
    .B1(_08195_),
    .B2(_08206_),
    .X(_08207_));
 sky130_fd_sc_hd__a2bb2o_1 _24107_ (.A1_N(_08194_),
    .A2_N(_08207_),
    .B1(_08194_),
    .B2(_08207_),
    .X(_08208_));
 sky130_fd_sc_hd__o22a_1 _24108_ (.A1(_08046_),
    .A2(_08061_),
    .B1(_08045_),
    .B2(_08062_),
    .X(_08209_));
 sky130_fd_sc_hd__a2bb2o_1 _24109_ (.A1_N(_08208_),
    .A2_N(_08209_),
    .B1(_08208_),
    .B2(_08209_),
    .X(_08210_));
 sky130_fd_sc_hd__a2bb2o_2 _24110_ (.A1_N(_08193_),
    .A2_N(_08210_),
    .B1(_08193_),
    .B2(_08210_),
    .X(_08211_));
 sky130_fd_sc_hd__a2bb2o_1 _24111_ (.A1_N(_08169_),
    .A2_N(_08211_),
    .B1(_08169_),
    .B2(_08211_),
    .X(_08212_));
 sky130_fd_sc_hd__a2bb2o_1 _24112_ (.A1_N(_08168_),
    .A2_N(_08212_),
    .B1(_08168_),
    .B2(_08212_),
    .X(_08213_));
 sky130_fd_sc_hd__o22a_1 _24113_ (.A1(_08092_),
    .A2(_08093_),
    .B1(_08083_),
    .B2(_08094_),
    .X(_08214_));
 sky130_fd_sc_hd__o22a_1 _24114_ (.A1(_08099_),
    .A2(_08113_),
    .B1(_08098_),
    .B2(_08114_),
    .X(_08215_));
 sky130_fd_sc_hd__or2_1 _24115_ (.A(_05537_),
    .B(_07170_),
    .X(_08216_));
 sky130_fd_sc_hd__clkbuf_2 _24116_ (.A(_05714_),
    .X(_08217_));
 sky130_fd_sc_hd__o22a_1 _24117_ (.A1(_08217_),
    .A2(_06649_),
    .B1(_05588_),
    .B2(_06880_),
    .X(_08218_));
 sky130_fd_sc_hd__and4_1 _24118_ (.A(_07363_),
    .B(_07190_),
    .C(_07364_),
    .D(_13545_),
    .X(_08219_));
 sky130_fd_sc_hd__or2_1 _24119_ (.A(_08218_),
    .B(_08219_),
    .X(_08220_));
 sky130_fd_sc_hd__a2bb2o_1 _24120_ (.A1_N(_08216_),
    .A2_N(_08220_),
    .B1(_08216_),
    .B2(_08220_),
    .X(_08221_));
 sky130_fd_sc_hd__or2_1 _24121_ (.A(_07369_),
    .B(_07780_),
    .X(_08222_));
 sky130_fd_sc_hd__buf_2 _24122_ (.A(_06110_),
    .X(_08223_));
 sky130_fd_sc_hd__o22a_1 _24123_ (.A1(_08223_),
    .A2(_06338_),
    .B1(_07930_),
    .B2(_06565_),
    .X(_08224_));
 sky130_fd_sc_hd__and4_1 _24124_ (.A(_07234_),
    .B(_06898_),
    .C(_07235_),
    .D(_07484_),
    .X(_08225_));
 sky130_fd_sc_hd__or2_1 _24125_ (.A(_08224_),
    .B(_08225_),
    .X(_08226_));
 sky130_fd_sc_hd__a2bb2o_1 _24126_ (.A1_N(_08222_),
    .A2_N(_08226_),
    .B1(_08222_),
    .B2(_08226_),
    .X(_08227_));
 sky130_fd_sc_hd__o21ba_1 _24127_ (.A1(_08076_),
    .A2(_08079_),
    .B1_N(_08078_),
    .X(_08228_));
 sky130_fd_sc_hd__a2bb2o_1 _24128_ (.A1_N(_08227_),
    .A2_N(_08228_),
    .B1(_08227_),
    .B2(_08228_),
    .X(_08229_));
 sky130_fd_sc_hd__a2bb2o_2 _24129_ (.A1_N(_08221_),
    .A2_N(_08229_),
    .B1(_08221_),
    .B2(_08229_),
    .X(_08230_));
 sky130_fd_sc_hd__o21ba_1 _24130_ (.A1(_08086_),
    .A2(_08089_),
    .B1_N(_08088_),
    .X(_08231_));
 sky130_fd_sc_hd__o21ba_1 _24131_ (.A1(_08100_),
    .A2(_08104_),
    .B1_N(_08103_),
    .X(_08232_));
 sky130_fd_sc_hd__clkbuf_2 _24132_ (.A(_07128_),
    .X(_08233_));
 sky130_fd_sc_hd__buf_1 _24133_ (.A(_06039_),
    .X(_08234_));
 sky130_fd_sc_hd__o22a_1 _24134_ (.A1(_08233_),
    .A2(_08234_),
    .B1(_06094_),
    .B2(_06218_),
    .X(_08235_));
 sky130_fd_sc_hd__clkbuf_2 _24135_ (.A(_13117_),
    .X(_08236_));
 sky130_fd_sc_hd__buf_1 _24136_ (.A(_13569_),
    .X(_08237_));
 sky130_fd_sc_hd__clkbuf_2 _24137_ (.A(_13121_),
    .X(_08238_));
 sky130_fd_sc_hd__and4_1 _24138_ (.A(_08236_),
    .B(_08237_),
    .C(_08238_),
    .D(_13567_),
    .X(_08239_));
 sky130_fd_sc_hd__nor2_2 _24139_ (.A(_08235_),
    .B(_08239_),
    .Y(_08240_));
 sky130_fd_sc_hd__clkbuf_2 _24140_ (.A(_06096_),
    .X(_08241_));
 sky130_fd_sc_hd__nor2_2 _24141_ (.A(_08241_),
    .B(_06330_),
    .Y(_08242_));
 sky130_fd_sc_hd__a2bb2o_2 _24142_ (.A1_N(_08240_),
    .A2_N(_08242_),
    .B1(_08240_),
    .B2(_08242_),
    .X(_08243_));
 sky130_fd_sc_hd__a2bb2o_1 _24143_ (.A1_N(_08232_),
    .A2_N(_08243_),
    .B1(_08232_),
    .B2(_08243_),
    .X(_08244_));
 sky130_fd_sc_hd__a2bb2o_1 _24144_ (.A1_N(_08231_),
    .A2_N(_08244_),
    .B1(_08231_),
    .B2(_08244_),
    .X(_08245_));
 sky130_fd_sc_hd__o22a_1 _24145_ (.A1(_08085_),
    .A2(_08090_),
    .B1(_08084_),
    .B2(_08091_),
    .X(_08246_));
 sky130_fd_sc_hd__a2bb2o_1 _24146_ (.A1_N(_08245_),
    .A2_N(_08246_),
    .B1(_08245_),
    .B2(_08246_),
    .X(_08247_));
 sky130_fd_sc_hd__a2bb2o_1 _24147_ (.A1_N(_08230_),
    .A2_N(_08247_),
    .B1(_08230_),
    .B2(_08247_),
    .X(_08248_));
 sky130_fd_sc_hd__a2bb2o_1 _24148_ (.A1_N(_08215_),
    .A2_N(_08248_),
    .B1(_08215_),
    .B2(_08248_),
    .X(_08249_));
 sky130_fd_sc_hd__a2bb2o_1 _24149_ (.A1_N(_08214_),
    .A2_N(_08249_),
    .B1(_08214_),
    .B2(_08249_),
    .X(_08250_));
 sky130_fd_sc_hd__o22a_1 _24150_ (.A1(_08110_),
    .A2(_08111_),
    .B1(_08105_),
    .B2(_08112_),
    .X(_08251_));
 sky130_fd_sc_hd__o22a_1 _24151_ (.A1(_08117_),
    .A2(_08127_),
    .B1(_08116_),
    .B2(_08128_),
    .X(_08252_));
 sky130_fd_sc_hd__clkbuf_2 _24152_ (.A(_06284_),
    .X(_08253_));
 sky130_fd_sc_hd__or2_1 _24153_ (.A(_08253_),
    .B(_06130_),
    .X(_08254_));
 sky130_fd_sc_hd__o22a_1 _24154_ (.A1(_07812_),
    .A2(_06356_),
    .B1(_06390_),
    .B2(_06028_),
    .X(_08255_));
 sky130_fd_sc_hd__clkbuf_2 _24155_ (.A(_13105_),
    .X(_08256_));
 sky130_fd_sc_hd__and4_1 _24156_ (.A(_08256_),
    .B(_13582_),
    .C(_08102_),
    .D(_13579_),
    .X(_08257_));
 sky130_fd_sc_hd__or2_1 _24157_ (.A(_08255_),
    .B(_08257_),
    .X(_08258_));
 sky130_fd_sc_hd__a2bb2o_2 _24158_ (.A1_N(_08254_),
    .A2_N(_08258_),
    .B1(_08254_),
    .B2(_08258_),
    .X(_08259_));
 sky130_fd_sc_hd__or2_1 _24159_ (.A(_06688_),
    .B(_06520_),
    .X(_08260_));
 sky130_fd_sc_hd__clkbuf_2 _24160_ (.A(_06947_),
    .X(_08261_));
 sky130_fd_sc_hd__clkbuf_2 _24161_ (.A(_08261_),
    .X(_08262_));
 sky130_fd_sc_hd__buf_1 _24162_ (.A(_05829_),
    .X(_08263_));
 sky130_fd_sc_hd__o22a_1 _24163_ (.A1(_08262_),
    .A2(_07255_),
    .B1(_07818_),
    .B2(_08263_),
    .X(_08264_));
 sky130_fd_sc_hd__buf_1 _24164_ (.A(_13587_),
    .X(_08265_));
 sky130_fd_sc_hd__and4_1 _24165_ (.A(_13097_),
    .B(_13592_),
    .C(_13102_),
    .D(_08265_),
    .X(_08266_));
 sky130_fd_sc_hd__or2_1 _24166_ (.A(_08264_),
    .B(_08266_),
    .X(_08267_));
 sky130_fd_sc_hd__a2bb2o_1 _24167_ (.A1_N(_08260_),
    .A2_N(_08267_),
    .B1(_08260_),
    .B2(_08267_),
    .X(_08268_));
 sky130_fd_sc_hd__o21ba_1 _24168_ (.A1(_08106_),
    .A2(_08109_),
    .B1_N(_08108_),
    .X(_08269_));
 sky130_fd_sc_hd__a2bb2o_1 _24169_ (.A1_N(_08268_),
    .A2_N(_08269_),
    .B1(_08268_),
    .B2(_08269_),
    .X(_08270_));
 sky130_fd_sc_hd__a2bb2o_1 _24170_ (.A1_N(_08259_),
    .A2_N(_08270_),
    .B1(_08259_),
    .B2(_08270_),
    .X(_08271_));
 sky130_fd_sc_hd__a2bb2o_1 _24171_ (.A1_N(_08252_),
    .A2_N(_08271_),
    .B1(_08252_),
    .B2(_08271_),
    .X(_08272_));
 sky130_fd_sc_hd__a2bb2o_1 _24172_ (.A1_N(_08251_),
    .A2_N(_08272_),
    .B1(_08251_),
    .B2(_08272_),
    .X(_08273_));
 sky130_fd_sc_hd__o21ba_1 _24173_ (.A1(_08119_),
    .A2(_08126_),
    .B1_N(_08125_),
    .X(_08274_));
 sky130_fd_sc_hd__o21ba_1 _24174_ (.A1(_08137_),
    .A2(_08140_),
    .B1_N(_08138_),
    .X(_08275_));
 sky130_fd_sc_hd__or2_1 _24175_ (.A(_08118_),
    .B(_07403_),
    .X(_08276_));
 sky130_fd_sc_hd__o22a_1 _24176_ (.A1(_08120_),
    .A2(_07983_),
    .B1(_08121_),
    .B2(_05862_),
    .X(_08277_));
 sky130_fd_sc_hd__and4_1 _24177_ (.A(_08123_),
    .B(_13604_),
    .C(_08124_),
    .D(_07820_),
    .X(_08278_));
 sky130_fd_sc_hd__or2_1 _24178_ (.A(_08277_),
    .B(_08278_),
    .X(_08279_));
 sky130_fd_sc_hd__a2bb2o_1 _24179_ (.A1_N(_08276_),
    .A2_N(_08279_),
    .B1(_08276_),
    .B2(_08279_),
    .X(_08280_));
 sky130_fd_sc_hd__a2bb2o_1 _24180_ (.A1_N(_08275_),
    .A2_N(_08280_),
    .B1(_08275_),
    .B2(_08280_),
    .X(_08281_));
 sky130_fd_sc_hd__a2bb2o_1 _24181_ (.A1_N(_08274_),
    .A2_N(_08281_),
    .B1(_08274_),
    .B2(_08281_),
    .X(_08282_));
 sky130_fd_sc_hd__buf_1 _24182_ (.A(_06544_),
    .X(_08283_));
 sky130_fd_sc_hd__or2_1 _24183_ (.A(_07681_),
    .B(_08283_),
    .X(_08284_));
 sky130_fd_sc_hd__buf_1 _24184_ (.A(_07832_),
    .X(_08285_));
 sky130_fd_sc_hd__buf_1 _24185_ (.A(_08285_),
    .X(_08286_));
 sky130_fd_sc_hd__buf_1 _24186_ (.A(_07678_),
    .X(_08287_));
 sky130_fd_sc_hd__o22a_1 _24187_ (.A1(_08286_),
    .A2(_05340_),
    .B1(_08287_),
    .B2(_08136_),
    .X(_08288_));
 sky130_fd_sc_hd__and4_1 _24188_ (.A(_13073_),
    .B(_13616_),
    .C(_13078_),
    .D(_13613_),
    .X(_08289_));
 sky130_fd_sc_hd__or2_1 _24189_ (.A(_08288_),
    .B(_08289_),
    .X(_08290_));
 sky130_fd_sc_hd__a2bb2o_1 _24190_ (.A1_N(_08284_),
    .A2_N(_08290_),
    .B1(_08284_),
    .B2(_08290_),
    .X(_08291_));
 sky130_fd_sc_hd__buf_2 _24191_ (.A(_07970_),
    .X(_08292_));
 sky130_fd_sc_hd__or2_1 _24192_ (.A(_08292_),
    .B(_05316_),
    .X(_08293_));
 sky130_fd_sc_hd__buf_1 _24193_ (.A(\pcpi_mul.rs2[32] ),
    .X(_08294_));
 sky130_fd_sc_hd__buf_1 _24194_ (.A(_08294_),
    .X(_08295_));
 sky130_fd_sc_hd__and4_1 _24195_ (.A(_13064_),
    .B(_13624_),
    .C(_08295_),
    .D(_05148_),
    .X(_08296_));
 sky130_fd_sc_hd__o22a_1 _24196_ (.A1(_08131_),
    .A2(_05318_),
    .B1(_11717_),
    .B2(_13626_),
    .X(_08297_));
 sky130_fd_sc_hd__or2_1 _24197_ (.A(_08296_),
    .B(_08297_),
    .X(_08298_));
 sky130_fd_sc_hd__a2bb2o_1 _24198_ (.A1_N(_08293_),
    .A2_N(_08298_),
    .B1(_08293_),
    .B2(_08298_),
    .X(_08299_));
 sky130_fd_sc_hd__a2bb2o_1 _24199_ (.A1_N(_08134_),
    .A2_N(_08299_),
    .B1(_08134_),
    .B2(_08299_),
    .X(_08300_));
 sky130_fd_sc_hd__a2bb2o_1 _24200_ (.A1_N(_08291_),
    .A2_N(_08300_),
    .B1(_08291_),
    .B2(_08300_),
    .X(_08301_));
 sky130_fd_sc_hd__a2bb2o_1 _24201_ (.A1_N(_08142_),
    .A2_N(_08301_),
    .B1(_08142_),
    .B2(_08301_),
    .X(_08302_));
 sky130_fd_sc_hd__a2bb2o_1 _24202_ (.A1_N(_08282_),
    .A2_N(_08302_),
    .B1(_08282_),
    .B2(_08302_),
    .X(_08303_));
 sky130_fd_sc_hd__o22a_1 _24203_ (.A1(_07979_),
    .A2(_08143_),
    .B1(_08129_),
    .B2(_08144_),
    .X(_08304_));
 sky130_fd_sc_hd__a2bb2o_1 _24204_ (.A1_N(_08303_),
    .A2_N(_08304_),
    .B1(_08303_),
    .B2(_08304_),
    .X(_08305_));
 sky130_fd_sc_hd__a2bb2o_1 _24205_ (.A1_N(_08273_),
    .A2_N(_08305_),
    .B1(_08273_),
    .B2(_08305_),
    .X(_08306_));
 sky130_fd_sc_hd__o22a_1 _24206_ (.A1(_07991_),
    .A2(_08145_),
    .B1(_08115_),
    .B2(_08146_),
    .X(_08307_));
 sky130_fd_sc_hd__a2bb2o_1 _24207_ (.A1_N(_08306_),
    .A2_N(_08307_),
    .B1(_08306_),
    .B2(_08307_),
    .X(_08308_));
 sky130_fd_sc_hd__a2bb2o_1 _24208_ (.A1_N(_08250_),
    .A2_N(_08308_),
    .B1(_08250_),
    .B2(_08308_),
    .X(_08309_));
 sky130_fd_sc_hd__o22a_1 _24209_ (.A1(_08147_),
    .A2(_08148_),
    .B1(_08097_),
    .B2(_08149_),
    .X(_08310_));
 sky130_fd_sc_hd__a2bb2o_1 _24210_ (.A1_N(_08309_),
    .A2_N(_08310_),
    .B1(_08309_),
    .B2(_08310_),
    .X(_08311_));
 sky130_fd_sc_hd__a2bb2o_1 _24211_ (.A1_N(_08213_),
    .A2_N(_08311_),
    .B1(_08213_),
    .B2(_08311_),
    .X(_08312_));
 sky130_fd_sc_hd__o22a_1 _24212_ (.A1(_08150_),
    .A2(_08151_),
    .B1(_08068_),
    .B2(_08152_),
    .X(_08313_));
 sky130_fd_sc_hd__a2bb2o_1 _24213_ (.A1_N(_08312_),
    .A2_N(_08313_),
    .B1(_08312_),
    .B2(_08313_),
    .X(_08314_));
 sky130_fd_sc_hd__a2bb2o_1 _24214_ (.A1_N(_08167_),
    .A2_N(_08314_),
    .B1(_08167_),
    .B2(_08314_),
    .X(_08315_));
 sky130_fd_sc_hd__o22a_1 _24215_ (.A1(_08153_),
    .A2(_08154_),
    .B1(_08016_),
    .B2(_08155_),
    .X(_08316_));
 sky130_fd_sc_hd__a2bb2o_1 _24216_ (.A1_N(_08315_),
    .A2_N(_08316_),
    .B1(_08315_),
    .B2(_08316_),
    .X(_08317_));
 sky130_fd_sc_hd__a2bb2o_1 _24217_ (.A1_N(_08015_),
    .A2_N(_08317_),
    .B1(_08015_),
    .B2(_08317_),
    .X(_08318_));
 sky130_fd_sc_hd__o22a_4 _24218_ (.A1(_08156_),
    .A2(_08157_),
    .B1(_07865_),
    .B2(_08158_),
    .X(_08319_));
 sky130_fd_sc_hd__or2_2 _24219_ (.A(_08318_),
    .B(_08319_),
    .X(_08320_));
 sky130_fd_sc_hd__a21bo_1 _24220_ (.A1(_08318_),
    .A2(_08319_),
    .B1_N(_08320_),
    .X(_08321_));
 sky130_fd_sc_hd__buf_2 _24221_ (.A(_08321_),
    .X(_08322_));
 sky130_fd_sc_hd__or2_1 _24222_ (.A(_08009_),
    .B(_08162_),
    .X(_08323_));
 sky130_fd_sc_hd__or3_1 _24223_ (.A(_07715_),
    .B(_07861_),
    .C(_08323_),
    .X(_08324_));
 sky130_fd_sc_hd__or2_2 _24224_ (.A(_07718_),
    .B(_08324_),
    .X(_08325_));
 sky130_fd_sc_hd__o221a_1 _24225_ (.A1(_08008_),
    .A2(_08160_),
    .B1(_08010_),
    .B2(_08323_),
    .C1(_08161_),
    .X(_08326_));
 sky130_fd_sc_hd__o21a_1 _24226_ (.A1(_07719_),
    .A2(_08324_),
    .B1(_08326_),
    .X(_08327_));
 sky130_fd_sc_hd__o221a_4 _24227_ (.A1(_07158_),
    .A2(_08325_),
    .B1(_07156_),
    .B2(_08325_),
    .C1(_08327_),
    .X(_08328_));
 sky130_fd_sc_hd__buf_2 _24228_ (.A(_08328_),
    .X(_08329_));
 sky130_fd_sc_hd__a2bb2oi_4 _24229_ (.A1_N(_08322_),
    .A2_N(_08329_),
    .B1(_08322_),
    .B2(_08329_),
    .Y(_02651_));
 sky130_fd_sc_hd__o21ai_2 _24230_ (.A1(_08322_),
    .A2(_08329_),
    .B1(_08320_),
    .Y(_08330_));
 sky130_fd_sc_hd__o22a_4 _24231_ (.A1(_08164_),
    .A2(_08165_),
    .B1(_11723_),
    .B2(_08166_),
    .X(_08331_));
 sky130_fd_sc_hd__o22a_1 _24232_ (.A1(_08169_),
    .A2(_08211_),
    .B1(_08168_),
    .B2(_08212_),
    .X(_08332_));
 sky130_fd_sc_hd__o22a_4 _24233_ (.A1(_08190_),
    .A2(_08191_),
    .B1(_08170_),
    .B2(_08192_),
    .X(_08333_));
 sky130_fd_sc_hd__or2_1 _24234_ (.A(_08332_),
    .B(_08333_),
    .X(_08334_));
 sky130_fd_sc_hd__a21bo_1 _24235_ (.A1(_08332_),
    .A2(_08333_),
    .B1_N(_08334_),
    .X(_08335_));
 sky130_fd_sc_hd__o22a_4 _24236_ (.A1(_08208_),
    .A2(_08209_),
    .B1(_08193_),
    .B2(_08210_),
    .X(_08336_));
 sky130_fd_sc_hd__o22a_1 _24237_ (.A1(_08215_),
    .A2(_08248_),
    .B1(_08214_),
    .B2(_08249_),
    .X(_08337_));
 sky130_fd_sc_hd__a21oi_4 _24238_ (.A1(_08174_),
    .A2(_08176_),
    .B1(_08173_),
    .Y(_08338_));
 sky130_fd_sc_hd__or2_1 _24239_ (.A(_06217_),
    .B(_08035_),
    .X(_08339_));
 sky130_fd_sc_hd__clkbuf_2 _24240_ (.A(_11701_),
    .X(_08340_));
 sky130_fd_sc_hd__or2_4 _24241_ (.A(_08340_),
    .B(_05305_),
    .X(_08341_));
 sky130_fd_sc_hd__clkbuf_2 _24242_ (.A(_08341_),
    .X(_08342_));
 sky130_fd_sc_hd__o2bb2a_1 _24243_ (.A1_N(_08339_),
    .A2_N(_08342_),
    .B1(_08339_),
    .B2(_08342_),
    .X(_08343_));
 sky130_vsdinv _24244_ (.A(_08343_),
    .Y(_08344_));
 sky130_fd_sc_hd__or2_1 _24245_ (.A(_07456_),
    .B(_07892_),
    .X(_08345_));
 sky130_fd_sc_hd__a32o_2 _24246_ (.A1(\pcpi_mul.rs2[3] ),
    .A2(_13512_),
    .A3(_08343_),
    .B1(_08344_),
    .B2(_08345_),
    .X(_08346_));
 sky130_fd_sc_hd__buf_1 _24247_ (.A(_08185_),
    .X(_08347_));
 sky130_fd_sc_hd__o22a_1 _24248_ (.A1(_07181_),
    .A2(_08179_),
    .B1(_07183_),
    .B2(_07872_),
    .X(_08348_));
 sky130_fd_sc_hd__and4_1 _24249_ (.A(_13161_),
    .B(_07876_),
    .C(_13167_),
    .D(_08022_),
    .X(_08349_));
 sky130_fd_sc_hd__or2_1 _24250_ (.A(_08348_),
    .B(_08349_),
    .X(_08350_));
 sky130_vsdinv _24251_ (.A(_08350_),
    .Y(_08351_));
 sky130_fd_sc_hd__a22o_1 _24252_ (.A1(_08347_),
    .A2(_08351_),
    .B1(_08184_),
    .B2(_08350_),
    .X(_08352_));
 sky130_fd_sc_hd__clkbuf_2 _24253_ (.A(_08185_),
    .X(_08353_));
 sky130_fd_sc_hd__a21oi_2 _24254_ (.A1(_08183_),
    .A2(_08353_),
    .B1(_08182_),
    .Y(_08354_));
 sky130_fd_sc_hd__a2bb2o_1 _24255_ (.A1_N(_08352_),
    .A2_N(_08354_),
    .B1(_08352_),
    .B2(_08354_),
    .X(_08355_));
 sky130_fd_sc_hd__a2bb2o_1 _24256_ (.A1_N(_08346_),
    .A2_N(_08355_),
    .B1(_08346_),
    .B2(_08355_),
    .X(_08356_));
 sky130_fd_sc_hd__o22a_1 _24257_ (.A1(_08187_),
    .A2(_08188_),
    .B1(_08177_),
    .B2(_08189_),
    .X(_08357_));
 sky130_fd_sc_hd__a2bb2o_1 _24258_ (.A1_N(_08356_),
    .A2_N(_08357_),
    .B1(_08356_),
    .B2(_08357_),
    .X(_08358_));
 sky130_fd_sc_hd__a2bb2o_2 _24259_ (.A1_N(_08338_),
    .A2_N(_08358_),
    .B1(_08338_),
    .B2(_08358_),
    .X(_08359_));
 sky130_fd_sc_hd__o22a_1 _24260_ (.A1(_08197_),
    .A2(_08204_),
    .B1(_08196_),
    .B2(_08205_),
    .X(_08360_));
 sky130_fd_sc_hd__o22a_1 _24261_ (.A1(_08227_),
    .A2(_08228_),
    .B1(_08221_),
    .B2(_08229_),
    .X(_08361_));
 sky130_fd_sc_hd__a21oi_2 _24262_ (.A1(_08202_),
    .A2(_08203_),
    .B1(_08201_),
    .Y(_08362_));
 sky130_fd_sc_hd__o21ba_1 _24263_ (.A1(_08216_),
    .A2(_08220_),
    .B1_N(_08219_),
    .X(_08363_));
 sky130_fd_sc_hd__buf_1 _24264_ (.A(_07324_),
    .X(_08364_));
 sky130_fd_sc_hd__o22a_1 _24265_ (.A1(_08049_),
    .A2(_08198_),
    .B1(_05458_),
    .B2(_08364_),
    .X(_08365_));
 sky130_fd_sc_hd__and4_1 _24266_ (.A(_08052_),
    .B(_07742_),
    .C(_08054_),
    .D(_13528_),
    .X(_08366_));
 sky130_fd_sc_hd__nor2_2 _24267_ (.A(_08365_),
    .B(_08366_),
    .Y(_08367_));
 sky130_fd_sc_hd__nor2_2 _24268_ (.A(_08057_),
    .B(_07464_),
    .Y(_08368_));
 sky130_fd_sc_hd__a2bb2o_1 _24269_ (.A1_N(_08367_),
    .A2_N(_08368_),
    .B1(_08367_),
    .B2(_08368_),
    .X(_08369_));
 sky130_fd_sc_hd__a2bb2o_1 _24270_ (.A1_N(_08363_),
    .A2_N(_08369_),
    .B1(_08363_),
    .B2(_08369_),
    .X(_08370_));
 sky130_fd_sc_hd__a2bb2o_1 _24271_ (.A1_N(_08362_),
    .A2_N(_08370_),
    .B1(_08362_),
    .B2(_08370_),
    .X(_08371_));
 sky130_fd_sc_hd__a2bb2o_1 _24272_ (.A1_N(_08361_),
    .A2_N(_08371_),
    .B1(_08361_),
    .B2(_08371_),
    .X(_08372_));
 sky130_fd_sc_hd__a2bb2o_1 _24273_ (.A1_N(_08360_),
    .A2_N(_08372_),
    .B1(_08360_),
    .B2(_08372_),
    .X(_08373_));
 sky130_fd_sc_hd__o22a_1 _24274_ (.A1(_08195_),
    .A2(_08206_),
    .B1(_08194_),
    .B2(_08207_),
    .X(_08374_));
 sky130_fd_sc_hd__a2bb2o_1 _24275_ (.A1_N(_08373_),
    .A2_N(_08374_),
    .B1(_08373_),
    .B2(_08374_),
    .X(_08375_));
 sky130_fd_sc_hd__a2bb2o_2 _24276_ (.A1_N(_08359_),
    .A2_N(_08375_),
    .B1(_08359_),
    .B2(_08375_),
    .X(_08376_));
 sky130_fd_sc_hd__a2bb2o_1 _24277_ (.A1_N(_08337_),
    .A2_N(_08376_),
    .B1(_08337_),
    .B2(_08376_),
    .X(_08377_));
 sky130_fd_sc_hd__a2bb2o_1 _24278_ (.A1_N(_08336_),
    .A2_N(_08377_),
    .B1(_08336_),
    .B2(_08377_),
    .X(_08378_));
 sky130_fd_sc_hd__o22a_1 _24279_ (.A1(_08245_),
    .A2(_08246_),
    .B1(_08230_),
    .B2(_08247_),
    .X(_08379_));
 sky130_fd_sc_hd__o22a_1 _24280_ (.A1(_08252_),
    .A2(_08271_),
    .B1(_08251_),
    .B2(_08272_),
    .X(_08380_));
 sky130_fd_sc_hd__or2_1 _24281_ (.A(_05537_),
    .B(_07172_),
    .X(_08381_));
 sky130_fd_sc_hd__o22a_1 _24282_ (.A1(_08217_),
    .A2(_07905_),
    .B1(_05588_),
    .B2(_07018_),
    .X(_08382_));
 sky130_fd_sc_hd__and4_1 _24283_ (.A(_07363_),
    .B(_07907_),
    .C(_07364_),
    .D(_13541_),
    .X(_08383_));
 sky130_fd_sc_hd__or2_1 _24284_ (.A(_08382_),
    .B(_08383_),
    .X(_08384_));
 sky130_fd_sc_hd__a2bb2o_1 _24285_ (.A1_N(_08381_),
    .A2_N(_08384_),
    .B1(_08381_),
    .B2(_08384_),
    .X(_08385_));
 sky130_fd_sc_hd__clkbuf_2 _24286_ (.A(_05794_),
    .X(_08386_));
 sky130_fd_sc_hd__or2_1 _24287_ (.A(_08386_),
    .B(_07482_),
    .X(_08387_));
 sky130_fd_sc_hd__clkbuf_2 _24288_ (.A(_06573_),
    .X(_08388_));
 sky130_fd_sc_hd__o22a_1 _24289_ (.A1(_08223_),
    .A2(_07348_),
    .B1(_07930_),
    .B2(_08388_),
    .X(_08389_));
 sky130_fd_sc_hd__buf_1 _24290_ (.A(_06535_),
    .X(_08390_));
 sky130_fd_sc_hd__buf_1 _24291_ (.A(_06536_),
    .X(_08391_));
 sky130_fd_sc_hd__and4_1 _24292_ (.A(_08390_),
    .B(_07485_),
    .C(_08391_),
    .D(_13552_),
    .X(_08392_));
 sky130_fd_sc_hd__or2_1 _24293_ (.A(_08389_),
    .B(_08392_),
    .X(_08393_));
 sky130_fd_sc_hd__a2bb2o_1 _24294_ (.A1_N(_08387_),
    .A2_N(_08393_),
    .B1(_08387_),
    .B2(_08393_),
    .X(_08394_));
 sky130_fd_sc_hd__o21ba_1 _24295_ (.A1(_08222_),
    .A2(_08226_),
    .B1_N(_08225_),
    .X(_08395_));
 sky130_fd_sc_hd__a2bb2o_1 _24296_ (.A1_N(_08394_),
    .A2_N(_08395_),
    .B1(_08394_),
    .B2(_08395_),
    .X(_08396_));
 sky130_fd_sc_hd__a2bb2o_2 _24297_ (.A1_N(_08385_),
    .A2_N(_08396_),
    .B1(_08385_),
    .B2(_08396_),
    .X(_08397_));
 sky130_fd_sc_hd__a21oi_2 _24298_ (.A1(_08240_),
    .A2(_08242_),
    .B1(_08239_),
    .Y(_08398_));
 sky130_fd_sc_hd__o21ba_1 _24299_ (.A1(_08254_),
    .A2(_08258_),
    .B1_N(_08257_),
    .X(_08399_));
 sky130_fd_sc_hd__or2_1 _24300_ (.A(_08241_),
    .B(_06438_),
    .X(_08400_));
 sky130_fd_sc_hd__buf_2 _24301_ (.A(_06088_),
    .X(_08401_));
 sky130_fd_sc_hd__o22a_1 _24302_ (.A1(_07941_),
    .A2(_06921_),
    .B1(_08401_),
    .B2(_06329_),
    .X(_08402_));
 sky130_fd_sc_hd__and4_1 _24303_ (.A(_13118_),
    .B(_06925_),
    .C(_13122_),
    .D(_07059_),
    .X(_08403_));
 sky130_fd_sc_hd__or2_1 _24304_ (.A(_08402_),
    .B(_08403_),
    .X(_08404_));
 sky130_fd_sc_hd__a2bb2o_1 _24305_ (.A1_N(_08400_),
    .A2_N(_08404_),
    .B1(_08400_),
    .B2(_08404_),
    .X(_08405_));
 sky130_fd_sc_hd__a2bb2o_1 _24306_ (.A1_N(_08399_),
    .A2_N(_08405_),
    .B1(_08399_),
    .B2(_08405_),
    .X(_08406_));
 sky130_fd_sc_hd__a2bb2o_1 _24307_ (.A1_N(_08398_),
    .A2_N(_08406_),
    .B1(_08398_),
    .B2(_08406_),
    .X(_08407_));
 sky130_fd_sc_hd__o22a_1 _24308_ (.A1(_08232_),
    .A2(_08243_),
    .B1(_08231_),
    .B2(_08244_),
    .X(_08408_));
 sky130_fd_sc_hd__a2bb2o_1 _24309_ (.A1_N(_08407_),
    .A2_N(_08408_),
    .B1(_08407_),
    .B2(_08408_),
    .X(_08409_));
 sky130_fd_sc_hd__a2bb2o_1 _24310_ (.A1_N(_08397_),
    .A2_N(_08409_),
    .B1(_08397_),
    .B2(_08409_),
    .X(_08410_));
 sky130_fd_sc_hd__a2bb2o_1 _24311_ (.A1_N(_08380_),
    .A2_N(_08410_),
    .B1(_08380_),
    .B2(_08410_),
    .X(_08411_));
 sky130_fd_sc_hd__a2bb2o_1 _24312_ (.A1_N(_08379_),
    .A2_N(_08411_),
    .B1(_08379_),
    .B2(_08411_),
    .X(_08412_));
 sky130_fd_sc_hd__o22a_1 _24313_ (.A1(_08268_),
    .A2(_08269_),
    .B1(_08259_),
    .B2(_08270_),
    .X(_08413_));
 sky130_fd_sc_hd__o22a_1 _24314_ (.A1(_08275_),
    .A2(_08280_),
    .B1(_08274_),
    .B2(_08281_),
    .X(_08414_));
 sky130_fd_sc_hd__or2_1 _24315_ (.A(_08253_),
    .B(_06132_),
    .X(_08415_));
 sky130_fd_sc_hd__clkbuf_2 _24316_ (.A(_07081_),
    .X(_08416_));
 sky130_fd_sc_hd__buf_1 _24317_ (.A(_06030_),
    .X(_08417_));
 sky130_fd_sc_hd__o22a_1 _24318_ (.A1(_08416_),
    .A2(_06028_),
    .B1(_06390_),
    .B2(_08417_),
    .X(_08418_));
 sky130_fd_sc_hd__buf_1 _24319_ (.A(_13574_),
    .X(_08419_));
 sky130_fd_sc_hd__and4_1 _24320_ (.A(_08256_),
    .B(_13579_),
    .C(_08102_),
    .D(_08419_),
    .X(_08420_));
 sky130_fd_sc_hd__or2_1 _24321_ (.A(_08418_),
    .B(_08420_),
    .X(_08421_));
 sky130_fd_sc_hd__a2bb2o_1 _24322_ (.A1_N(_08415_),
    .A2_N(_08421_),
    .B1(_08415_),
    .B2(_08421_),
    .X(_08422_));
 sky130_fd_sc_hd__or2_1 _24323_ (.A(_06688_),
    .B(_05928_),
    .X(_08423_));
 sky130_fd_sc_hd__clkbuf_2 _24324_ (.A(_06805_),
    .X(_08424_));
 sky130_fd_sc_hd__buf_1 _24325_ (.A(_05724_),
    .X(_08425_));
 sky130_fd_sc_hd__o22a_1 _24326_ (.A1(_08262_),
    .A2(_08263_),
    .B1(_08424_),
    .B2(_08425_),
    .X(_08426_));
 sky130_fd_sc_hd__buf_1 _24327_ (.A(_13584_),
    .X(_08427_));
 sky130_fd_sc_hd__and4_1 _24328_ (.A(_13097_),
    .B(_08265_),
    .C(_13102_),
    .D(_08427_),
    .X(_08428_));
 sky130_fd_sc_hd__or2_1 _24329_ (.A(_08426_),
    .B(_08428_),
    .X(_08429_));
 sky130_fd_sc_hd__a2bb2o_1 _24330_ (.A1_N(_08423_),
    .A2_N(_08429_),
    .B1(_08423_),
    .B2(_08429_),
    .X(_08430_));
 sky130_fd_sc_hd__o21ba_1 _24331_ (.A1(_08260_),
    .A2(_08267_),
    .B1_N(_08266_),
    .X(_08431_));
 sky130_fd_sc_hd__a2bb2o_1 _24332_ (.A1_N(_08430_),
    .A2_N(_08431_),
    .B1(_08430_),
    .B2(_08431_),
    .X(_08432_));
 sky130_fd_sc_hd__a2bb2o_1 _24333_ (.A1_N(_08422_),
    .A2_N(_08432_),
    .B1(_08422_),
    .B2(_08432_),
    .X(_08433_));
 sky130_fd_sc_hd__a2bb2o_1 _24334_ (.A1_N(_08414_),
    .A2_N(_08433_),
    .B1(_08414_),
    .B2(_08433_),
    .X(_08434_));
 sky130_fd_sc_hd__a2bb2o_1 _24335_ (.A1_N(_08413_),
    .A2_N(_08434_),
    .B1(_08413_),
    .B2(_08434_),
    .X(_08435_));
 sky130_fd_sc_hd__o21ba_1 _24336_ (.A1(_08276_),
    .A2(_08279_),
    .B1_N(_08278_),
    .X(_08436_));
 sky130_fd_sc_hd__o21ba_1 _24337_ (.A1(_08284_),
    .A2(_08290_),
    .B1_N(_08289_),
    .X(_08437_));
 sky130_fd_sc_hd__or2_1 _24338_ (.A(_08118_),
    .B(_05731_),
    .X(_08438_));
 sky130_fd_sc_hd__buf_1 _24339_ (.A(_06831_),
    .X(_08439_));
 sky130_fd_sc_hd__o22a_1 _24340_ (.A1(_08120_),
    .A2(_06099_),
    .B1(_08121_),
    .B2(_08439_),
    .X(_08440_));
 sky130_fd_sc_hd__buf_1 _24341_ (.A(_13091_),
    .X(_08441_));
 sky130_fd_sc_hd__and4_1 _24342_ (.A(_08123_),
    .B(_13599_),
    .C(_08441_),
    .D(_13595_),
    .X(_08442_));
 sky130_fd_sc_hd__or2_1 _24343_ (.A(_08440_),
    .B(_08442_),
    .X(_08443_));
 sky130_fd_sc_hd__a2bb2o_1 _24344_ (.A1_N(_08438_),
    .A2_N(_08443_),
    .B1(_08438_),
    .B2(_08443_),
    .X(_08444_));
 sky130_fd_sc_hd__a2bb2o_1 _24345_ (.A1_N(_08437_),
    .A2_N(_08444_),
    .B1(_08437_),
    .B2(_08444_),
    .X(_08445_));
 sky130_fd_sc_hd__a2bb2o_1 _24346_ (.A1_N(_08436_),
    .A2_N(_08445_),
    .B1(_08436_),
    .B2(_08445_),
    .X(_08446_));
 sky130_fd_sc_hd__or2_1 _24347_ (.A(_07681_),
    .B(_07079_),
    .X(_08447_));
 sky130_fd_sc_hd__buf_1 _24348_ (.A(_08285_),
    .X(_08448_));
 sky130_fd_sc_hd__buf_1 _24349_ (.A(_07678_),
    .X(_08449_));
 sky130_fd_sc_hd__o22a_1 _24350_ (.A1(_08448_),
    .A2(_08136_),
    .B1(_08449_),
    .B2(_08283_),
    .X(_08450_));
 sky130_fd_sc_hd__buf_1 _24351_ (.A(_13072_),
    .X(_08451_));
 sky130_fd_sc_hd__buf_1 _24352_ (.A(_07830_),
    .X(_08452_));
 sky130_fd_sc_hd__and4_1 _24353_ (.A(_08451_),
    .B(_13613_),
    .C(_08452_),
    .D(_13609_),
    .X(_08453_));
 sky130_fd_sc_hd__or2_1 _24354_ (.A(_08450_),
    .B(_08453_),
    .X(_08454_));
 sky130_fd_sc_hd__a2bb2o_1 _24355_ (.A1_N(_08447_),
    .A2_N(_08454_),
    .B1(_08447_),
    .B2(_08454_),
    .X(_08455_));
 sky130_fd_sc_hd__or2_1 _24356_ (.A(_08292_),
    .B(_05340_),
    .X(_08456_));
 sky130_fd_sc_hd__buf_1 _24357_ (.A(\pcpi_mul.rs2[31] ),
    .X(_08457_));
 sky130_fd_sc_hd__and4_1 _24358_ (.A(_08295_),
    .B(_05910_),
    .C(_08457_),
    .D(_13620_),
    .X(_08458_));
 sky130_fd_sc_hd__o22a_1 _24359_ (.A1(_11717_),
    .A2(_13624_),
    .B1(_08131_),
    .B2(_05315_),
    .X(_08459_));
 sky130_fd_sc_hd__or2_1 _24360_ (.A(_08458_),
    .B(_08459_),
    .X(_08460_));
 sky130_fd_sc_hd__a2bb2o_1 _24361_ (.A1_N(_08456_),
    .A2_N(_08460_),
    .B1(_08456_),
    .B2(_08460_),
    .X(_08461_));
 sky130_fd_sc_hd__o21ba_1 _24362_ (.A1(_08293_),
    .A2(_08298_),
    .B1_N(_08296_),
    .X(_08462_));
 sky130_fd_sc_hd__a2bb2o_1 _24363_ (.A1_N(_08461_),
    .A2_N(_08462_),
    .B1(_08461_),
    .B2(_08462_),
    .X(_08463_));
 sky130_fd_sc_hd__a2bb2o_1 _24364_ (.A1_N(_08455_),
    .A2_N(_08463_),
    .B1(_08455_),
    .B2(_08463_),
    .X(_08464_));
 sky130_fd_sc_hd__o22a_1 _24365_ (.A1(_08134_),
    .A2(_08299_),
    .B1(_08291_),
    .B2(_08300_),
    .X(_08465_));
 sky130_fd_sc_hd__a2bb2o_1 _24366_ (.A1_N(_08464_),
    .A2_N(_08465_),
    .B1(_08464_),
    .B2(_08465_),
    .X(_08466_));
 sky130_fd_sc_hd__a2bb2o_1 _24367_ (.A1_N(_08446_),
    .A2_N(_08466_),
    .B1(_08446_),
    .B2(_08466_),
    .X(_08467_));
 sky130_fd_sc_hd__o22a_1 _24368_ (.A1(_08142_),
    .A2(_08301_),
    .B1(_08282_),
    .B2(_08302_),
    .X(_08468_));
 sky130_fd_sc_hd__a2bb2o_1 _24369_ (.A1_N(_08467_),
    .A2_N(_08468_),
    .B1(_08467_),
    .B2(_08468_),
    .X(_08469_));
 sky130_fd_sc_hd__a2bb2o_1 _24370_ (.A1_N(_08435_),
    .A2_N(_08469_),
    .B1(_08435_),
    .B2(_08469_),
    .X(_08470_));
 sky130_fd_sc_hd__o22a_1 _24371_ (.A1(_08303_),
    .A2(_08304_),
    .B1(_08273_),
    .B2(_08305_),
    .X(_08471_));
 sky130_fd_sc_hd__a2bb2o_1 _24372_ (.A1_N(_08470_),
    .A2_N(_08471_),
    .B1(_08470_),
    .B2(_08471_),
    .X(_08472_));
 sky130_fd_sc_hd__a2bb2o_1 _24373_ (.A1_N(_08412_),
    .A2_N(_08472_),
    .B1(_08412_),
    .B2(_08472_),
    .X(_08473_));
 sky130_fd_sc_hd__o22a_1 _24374_ (.A1(_08306_),
    .A2(_08307_),
    .B1(_08250_),
    .B2(_08308_),
    .X(_08474_));
 sky130_fd_sc_hd__a2bb2o_1 _24375_ (.A1_N(_08473_),
    .A2_N(_08474_),
    .B1(_08473_),
    .B2(_08474_),
    .X(_08475_));
 sky130_fd_sc_hd__a2bb2o_1 _24376_ (.A1_N(_08378_),
    .A2_N(_08475_),
    .B1(_08378_),
    .B2(_08475_),
    .X(_08476_));
 sky130_fd_sc_hd__o22a_1 _24377_ (.A1(_08309_),
    .A2(_08310_),
    .B1(_08213_),
    .B2(_08311_),
    .X(_08477_));
 sky130_fd_sc_hd__a2bb2o_1 _24378_ (.A1_N(_08476_),
    .A2_N(_08477_),
    .B1(_08476_),
    .B2(_08477_),
    .X(_08478_));
 sky130_fd_sc_hd__a2bb2o_1 _24379_ (.A1_N(_08335_),
    .A2_N(_08478_),
    .B1(_08335_),
    .B2(_08478_),
    .X(_08479_));
 sky130_fd_sc_hd__o22a_1 _24380_ (.A1(_08312_),
    .A2(_08313_),
    .B1(_08167_),
    .B2(_08314_),
    .X(_08480_));
 sky130_fd_sc_hd__a2bb2o_1 _24381_ (.A1_N(_08479_),
    .A2_N(_08480_),
    .B1(_08479_),
    .B2(_08480_),
    .X(_08481_));
 sky130_fd_sc_hd__a2bb2o_1 _24382_ (.A1_N(_08331_),
    .A2_N(_08481_),
    .B1(_08331_),
    .B2(_08481_),
    .X(_08482_));
 sky130_fd_sc_hd__o22a_1 _24383_ (.A1(_08315_),
    .A2(_08316_),
    .B1(_08015_),
    .B2(_08317_),
    .X(_08483_));
 sky130_fd_sc_hd__or2_1 _24384_ (.A(_08482_),
    .B(_08483_),
    .X(_08484_));
 sky130_fd_sc_hd__a21bo_1 _24385_ (.A1(_08482_),
    .A2(_08483_),
    .B1_N(_08484_),
    .X(_08485_));
 sky130_fd_sc_hd__a2bb2o_4 _24386_ (.A1_N(_08330_),
    .A2_N(_08485_),
    .B1(_08330_),
    .B2(_08485_),
    .X(_02652_));
 sky130_fd_sc_hd__o22a_1 _24387_ (.A1(_08337_),
    .A2(_08376_),
    .B1(_08336_),
    .B2(_08377_),
    .X(_08486_));
 sky130_fd_sc_hd__o22a_4 _24388_ (.A1(_08356_),
    .A2(_08357_),
    .B1(_08338_),
    .B2(_08358_),
    .X(_08487_));
 sky130_fd_sc_hd__or2_1 _24389_ (.A(_08486_),
    .B(_08487_),
    .X(_08488_));
 sky130_fd_sc_hd__a21bo_1 _24390_ (.A1(_08486_),
    .A2(_08487_),
    .B1_N(_08488_),
    .X(_08489_));
 sky130_fd_sc_hd__o22a_2 _24391_ (.A1(_08373_),
    .A2(_08374_),
    .B1(_08359_),
    .B2(_08375_),
    .X(_08490_));
 sky130_fd_sc_hd__o22a_1 _24392_ (.A1(_08380_),
    .A2(_08410_),
    .B1(_08379_),
    .B2(_08411_),
    .X(_08491_));
 sky130_fd_sc_hd__o22a_2 _24393_ (.A1(_08339_),
    .A2(_08342_),
    .B1(_08344_),
    .B2(_08345_),
    .X(_08492_));
 sky130_fd_sc_hd__or2_4 _24394_ (.A(_08340_),
    .B(_05322_),
    .X(_08493_));
 sky130_fd_sc_hd__nor2_8 _24395_ (.A(_08341_),
    .B(_08493_),
    .Y(_08494_));
 sky130_fd_sc_hd__a21oi_4 _24396_ (.A1(_08342_),
    .A2(_08493_),
    .B1(_08494_),
    .Y(_08495_));
 sky130_fd_sc_hd__buf_1 _24397_ (.A(_08495_),
    .X(_08496_));
 sky130_fd_sc_hd__clkbuf_2 _24398_ (.A(_08033_),
    .X(_08497_));
 sky130_fd_sc_hd__clkbuf_2 _24399_ (.A(_08497_),
    .X(_08498_));
 sky130_fd_sc_hd__buf_1 _24400_ (.A(_08498_),
    .X(_08499_));
 sky130_fd_sc_hd__clkbuf_4 _24401_ (.A(_08499_),
    .X(_08500_));
 sky130_fd_sc_hd__nor2_4 _24402_ (.A(_06887_),
    .B(_08500_),
    .Y(_08501_));
 sky130_fd_sc_hd__a2bb2o_1 _24403_ (.A1_N(_08496_),
    .A2_N(_08501_),
    .B1(_08496_),
    .B2(_08501_),
    .X(_08502_));
 sky130_fd_sc_hd__o22a_1 _24404_ (.A1(_07181_),
    .A2(_07872_),
    .B1(_07183_),
    .B2(_07890_),
    .X(_08503_));
 sky130_fd_sc_hd__and4_1 _24405_ (.A(_13161_),
    .B(_08022_),
    .C(_13167_),
    .D(_13509_),
    .X(_08504_));
 sky130_fd_sc_hd__or2_1 _24406_ (.A(_08503_),
    .B(_08504_),
    .X(_08505_));
 sky130_vsdinv _24407_ (.A(_08505_),
    .Y(_08506_));
 sky130_fd_sc_hd__a22o_1 _24408_ (.A1(_08186_),
    .A2(_08506_),
    .B1(_08184_),
    .B2(_08505_),
    .X(_08507_));
 sky130_fd_sc_hd__a21oi_2 _24409_ (.A1(_08353_),
    .A2(_08351_),
    .B1(_08349_),
    .Y(_08508_));
 sky130_fd_sc_hd__a2bb2o_1 _24410_ (.A1_N(_08507_),
    .A2_N(_08508_),
    .B1(_08507_),
    .B2(_08508_),
    .X(_08509_));
 sky130_fd_sc_hd__a2bb2o_1 _24411_ (.A1_N(_08502_),
    .A2_N(_08509_),
    .B1(_08502_),
    .B2(_08509_),
    .X(_08510_));
 sky130_fd_sc_hd__o22a_1 _24412_ (.A1(_08352_),
    .A2(_08354_),
    .B1(_08346_),
    .B2(_08355_),
    .X(_08511_));
 sky130_fd_sc_hd__a2bb2o_1 _24413_ (.A1_N(_08510_),
    .A2_N(_08511_),
    .B1(_08510_),
    .B2(_08511_),
    .X(_08512_));
 sky130_fd_sc_hd__a2bb2o_2 _24414_ (.A1_N(_08492_),
    .A2_N(_08512_),
    .B1(_08492_),
    .B2(_08512_),
    .X(_08513_));
 sky130_fd_sc_hd__o22a_1 _24415_ (.A1(_08363_),
    .A2(_08369_),
    .B1(_08362_),
    .B2(_08370_),
    .X(_08514_));
 sky130_fd_sc_hd__o22a_1 _24416_ (.A1(_08394_),
    .A2(_08395_),
    .B1(_08385_),
    .B2(_08396_),
    .X(_08515_));
 sky130_fd_sc_hd__a21oi_2 _24417_ (.A1(_08367_),
    .A2(_08368_),
    .B1(_08366_),
    .Y(_08516_));
 sky130_fd_sc_hd__o21ba_1 _24418_ (.A1(_08381_),
    .A2(_08384_),
    .B1_N(_08383_),
    .X(_08517_));
 sky130_fd_sc_hd__clkbuf_2 _24419_ (.A(_05457_),
    .X(_08518_));
 sky130_fd_sc_hd__o22a_1 _24420_ (.A1(_08049_),
    .A2(_08364_),
    .B1(_08518_),
    .B2(_07463_),
    .X(_08519_));
 sky130_fd_sc_hd__and4_1 _24421_ (.A(_08052_),
    .B(_13528_),
    .C(_08054_),
    .D(_07587_),
    .X(_08520_));
 sky130_fd_sc_hd__nor2_2 _24422_ (.A(_08519_),
    .B(_08520_),
    .Y(_08521_));
 sky130_fd_sc_hd__nor2_2 _24423_ (.A(_08057_),
    .B(_07596_),
    .Y(_08522_));
 sky130_fd_sc_hd__a2bb2o_1 _24424_ (.A1_N(_08521_),
    .A2_N(_08522_),
    .B1(_08521_),
    .B2(_08522_),
    .X(_08523_));
 sky130_fd_sc_hd__a2bb2o_1 _24425_ (.A1_N(_08517_),
    .A2_N(_08523_),
    .B1(_08517_),
    .B2(_08523_),
    .X(_08524_));
 sky130_fd_sc_hd__a2bb2o_1 _24426_ (.A1_N(_08516_),
    .A2_N(_08524_),
    .B1(_08516_),
    .B2(_08524_),
    .X(_08525_));
 sky130_fd_sc_hd__a2bb2o_1 _24427_ (.A1_N(_08515_),
    .A2_N(_08525_),
    .B1(_08515_),
    .B2(_08525_),
    .X(_08526_));
 sky130_fd_sc_hd__a2bb2o_1 _24428_ (.A1_N(_08514_),
    .A2_N(_08526_),
    .B1(_08514_),
    .B2(_08526_),
    .X(_08527_));
 sky130_fd_sc_hd__o22a_1 _24429_ (.A1(_08361_),
    .A2(_08371_),
    .B1(_08360_),
    .B2(_08372_),
    .X(_08528_));
 sky130_fd_sc_hd__a2bb2o_1 _24430_ (.A1_N(_08527_),
    .A2_N(_08528_),
    .B1(_08527_),
    .B2(_08528_),
    .X(_08529_));
 sky130_fd_sc_hd__a2bb2o_2 _24431_ (.A1_N(_08513_),
    .A2_N(_08529_),
    .B1(_08513_),
    .B2(_08529_),
    .X(_08530_));
 sky130_fd_sc_hd__a2bb2o_1 _24432_ (.A1_N(_08491_),
    .A2_N(_08530_),
    .B1(_08491_),
    .B2(_08530_),
    .X(_08531_));
 sky130_fd_sc_hd__a2bb2o_1 _24433_ (.A1_N(_08490_),
    .A2_N(_08531_),
    .B1(_08490_),
    .B2(_08531_),
    .X(_08532_));
 sky130_fd_sc_hd__o22a_1 _24434_ (.A1(_08407_),
    .A2(_08408_),
    .B1(_08397_),
    .B2(_08409_),
    .X(_08533_));
 sky130_fd_sc_hd__o22a_1 _24435_ (.A1(_08414_),
    .A2(_08433_),
    .B1(_08413_),
    .B2(_08434_),
    .X(_08534_));
 sky130_fd_sc_hd__clkbuf_4 _24436_ (.A(_05711_),
    .X(_08535_));
 sky130_fd_sc_hd__or2_1 _24437_ (.A(_08535_),
    .B(_07197_),
    .X(_08536_));
 sky130_fd_sc_hd__clkbuf_2 _24438_ (.A(_06300_),
    .X(_08537_));
 sky130_fd_sc_hd__clkbuf_2 _24439_ (.A(_05592_),
    .X(_08538_));
 sky130_fd_sc_hd__o22a_1 _24440_ (.A1(_08537_),
    .A2(_08050_),
    .B1(_08538_),
    .B2(_07457_),
    .X(_08539_));
 sky130_fd_sc_hd__and4_1 _24441_ (.A(_13137_),
    .B(_07908_),
    .C(_13143_),
    .D(_08200_),
    .X(_08540_));
 sky130_fd_sc_hd__or2_1 _24442_ (.A(_08539_),
    .B(_08540_),
    .X(_08541_));
 sky130_fd_sc_hd__a2bb2o_1 _24443_ (.A1_N(_08536_),
    .A2_N(_08541_),
    .B1(_08536_),
    .B2(_08541_),
    .X(_08542_));
 sky130_fd_sc_hd__or2_1 _24444_ (.A(_08386_),
    .B(_06881_),
    .X(_08543_));
 sky130_fd_sc_hd__clkbuf_2 _24445_ (.A(_06710_),
    .X(_08544_));
 sky130_fd_sc_hd__buf_1 _24446_ (.A(_06533_),
    .X(_08545_));
 sky130_fd_sc_hd__o22a_1 _24447_ (.A1(_08544_),
    .A2(_08388_),
    .B1(_08545_),
    .B2(_07762_),
    .X(_08546_));
 sky130_fd_sc_hd__buf_1 _24448_ (.A(_06535_),
    .X(_08547_));
 sky130_fd_sc_hd__buf_1 _24449_ (.A(_06536_),
    .X(_08548_));
 sky130_fd_sc_hd__and4_1 _24450_ (.A(_08547_),
    .B(_07187_),
    .C(_08548_),
    .D(_13549_),
    .X(_08549_));
 sky130_fd_sc_hd__or2_1 _24451_ (.A(_08546_),
    .B(_08549_),
    .X(_08550_));
 sky130_fd_sc_hd__a2bb2o_1 _24452_ (.A1_N(_08543_),
    .A2_N(_08550_),
    .B1(_08543_),
    .B2(_08550_),
    .X(_08551_));
 sky130_fd_sc_hd__o21ba_1 _24453_ (.A1(_08387_),
    .A2(_08393_),
    .B1_N(_08392_),
    .X(_08552_));
 sky130_fd_sc_hd__a2bb2o_1 _24454_ (.A1_N(_08551_),
    .A2_N(_08552_),
    .B1(_08551_),
    .B2(_08552_),
    .X(_08553_));
 sky130_fd_sc_hd__a2bb2o_2 _24455_ (.A1_N(_08542_),
    .A2_N(_08553_),
    .B1(_08542_),
    .B2(_08553_),
    .X(_08554_));
 sky130_fd_sc_hd__o21ba_1 _24456_ (.A1(_08400_),
    .A2(_08404_),
    .B1_N(_08403_),
    .X(_08555_));
 sky130_fd_sc_hd__o21ba_1 _24457_ (.A1(_08415_),
    .A2(_08421_),
    .B1_N(_08420_),
    .X(_08556_));
 sky130_fd_sc_hd__buf_2 _24458_ (.A(_07348_),
    .X(_08557_));
 sky130_fd_sc_hd__or2_1 _24459_ (.A(_08241_),
    .B(_08557_),
    .X(_08558_));
 sky130_fd_sc_hd__buf_1 _24460_ (.A(_06765_),
    .X(_08559_));
 sky130_fd_sc_hd__o22a_1 _24461_ (.A1(_08233_),
    .A2(_06329_),
    .B1(_08401_),
    .B2(_08559_),
    .X(_08560_));
 sky130_fd_sc_hd__and4_1 _24462_ (.A(_08236_),
    .B(_13564_),
    .C(_08238_),
    .D(_13560_),
    .X(_08561_));
 sky130_fd_sc_hd__or2_1 _24463_ (.A(_08560_),
    .B(_08561_),
    .X(_08562_));
 sky130_fd_sc_hd__a2bb2o_1 _24464_ (.A1_N(_08558_),
    .A2_N(_08562_),
    .B1(_08558_),
    .B2(_08562_),
    .X(_08563_));
 sky130_fd_sc_hd__a2bb2o_1 _24465_ (.A1_N(_08556_),
    .A2_N(_08563_),
    .B1(_08556_),
    .B2(_08563_),
    .X(_08564_));
 sky130_fd_sc_hd__a2bb2o_1 _24466_ (.A1_N(_08555_),
    .A2_N(_08564_),
    .B1(_08555_),
    .B2(_08564_),
    .X(_08565_));
 sky130_fd_sc_hd__o22a_1 _24467_ (.A1(_08399_),
    .A2(_08405_),
    .B1(_08398_),
    .B2(_08406_),
    .X(_08566_));
 sky130_fd_sc_hd__a2bb2o_1 _24468_ (.A1_N(_08565_),
    .A2_N(_08566_),
    .B1(_08565_),
    .B2(_08566_),
    .X(_08567_));
 sky130_fd_sc_hd__a2bb2o_1 _24469_ (.A1_N(_08554_),
    .A2_N(_08567_),
    .B1(_08554_),
    .B2(_08567_),
    .X(_08568_));
 sky130_fd_sc_hd__a2bb2o_1 _24470_ (.A1_N(_08534_),
    .A2_N(_08568_),
    .B1(_08534_),
    .B2(_08568_),
    .X(_08569_));
 sky130_fd_sc_hd__a2bb2o_1 _24471_ (.A1_N(_08533_),
    .A2_N(_08569_),
    .B1(_08533_),
    .B2(_08569_),
    .X(_08570_));
 sky130_fd_sc_hd__o22a_1 _24472_ (.A1(_08430_),
    .A2(_08431_),
    .B1(_08422_),
    .B2(_08432_),
    .X(_08571_));
 sky130_fd_sc_hd__o22a_1 _24473_ (.A1(_08437_),
    .A2(_08444_),
    .B1(_08436_),
    .B2(_08445_),
    .X(_08572_));
 sky130_fd_sc_hd__or2_1 _24474_ (.A(_06285_),
    .B(_06327_),
    .X(_08573_));
 sky130_fd_sc_hd__buf_1 _24475_ (.A(_07081_),
    .X(_08574_));
 sky130_fd_sc_hd__clkbuf_2 _24476_ (.A(_06389_),
    .X(_08575_));
 sky130_fd_sc_hd__o22a_1 _24477_ (.A1(_08574_),
    .A2(_06031_),
    .B1(_08575_),
    .B2(_08234_),
    .X(_08576_));
 sky130_fd_sc_hd__buf_1 _24478_ (.A(_13105_),
    .X(_08577_));
 sky130_fd_sc_hd__buf_1 _24479_ (.A(_06941_),
    .X(_08578_));
 sky130_fd_sc_hd__and4_1 _24480_ (.A(_08577_),
    .B(_08419_),
    .C(_08578_),
    .D(_13570_),
    .X(_08579_));
 sky130_fd_sc_hd__or2_1 _24481_ (.A(_08576_),
    .B(_08579_),
    .X(_08580_));
 sky130_fd_sc_hd__a2bb2o_2 _24482_ (.A1_N(_08573_),
    .A2_N(_08580_),
    .B1(_08573_),
    .B2(_08580_),
    .X(_08581_));
 sky130_fd_sc_hd__buf_1 _24483_ (.A(_07663_),
    .X(_08582_));
 sky130_fd_sc_hd__or2_1 _24484_ (.A(_08582_),
    .B(_05932_),
    .X(_08583_));
 sky130_fd_sc_hd__o22a_1 _24485_ (.A1(_08262_),
    .A2(_08425_),
    .B1(_08424_),
    .B2(_05820_),
    .X(_08584_));
 sky130_fd_sc_hd__buf_1 _24486_ (.A(_13096_),
    .X(_08585_));
 sky130_fd_sc_hd__buf_1 _24487_ (.A(_13101_),
    .X(_08586_));
 sky130_fd_sc_hd__buf_1 _24488_ (.A(_13581_),
    .X(_08587_));
 sky130_fd_sc_hd__and4_1 _24489_ (.A(_08585_),
    .B(_08427_),
    .C(_08586_),
    .D(_08587_),
    .X(_08588_));
 sky130_fd_sc_hd__or2_1 _24490_ (.A(_08584_),
    .B(_08588_),
    .X(_08589_));
 sky130_fd_sc_hd__a2bb2o_1 _24491_ (.A1_N(_08583_),
    .A2_N(_08589_),
    .B1(_08583_),
    .B2(_08589_),
    .X(_08590_));
 sky130_fd_sc_hd__o21ba_1 _24492_ (.A1(_08423_),
    .A2(_08429_),
    .B1_N(_08428_),
    .X(_08591_));
 sky130_fd_sc_hd__a2bb2o_1 _24493_ (.A1_N(_08590_),
    .A2_N(_08591_),
    .B1(_08590_),
    .B2(_08591_),
    .X(_08592_));
 sky130_fd_sc_hd__a2bb2o_1 _24494_ (.A1_N(_08581_),
    .A2_N(_08592_),
    .B1(_08581_),
    .B2(_08592_),
    .X(_08593_));
 sky130_fd_sc_hd__a2bb2o_1 _24495_ (.A1_N(_08572_),
    .A2_N(_08593_),
    .B1(_08572_),
    .B2(_08593_),
    .X(_08594_));
 sky130_fd_sc_hd__a2bb2o_1 _24496_ (.A1_N(_08571_),
    .A2_N(_08594_),
    .B1(_08571_),
    .B2(_08594_),
    .X(_08595_));
 sky130_fd_sc_hd__o21ba_1 _24497_ (.A1(_08438_),
    .A2(_08443_),
    .B1_N(_08442_),
    .X(_08596_));
 sky130_fd_sc_hd__o21ba_1 _24498_ (.A1(_08447_),
    .A2(_08454_),
    .B1_N(_08453_),
    .X(_08597_));
 sky130_fd_sc_hd__or2_1 _24499_ (.A(_07273_),
    .B(_05831_),
    .X(_08598_));
 sky130_fd_sc_hd__clkbuf_2 _24500_ (.A(_07397_),
    .X(_08599_));
 sky130_fd_sc_hd__buf_1 _24501_ (.A(_08599_),
    .X(_08600_));
 sky130_fd_sc_hd__buf_1 _24502_ (.A(_07267_),
    .X(_08601_));
 sky130_fd_sc_hd__o22a_1 _24503_ (.A1(_08600_),
    .A2(_08439_),
    .B1(_08601_),
    .B2(_07126_),
    .X(_08602_));
 sky130_fd_sc_hd__buf_1 _24504_ (.A(_13087_),
    .X(_08603_));
 sky130_fd_sc_hd__and4_1 _24505_ (.A(_08603_),
    .B(_13595_),
    .C(_08441_),
    .D(_13592_),
    .X(_08604_));
 sky130_fd_sc_hd__or2_1 _24506_ (.A(_08602_),
    .B(_08604_),
    .X(_08605_));
 sky130_fd_sc_hd__a2bb2o_1 _24507_ (.A1_N(_08598_),
    .A2_N(_08605_),
    .B1(_08598_),
    .B2(_08605_),
    .X(_08606_));
 sky130_fd_sc_hd__a2bb2o_1 _24508_ (.A1_N(_08597_),
    .A2_N(_08606_),
    .B1(_08597_),
    .B2(_08606_),
    .X(_08607_));
 sky130_fd_sc_hd__a2bb2o_1 _24509_ (.A1_N(_08596_),
    .A2_N(_08607_),
    .B1(_08596_),
    .B2(_08607_),
    .X(_08608_));
 sky130_fd_sc_hd__clkbuf_2 _24510_ (.A(_07530_),
    .X(_08609_));
 sky130_fd_sc_hd__or2_1 _24511_ (.A(_08609_),
    .B(_07278_),
    .X(_08610_));
 sky130_fd_sc_hd__clkbuf_2 _24512_ (.A(_08285_),
    .X(_08611_));
 sky130_fd_sc_hd__o22a_1 _24513_ (.A1(_08611_),
    .A2(_08283_),
    .B1(_07684_),
    .B2(_07079_),
    .X(_08612_));
 sky130_fd_sc_hd__buf_1 _24514_ (.A(_13072_),
    .X(_08613_));
 sky130_fd_sc_hd__buf_1 _24515_ (.A(_13078_),
    .X(_08614_));
 sky130_fd_sc_hd__and4_1 _24516_ (.A(_08613_),
    .B(_13609_),
    .C(_08614_),
    .D(_13604_),
    .X(_08615_));
 sky130_fd_sc_hd__or2_1 _24517_ (.A(_08612_),
    .B(_08615_),
    .X(_08616_));
 sky130_fd_sc_hd__a2bb2o_1 _24518_ (.A1_N(_08610_),
    .A2_N(_08616_),
    .B1(_08610_),
    .B2(_08616_),
    .X(_08617_));
 sky130_fd_sc_hd__or2_1 _24519_ (.A(_08292_),
    .B(_08136_),
    .X(_08618_));
 sky130_fd_sc_hd__and4_1 _24520_ (.A(_08295_),
    .B(_06015_),
    .C(_13064_),
    .D(_13616_),
    .X(_08619_));
 sky130_fd_sc_hd__clkbuf_2 _24521_ (.A(_11716_),
    .X(_08620_));
 sky130_fd_sc_hd__o22a_1 _24522_ (.A1(_08620_),
    .A2(_13620_),
    .B1(_08131_),
    .B2(_05339_),
    .X(_08621_));
 sky130_fd_sc_hd__or2_1 _24523_ (.A(_08619_),
    .B(_08621_),
    .X(_08622_));
 sky130_fd_sc_hd__a2bb2o_1 _24524_ (.A1_N(_08618_),
    .A2_N(_08622_),
    .B1(_08618_),
    .B2(_08622_),
    .X(_08623_));
 sky130_fd_sc_hd__o21ba_1 _24525_ (.A1(_08456_),
    .A2(_08460_),
    .B1_N(_08458_),
    .X(_08624_));
 sky130_fd_sc_hd__a2bb2o_1 _24526_ (.A1_N(_08623_),
    .A2_N(_08624_),
    .B1(_08623_),
    .B2(_08624_),
    .X(_08625_));
 sky130_fd_sc_hd__a2bb2o_1 _24527_ (.A1_N(_08617_),
    .A2_N(_08625_),
    .B1(_08617_),
    .B2(_08625_),
    .X(_08626_));
 sky130_fd_sc_hd__o22a_1 _24528_ (.A1(_08461_),
    .A2(_08462_),
    .B1(_08455_),
    .B2(_08463_),
    .X(_08627_));
 sky130_fd_sc_hd__a2bb2o_1 _24529_ (.A1_N(_08626_),
    .A2_N(_08627_),
    .B1(_08626_),
    .B2(_08627_),
    .X(_08628_));
 sky130_fd_sc_hd__a2bb2o_1 _24530_ (.A1_N(_08608_),
    .A2_N(_08628_),
    .B1(_08608_),
    .B2(_08628_),
    .X(_08629_));
 sky130_fd_sc_hd__o22a_1 _24531_ (.A1(_08464_),
    .A2(_08465_),
    .B1(_08446_),
    .B2(_08466_),
    .X(_08630_));
 sky130_fd_sc_hd__a2bb2o_1 _24532_ (.A1_N(_08629_),
    .A2_N(_08630_),
    .B1(_08629_),
    .B2(_08630_),
    .X(_08631_));
 sky130_fd_sc_hd__a2bb2o_1 _24533_ (.A1_N(_08595_),
    .A2_N(_08631_),
    .B1(_08595_),
    .B2(_08631_),
    .X(_08632_));
 sky130_fd_sc_hd__o22a_1 _24534_ (.A1(_08467_),
    .A2(_08468_),
    .B1(_08435_),
    .B2(_08469_),
    .X(_08633_));
 sky130_fd_sc_hd__a2bb2o_1 _24535_ (.A1_N(_08632_),
    .A2_N(_08633_),
    .B1(_08632_),
    .B2(_08633_),
    .X(_08634_));
 sky130_fd_sc_hd__a2bb2o_1 _24536_ (.A1_N(_08570_),
    .A2_N(_08634_),
    .B1(_08570_),
    .B2(_08634_),
    .X(_08635_));
 sky130_fd_sc_hd__o22a_1 _24537_ (.A1(_08470_),
    .A2(_08471_),
    .B1(_08412_),
    .B2(_08472_),
    .X(_08636_));
 sky130_fd_sc_hd__a2bb2o_1 _24538_ (.A1_N(_08635_),
    .A2_N(_08636_),
    .B1(_08635_),
    .B2(_08636_),
    .X(_08637_));
 sky130_fd_sc_hd__a2bb2o_1 _24539_ (.A1_N(_08532_),
    .A2_N(_08637_),
    .B1(_08532_),
    .B2(_08637_),
    .X(_08638_));
 sky130_fd_sc_hd__o22a_1 _24540_ (.A1(_08473_),
    .A2(_08474_),
    .B1(_08378_),
    .B2(_08475_),
    .X(_08639_));
 sky130_fd_sc_hd__a2bb2o_1 _24541_ (.A1_N(_08638_),
    .A2_N(_08639_),
    .B1(_08638_),
    .B2(_08639_),
    .X(_08640_));
 sky130_fd_sc_hd__a2bb2o_1 _24542_ (.A1_N(_08489_),
    .A2_N(_08640_),
    .B1(_08489_),
    .B2(_08640_),
    .X(_08641_));
 sky130_fd_sc_hd__o22a_1 _24543_ (.A1(_08476_),
    .A2(_08477_),
    .B1(_08335_),
    .B2(_08478_),
    .X(_08642_));
 sky130_fd_sc_hd__a2bb2o_1 _24544_ (.A1_N(_08641_),
    .A2_N(_08642_),
    .B1(_08641_),
    .B2(_08642_),
    .X(_08643_));
 sky130_fd_sc_hd__a2bb2o_1 _24545_ (.A1_N(_08334_),
    .A2_N(_08643_),
    .B1(_08334_),
    .B2(_08643_),
    .X(_08644_));
 sky130_fd_sc_hd__o22a_1 _24546_ (.A1(_08479_),
    .A2(_08480_),
    .B1(_08331_),
    .B2(_08481_),
    .X(_08645_));
 sky130_fd_sc_hd__or2_1 _24547_ (.A(_08644_),
    .B(_08645_),
    .X(_08646_));
 sky130_vsdinv _24548_ (.A(_08646_),
    .Y(_08647_));
 sky130_fd_sc_hd__a21o_2 _24549_ (.A1(_08644_),
    .A2(_08645_),
    .B1(_08647_),
    .X(_08648_));
 sky130_fd_sc_hd__a22o_1 _24550_ (.A1(_08482_),
    .A2(_08483_),
    .B1(_08320_),
    .B2(_08484_),
    .X(_08649_));
 sky130_fd_sc_hd__o31a_2 _24551_ (.A1(_08322_),
    .A2(_08485_),
    .A3(_08329_),
    .B1(_08649_),
    .X(_08650_));
 sky130_fd_sc_hd__a2bb2oi_4 _24552_ (.A1_N(_08648_),
    .A2_N(_08650_),
    .B1(_08648_),
    .B2(_08650_),
    .Y(_02653_));
 sky130_fd_sc_hd__o22a_1 _24553_ (.A1(_08641_),
    .A2(_08642_),
    .B1(_08334_),
    .B2(_08643_),
    .X(_08651_));
 sky130_vsdinv _24554_ (.A(_08651_),
    .Y(_08652_));
 sky130_fd_sc_hd__o22a_1 _24555_ (.A1(_08491_),
    .A2(_08530_),
    .B1(_08490_),
    .B2(_08531_),
    .X(_08653_));
 sky130_fd_sc_hd__o22a_4 _24556_ (.A1(_08510_),
    .A2(_08511_),
    .B1(_08492_),
    .B2(_08512_),
    .X(_08654_));
 sky130_fd_sc_hd__or2_1 _24557_ (.A(_08653_),
    .B(_08654_),
    .X(_08655_));
 sky130_fd_sc_hd__a21bo_1 _24558_ (.A1(_08653_),
    .A2(_08654_),
    .B1_N(_08655_),
    .X(_08656_));
 sky130_fd_sc_hd__o22a_2 _24559_ (.A1(_08527_),
    .A2(_08528_),
    .B1(_08513_),
    .B2(_08529_),
    .X(_08657_));
 sky130_fd_sc_hd__o22a_1 _24560_ (.A1(_08534_),
    .A2(_08568_),
    .B1(_08533_),
    .B2(_08569_),
    .X(_08658_));
 sky130_fd_sc_hd__a21oi_1 _24561_ (.A1(_08496_),
    .A2(_08501_),
    .B1(_08494_),
    .Y(_08659_));
 sky130_fd_sc_hd__buf_1 _24562_ (.A(_08340_),
    .X(_08660_));
 sky130_fd_sc_hd__buf_2 _24563_ (.A(_08660_),
    .X(_08661_));
 sky130_fd_sc_hd__nor2_4 _24564_ (.A(_08661_),
    .B(_05827_),
    .Y(_08662_));
 sky130_fd_sc_hd__a2bb2o_1 _24565_ (.A1_N(_08495_),
    .A2_N(_08662_),
    .B1(_08495_),
    .B2(_08662_),
    .X(_08663_));
 sky130_fd_sc_hd__buf_1 _24566_ (.A(_08663_),
    .X(_08664_));
 sky130_fd_sc_hd__buf_1 _24567_ (.A(_08664_),
    .X(_08665_));
 sky130_fd_sc_hd__o22a_1 _24568_ (.A1(_07181_),
    .A2(_07890_),
    .B1(_07183_),
    .B2(_08034_),
    .X(_08666_));
 sky130_fd_sc_hd__buf_1 _24569_ (.A(\pcpi_mul.rs1[30] ),
    .X(_08667_));
 sky130_fd_sc_hd__buf_1 _24570_ (.A(\pcpi_mul.rs1[31] ),
    .X(_08668_));
 sky130_fd_sc_hd__and4_1 _24571_ (.A(_06233_),
    .B(_08667_),
    .C(_06235_),
    .D(_08668_),
    .X(_08669_));
 sky130_fd_sc_hd__or2_1 _24572_ (.A(_08666_),
    .B(_08669_),
    .X(_08670_));
 sky130_vsdinv _24573_ (.A(_08670_),
    .Y(_08671_));
 sky130_fd_sc_hd__a22o_1 _24574_ (.A1(_08186_),
    .A2(_08671_),
    .B1(_08184_),
    .B2(_08670_),
    .X(_08672_));
 sky130_fd_sc_hd__a21oi_2 _24575_ (.A1(_08353_),
    .A2(_08506_),
    .B1(_08504_),
    .Y(_08673_));
 sky130_fd_sc_hd__a2bb2o_1 _24576_ (.A1_N(_08672_),
    .A2_N(_08673_),
    .B1(_08672_),
    .B2(_08673_),
    .X(_08674_));
 sky130_fd_sc_hd__a2bb2o_1 _24577_ (.A1_N(_08665_),
    .A2_N(_08674_),
    .B1(_08665_),
    .B2(_08674_),
    .X(_08675_));
 sky130_fd_sc_hd__o22a_1 _24578_ (.A1(_08507_),
    .A2(_08508_),
    .B1(_08502_),
    .B2(_08509_),
    .X(_08676_));
 sky130_fd_sc_hd__a2bb2o_1 _24579_ (.A1_N(_08675_),
    .A2_N(_08676_),
    .B1(_08675_),
    .B2(_08676_),
    .X(_08677_));
 sky130_fd_sc_hd__a2bb2o_1 _24580_ (.A1_N(_08659_),
    .A2_N(_08677_),
    .B1(_08659_),
    .B2(_08677_),
    .X(_08678_));
 sky130_fd_sc_hd__o22a_1 _24581_ (.A1(_08517_),
    .A2(_08523_),
    .B1(_08516_),
    .B2(_08524_),
    .X(_08679_));
 sky130_fd_sc_hd__o22a_1 _24582_ (.A1(_08551_),
    .A2(_08552_),
    .B1(_08542_),
    .B2(_08553_),
    .X(_08680_));
 sky130_fd_sc_hd__a21oi_2 _24583_ (.A1(_08521_),
    .A2(_08522_),
    .B1(_08520_),
    .Y(_08681_));
 sky130_fd_sc_hd__o21ba_1 _24584_ (.A1(_08536_),
    .A2(_08541_),
    .B1_N(_08540_),
    .X(_08682_));
 sky130_fd_sc_hd__clkbuf_2 _24585_ (.A(_06671_),
    .X(_08683_));
 sky130_fd_sc_hd__buf_1 _24586_ (.A(_07462_),
    .X(_08684_));
 sky130_fd_sc_hd__o22a_1 _24587_ (.A1(_08683_),
    .A2(_08684_),
    .B1(_08518_),
    .B2(_07870_),
    .X(_08685_));
 sky130_fd_sc_hd__buf_1 _24588_ (.A(_13523_),
    .X(_08686_));
 sky130_fd_sc_hd__and4_1 _24589_ (.A(_13149_),
    .B(_08686_),
    .C(_13155_),
    .D(_07877_),
    .X(_08687_));
 sky130_fd_sc_hd__nor2_1 _24590_ (.A(_08685_),
    .B(_08687_),
    .Y(_08688_));
 sky130_fd_sc_hd__nor2_1 _24591_ (.A(_05425_),
    .B(_07749_),
    .Y(_08689_));
 sky130_fd_sc_hd__a2bb2o_1 _24592_ (.A1_N(_08688_),
    .A2_N(_08689_),
    .B1(_08688_),
    .B2(_08689_),
    .X(_08690_));
 sky130_fd_sc_hd__a2bb2o_1 _24593_ (.A1_N(_08682_),
    .A2_N(_08690_),
    .B1(_08682_),
    .B2(_08690_),
    .X(_08691_));
 sky130_fd_sc_hd__a2bb2o_1 _24594_ (.A1_N(_08681_),
    .A2_N(_08691_),
    .B1(_08681_),
    .B2(_08691_),
    .X(_08692_));
 sky130_fd_sc_hd__a2bb2o_1 _24595_ (.A1_N(_08680_),
    .A2_N(_08692_),
    .B1(_08680_),
    .B2(_08692_),
    .X(_08693_));
 sky130_fd_sc_hd__a2bb2o_1 _24596_ (.A1_N(_08679_),
    .A2_N(_08693_),
    .B1(_08679_),
    .B2(_08693_),
    .X(_08694_));
 sky130_fd_sc_hd__o22a_1 _24597_ (.A1(_08515_),
    .A2(_08525_),
    .B1(_08514_),
    .B2(_08526_),
    .X(_08695_));
 sky130_fd_sc_hd__a2bb2o_1 _24598_ (.A1_N(_08694_),
    .A2_N(_08695_),
    .B1(_08694_),
    .B2(_08695_),
    .X(_08696_));
 sky130_fd_sc_hd__a2bb2o_2 _24599_ (.A1_N(_08678_),
    .A2_N(_08696_),
    .B1(_08678_),
    .B2(_08696_),
    .X(_08697_));
 sky130_fd_sc_hd__a2bb2o_1 _24600_ (.A1_N(_08658_),
    .A2_N(_08697_),
    .B1(_08658_),
    .B2(_08697_),
    .X(_08698_));
 sky130_fd_sc_hd__a2bb2o_1 _24601_ (.A1_N(_08657_),
    .A2_N(_08698_),
    .B1(_08657_),
    .B2(_08698_),
    .X(_08699_));
 sky130_fd_sc_hd__o22a_1 _24602_ (.A1(_08565_),
    .A2(_08566_),
    .B1(_08554_),
    .B2(_08567_),
    .X(_08700_));
 sky130_fd_sc_hd__o22a_1 _24603_ (.A1(_08572_),
    .A2(_08593_),
    .B1(_08571_),
    .B2(_08594_),
    .X(_08701_));
 sky130_fd_sc_hd__or2_1 _24604_ (.A(_05537_),
    .B(_07884_),
    .X(_08702_));
 sky130_fd_sc_hd__o22a_1 _24605_ (.A1(_08217_),
    .A2(_07032_),
    .B1(_08538_),
    .B2(_08198_),
    .X(_08703_));
 sky130_fd_sc_hd__and4_1 _24606_ (.A(_07363_),
    .B(_13538_),
    .C(_07364_),
    .D(_07741_),
    .X(_08704_));
 sky130_fd_sc_hd__or2_1 _24607_ (.A(_08703_),
    .B(_08704_),
    .X(_08705_));
 sky130_fd_sc_hd__a2bb2o_1 _24608_ (.A1_N(_08702_),
    .A2_N(_08705_),
    .B1(_08702_),
    .B2(_08705_),
    .X(_08706_));
 sky130_fd_sc_hd__or2_1 _24609_ (.A(_08386_),
    .B(_07019_),
    .X(_08707_));
 sky130_fd_sc_hd__clkbuf_2 _24610_ (.A(_06533_),
    .X(_08708_));
 sky130_fd_sc_hd__o22a_1 _24611_ (.A1(_08544_),
    .A2(_06877_),
    .B1(_08708_),
    .B2(_07905_),
    .X(_08709_));
 sky130_fd_sc_hd__and4_1 _24612_ (.A(_08390_),
    .B(_13549_),
    .C(_08391_),
    .D(_07907_),
    .X(_08710_));
 sky130_fd_sc_hd__or2_1 _24613_ (.A(_08709_),
    .B(_08710_),
    .X(_08711_));
 sky130_fd_sc_hd__a2bb2o_1 _24614_ (.A1_N(_08707_),
    .A2_N(_08711_),
    .B1(_08707_),
    .B2(_08711_),
    .X(_08712_));
 sky130_fd_sc_hd__o21ba_1 _24615_ (.A1(_08543_),
    .A2(_08550_),
    .B1_N(_08549_),
    .X(_08713_));
 sky130_fd_sc_hd__a2bb2o_1 _24616_ (.A1_N(_08712_),
    .A2_N(_08713_),
    .B1(_08712_),
    .B2(_08713_),
    .X(_08714_));
 sky130_fd_sc_hd__a2bb2o_2 _24617_ (.A1_N(_08706_),
    .A2_N(_08714_),
    .B1(_08706_),
    .B2(_08714_),
    .X(_08715_));
 sky130_fd_sc_hd__o21ba_1 _24618_ (.A1(_08558_),
    .A2(_08562_),
    .B1_N(_08561_),
    .X(_08716_));
 sky130_fd_sc_hd__o21ba_1 _24619_ (.A1(_08573_),
    .A2(_08580_),
    .B1_N(_08579_),
    .X(_08717_));
 sky130_fd_sc_hd__or2_1 _24620_ (.A(_08241_),
    .B(_06641_),
    .X(_08718_));
 sky130_fd_sc_hd__buf_1 _24621_ (.A(_06450_),
    .X(_08719_));
 sky130_fd_sc_hd__o22a_1 _24622_ (.A1(_08233_),
    .A2(_08559_),
    .B1(_08401_),
    .B2(_08719_),
    .X(_08720_));
 sky130_fd_sc_hd__buf_1 _24623_ (.A(_07484_),
    .X(_08721_));
 sky130_fd_sc_hd__and4_1 _24624_ (.A(_08236_),
    .B(_13560_),
    .C(_08238_),
    .D(_08721_),
    .X(_08722_));
 sky130_fd_sc_hd__or2_1 _24625_ (.A(_08720_),
    .B(_08722_),
    .X(_08723_));
 sky130_fd_sc_hd__a2bb2o_1 _24626_ (.A1_N(_08718_),
    .A2_N(_08723_),
    .B1(_08718_),
    .B2(_08723_),
    .X(_08724_));
 sky130_fd_sc_hd__a2bb2o_1 _24627_ (.A1_N(_08717_),
    .A2_N(_08724_),
    .B1(_08717_),
    .B2(_08724_),
    .X(_08725_));
 sky130_fd_sc_hd__a2bb2o_1 _24628_ (.A1_N(_08716_),
    .A2_N(_08725_),
    .B1(_08716_),
    .B2(_08725_),
    .X(_08726_));
 sky130_fd_sc_hd__o22a_1 _24629_ (.A1(_08556_),
    .A2(_08563_),
    .B1(_08555_),
    .B2(_08564_),
    .X(_08727_));
 sky130_fd_sc_hd__a2bb2o_1 _24630_ (.A1_N(_08726_),
    .A2_N(_08727_),
    .B1(_08726_),
    .B2(_08727_),
    .X(_08728_));
 sky130_fd_sc_hd__a2bb2o_1 _24631_ (.A1_N(_08715_),
    .A2_N(_08728_),
    .B1(_08715_),
    .B2(_08728_),
    .X(_08729_));
 sky130_fd_sc_hd__a2bb2o_1 _24632_ (.A1_N(_08701_),
    .A2_N(_08729_),
    .B1(_08701_),
    .B2(_08729_),
    .X(_08730_));
 sky130_fd_sc_hd__a2bb2o_1 _24633_ (.A1_N(_08700_),
    .A2_N(_08730_),
    .B1(_08700_),
    .B2(_08730_),
    .X(_08731_));
 sky130_fd_sc_hd__o22a_1 _24634_ (.A1(_08590_),
    .A2(_08591_),
    .B1(_08581_),
    .B2(_08592_),
    .X(_08732_));
 sky130_fd_sc_hd__o22a_1 _24635_ (.A1(_08597_),
    .A2(_08606_),
    .B1(_08596_),
    .B2(_08607_),
    .X(_08733_));
 sky130_fd_sc_hd__clkbuf_4 _24636_ (.A(_06284_),
    .X(_08734_));
 sky130_fd_sc_hd__or2_1 _24637_ (.A(_08734_),
    .B(_06330_),
    .X(_08735_));
 sky130_fd_sc_hd__buf_2 _24638_ (.A(_06389_),
    .X(_08736_));
 sky130_fd_sc_hd__o22a_1 _24639_ (.A1(_08574_),
    .A2(_08234_),
    .B1(_08736_),
    .B2(_06218_),
    .X(_08737_));
 sky130_fd_sc_hd__buf_1 _24640_ (.A(_13566_),
    .X(_08738_));
 sky130_fd_sc_hd__and4_1 _24641_ (.A(_08577_),
    .B(_08237_),
    .C(_13112_),
    .D(_08738_),
    .X(_08739_));
 sky130_fd_sc_hd__or2_1 _24642_ (.A(_08737_),
    .B(_08739_),
    .X(_08740_));
 sky130_fd_sc_hd__a2bb2o_2 _24643_ (.A1_N(_08735_),
    .A2_N(_08740_),
    .B1(_08735_),
    .B2(_08740_),
    .X(_08741_));
 sky130_fd_sc_hd__or2_1 _24644_ (.A(_08582_),
    .B(_06032_),
    .X(_08742_));
 sky130_fd_sc_hd__buf_1 _24645_ (.A(_08261_),
    .X(_08743_));
 sky130_fd_sc_hd__o22a_1 _24646_ (.A1(_08743_),
    .A2(_05820_),
    .B1(_06806_),
    .B2(_05931_),
    .X(_08744_));
 sky130_fd_sc_hd__clkbuf_2 _24647_ (.A(_13096_),
    .X(_08745_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _24648_ (.A(_13101_),
    .X(_08746_));
 sky130_fd_sc_hd__buf_1 _24649_ (.A(_13578_),
    .X(_08747_));
 sky130_fd_sc_hd__and4_1 _24650_ (.A(_08745_),
    .B(_08587_),
    .C(_08746_),
    .D(_08747_),
    .X(_08748_));
 sky130_fd_sc_hd__or2_1 _24651_ (.A(_08744_),
    .B(_08748_),
    .X(_08749_));
 sky130_fd_sc_hd__a2bb2o_1 _24652_ (.A1_N(_08742_),
    .A2_N(_08749_),
    .B1(_08742_),
    .B2(_08749_),
    .X(_08750_));
 sky130_fd_sc_hd__o21ba_1 _24653_ (.A1(_08583_),
    .A2(_08589_),
    .B1_N(_08588_),
    .X(_08751_));
 sky130_fd_sc_hd__a2bb2o_1 _24654_ (.A1_N(_08750_),
    .A2_N(_08751_),
    .B1(_08750_),
    .B2(_08751_),
    .X(_08752_));
 sky130_fd_sc_hd__a2bb2o_1 _24655_ (.A1_N(_08741_),
    .A2_N(_08752_),
    .B1(_08741_),
    .B2(_08752_),
    .X(_08753_));
 sky130_fd_sc_hd__a2bb2o_1 _24656_ (.A1_N(_08733_),
    .A2_N(_08753_),
    .B1(_08733_),
    .B2(_08753_),
    .X(_08754_));
 sky130_fd_sc_hd__a2bb2o_1 _24657_ (.A1_N(_08732_),
    .A2_N(_08754_),
    .B1(_08732_),
    .B2(_08754_),
    .X(_08755_));
 sky130_fd_sc_hd__o21ba_1 _24658_ (.A1(_08598_),
    .A2(_08605_),
    .B1_N(_08604_),
    .X(_08756_));
 sky130_fd_sc_hd__o21ba_1 _24659_ (.A1(_08610_),
    .A2(_08616_),
    .B1_N(_08615_),
    .X(_08757_));
 sky130_fd_sc_hd__buf_2 _24660_ (.A(_07073_),
    .X(_08758_));
 sky130_fd_sc_hd__or2_1 _24661_ (.A(_08758_),
    .B(_05818_),
    .X(_08759_));
 sky130_fd_sc_hd__o22a_1 _24662_ (.A1(_08600_),
    .A2(_07126_),
    .B1(_08601_),
    .B2(_05723_),
    .X(_08760_));
 sky130_fd_sc_hd__buf_1 _24663_ (.A(_13087_),
    .X(_08761_));
 sky130_fd_sc_hd__and4_1 _24664_ (.A(_08761_),
    .B(_13592_),
    .C(_13092_),
    .D(_13588_),
    .X(_08762_));
 sky130_fd_sc_hd__or2_1 _24665_ (.A(_08760_),
    .B(_08762_),
    .X(_08763_));
 sky130_fd_sc_hd__a2bb2o_1 _24666_ (.A1_N(_08759_),
    .A2_N(_08763_),
    .B1(_08759_),
    .B2(_08763_),
    .X(_08764_));
 sky130_fd_sc_hd__a2bb2o_1 _24667_ (.A1_N(_08757_),
    .A2_N(_08764_),
    .B1(_08757_),
    .B2(_08764_),
    .X(_08765_));
 sky130_fd_sc_hd__a2bb2o_1 _24668_ (.A1_N(_08756_),
    .A2_N(_08765_),
    .B1(_08756_),
    .B2(_08765_),
    .X(_08766_));
 sky130_fd_sc_hd__or2_1 _24669_ (.A(_07531_),
    .B(_07403_),
    .X(_08767_));
 sky130_fd_sc_hd__o22a_1 _24670_ (.A1(_08611_),
    .A2(_07983_),
    .B1(_07684_),
    .B2(_05862_),
    .X(_08768_));
 sky130_fd_sc_hd__and4_1 _24671_ (.A(_08613_),
    .B(_13604_),
    .C(_08614_),
    .D(_13599_),
    .X(_08769_));
 sky130_fd_sc_hd__or2_1 _24672_ (.A(_08768_),
    .B(_08769_),
    .X(_08770_));
 sky130_fd_sc_hd__a2bb2o_1 _24673_ (.A1_N(_08767_),
    .A2_N(_08770_),
    .B1(_08767_),
    .B2(_08770_),
    .X(_08771_));
 sky130_fd_sc_hd__buf_1 _24674_ (.A(_07971_),
    .X(_08772_));
 sky130_fd_sc_hd__or2_1 _24675_ (.A(_08772_),
    .B(_08283_),
    .X(_08773_));
 sky130_fd_sc_hd__buf_1 _24676_ (.A(_08294_),
    .X(_08774_));
 sky130_fd_sc_hd__buf_1 _24677_ (.A(_08457_),
    .X(_08775_));
 sky130_fd_sc_hd__and4_1 _24678_ (.A(_08774_),
    .B(_05339_),
    .C(_08775_),
    .D(_07085_),
    .X(_08776_));
 sky130_fd_sc_hd__buf_1 _24679_ (.A(_11717_),
    .X(_08777_));
 sky130_fd_sc_hd__buf_1 _24680_ (.A(_08130_),
    .X(_08778_));
 sky130_fd_sc_hd__o22a_1 _24681_ (.A1(_08777_),
    .A2(_13616_),
    .B1(_08778_),
    .B2(_07082_),
    .X(_08779_));
 sky130_fd_sc_hd__or2_1 _24682_ (.A(_08776_),
    .B(_08779_),
    .X(_08780_));
 sky130_fd_sc_hd__a2bb2o_1 _24683_ (.A1_N(_08773_),
    .A2_N(_08780_),
    .B1(_08773_),
    .B2(_08780_),
    .X(_08781_));
 sky130_fd_sc_hd__o21ba_1 _24684_ (.A1(_08618_),
    .A2(_08622_),
    .B1_N(_08619_),
    .X(_08782_));
 sky130_fd_sc_hd__a2bb2o_1 _24685_ (.A1_N(_08781_),
    .A2_N(_08782_),
    .B1(_08781_),
    .B2(_08782_),
    .X(_08783_));
 sky130_fd_sc_hd__a2bb2o_1 _24686_ (.A1_N(_08771_),
    .A2_N(_08783_),
    .B1(_08771_),
    .B2(_08783_),
    .X(_08784_));
 sky130_fd_sc_hd__o22a_1 _24687_ (.A1(_08623_),
    .A2(_08624_),
    .B1(_08617_),
    .B2(_08625_),
    .X(_08785_));
 sky130_fd_sc_hd__a2bb2o_1 _24688_ (.A1_N(_08784_),
    .A2_N(_08785_),
    .B1(_08784_),
    .B2(_08785_),
    .X(_08786_));
 sky130_fd_sc_hd__a2bb2o_1 _24689_ (.A1_N(_08766_),
    .A2_N(_08786_),
    .B1(_08766_),
    .B2(_08786_),
    .X(_08787_));
 sky130_fd_sc_hd__o22a_1 _24690_ (.A1(_08626_),
    .A2(_08627_),
    .B1(_08608_),
    .B2(_08628_),
    .X(_08788_));
 sky130_fd_sc_hd__a2bb2o_1 _24691_ (.A1_N(_08787_),
    .A2_N(_08788_),
    .B1(_08787_),
    .B2(_08788_),
    .X(_08789_));
 sky130_fd_sc_hd__a2bb2o_1 _24692_ (.A1_N(_08755_),
    .A2_N(_08789_),
    .B1(_08755_),
    .B2(_08789_),
    .X(_08790_));
 sky130_fd_sc_hd__o22a_1 _24693_ (.A1(_08629_),
    .A2(_08630_),
    .B1(_08595_),
    .B2(_08631_),
    .X(_08791_));
 sky130_fd_sc_hd__a2bb2o_1 _24694_ (.A1_N(_08790_),
    .A2_N(_08791_),
    .B1(_08790_),
    .B2(_08791_),
    .X(_08792_));
 sky130_fd_sc_hd__a2bb2o_1 _24695_ (.A1_N(_08731_),
    .A2_N(_08792_),
    .B1(_08731_),
    .B2(_08792_),
    .X(_08793_));
 sky130_fd_sc_hd__o22a_1 _24696_ (.A1(_08632_),
    .A2(_08633_),
    .B1(_08570_),
    .B2(_08634_),
    .X(_08794_));
 sky130_fd_sc_hd__a2bb2o_1 _24697_ (.A1_N(_08793_),
    .A2_N(_08794_),
    .B1(_08793_),
    .B2(_08794_),
    .X(_08795_));
 sky130_fd_sc_hd__a2bb2o_1 _24698_ (.A1_N(_08699_),
    .A2_N(_08795_),
    .B1(_08699_),
    .B2(_08795_),
    .X(_08796_));
 sky130_fd_sc_hd__o22a_1 _24699_ (.A1(_08635_),
    .A2(_08636_),
    .B1(_08532_),
    .B2(_08637_),
    .X(_08797_));
 sky130_fd_sc_hd__a2bb2o_1 _24700_ (.A1_N(_08796_),
    .A2_N(_08797_),
    .B1(_08796_),
    .B2(_08797_),
    .X(_08798_));
 sky130_fd_sc_hd__a2bb2o_1 _24701_ (.A1_N(_08656_),
    .A2_N(_08798_),
    .B1(_08656_),
    .B2(_08798_),
    .X(_08799_));
 sky130_fd_sc_hd__o22a_1 _24702_ (.A1(_08638_),
    .A2(_08639_),
    .B1(_08489_),
    .B2(_08640_),
    .X(_08800_));
 sky130_fd_sc_hd__a2bb2o_1 _24703_ (.A1_N(_08799_),
    .A2_N(_08800_),
    .B1(_08799_),
    .B2(_08800_),
    .X(_08801_));
 sky130_fd_sc_hd__a2bb2o_1 _24704_ (.A1_N(_08488_),
    .A2_N(_08801_),
    .B1(_08488_),
    .B2(_08801_),
    .X(_08802_));
 sky130_vsdinv _24705_ (.A(_08802_),
    .Y(_08803_));
 sky130_fd_sc_hd__a22o_1 _24706_ (.A1(_08652_),
    .A2(_08803_),
    .B1(_08651_),
    .B2(_08802_),
    .X(_08804_));
 sky130_fd_sc_hd__o21ai_2 _24707_ (.A1(_08648_),
    .A2(_08650_),
    .B1(_08646_),
    .Y(_08805_));
 sky130_fd_sc_hd__a2bb2o_4 _24708_ (.A1_N(_08804_),
    .A2_N(_08805_),
    .B1(_08804_),
    .B2(_08805_),
    .X(_02654_));
 sky130_fd_sc_hd__o22a_1 _24709_ (.A1(_08658_),
    .A2(_08697_),
    .B1(_08657_),
    .B2(_08698_),
    .X(_08806_));
 sky130_fd_sc_hd__o22a_2 _24710_ (.A1(_08675_),
    .A2(_08676_),
    .B1(_08659_),
    .B2(_08677_),
    .X(_08807_));
 sky130_fd_sc_hd__or2_1 _24711_ (.A(_08806_),
    .B(_08807_),
    .X(_08808_));
 sky130_fd_sc_hd__a21bo_1 _24712_ (.A1(_08806_),
    .A2(_08807_),
    .B1_N(_08808_),
    .X(_08809_));
 sky130_fd_sc_hd__o22a_2 _24713_ (.A1(_08694_),
    .A2(_08695_),
    .B1(_08678_),
    .B2(_08696_),
    .X(_08810_));
 sky130_fd_sc_hd__o22a_1 _24714_ (.A1(_08701_),
    .A2(_08729_),
    .B1(_08700_),
    .B2(_08730_),
    .X(_08811_));
 sky130_fd_sc_hd__a21oi_2 _24715_ (.A1(_08496_),
    .A2(_08662_),
    .B1(_08494_),
    .Y(_08812_));
 sky130_fd_sc_hd__buf_1 _24716_ (.A(_08812_),
    .X(_08813_));
 sky130_fd_sc_hd__clkbuf_2 _24717_ (.A(\pcpi_mul.rs1[32] ),
    .X(_08814_));
 sky130_fd_sc_hd__buf_1 _24718_ (.A(_08814_),
    .X(_08815_));
 sky130_fd_sc_hd__buf_2 _24719_ (.A(_08815_),
    .X(_08816_));
 sky130_fd_sc_hd__a31o_1 _24720_ (.A1(_08816_),
    .A2(\pcpi_mul.rs2[0] ),
    .A3(_08671_),
    .B1(_08669_),
    .X(_08817_));
 sky130_vsdinv _24721_ (.A(_08817_),
    .Y(_08818_));
 sky130_fd_sc_hd__o22a_2 _24722_ (.A1(_06894_),
    .A2(_08035_),
    .B1(_11703_),
    .B2(_06895_),
    .X(_08819_));
 sky130_fd_sc_hd__clkbuf_2 _24723_ (.A(_13505_),
    .X(_08820_));
 sky130_fd_sc_hd__and4_1 _24724_ (.A(_07186_),
    .B(_08820_),
    .C(_08815_),
    .D(_07189_),
    .X(_08821_));
 sky130_fd_sc_hd__nor2_1 _24725_ (.A(_08819_),
    .B(_08821_),
    .Y(_08822_));
 sky130_fd_sc_hd__o2bb2a_1 _24726_ (.A1_N(_08347_),
    .A2_N(_08822_),
    .B1(_08347_),
    .B2(_08822_),
    .X(_08823_));
 sky130_vsdinv _24727_ (.A(_08823_),
    .Y(_08824_));
 sky130_fd_sc_hd__a22o_1 _24728_ (.A1(_08818_),
    .A2(_08824_),
    .B1(_08817_),
    .B2(_08823_),
    .X(_08825_));
 sky130_fd_sc_hd__a2bb2o_1 _24729_ (.A1_N(_08665_),
    .A2_N(_08825_),
    .B1(_08664_),
    .B2(_08825_),
    .X(_08826_));
 sky130_fd_sc_hd__o22a_1 _24730_ (.A1(_08672_),
    .A2(_08673_),
    .B1(_08665_),
    .B2(_08674_),
    .X(_08827_));
 sky130_fd_sc_hd__a2bb2o_1 _24731_ (.A1_N(_08826_),
    .A2_N(_08827_),
    .B1(_08826_),
    .B2(_08827_),
    .X(_08828_));
 sky130_fd_sc_hd__a2bb2o_1 _24732_ (.A1_N(_08813_),
    .A2_N(_08828_),
    .B1(_08813_),
    .B2(_08828_),
    .X(_08829_));
 sky130_fd_sc_hd__o22a_1 _24733_ (.A1(_08682_),
    .A2(_08690_),
    .B1(_08681_),
    .B2(_08691_),
    .X(_08830_));
 sky130_fd_sc_hd__o22a_1 _24734_ (.A1(_08712_),
    .A2(_08713_),
    .B1(_08706_),
    .B2(_08714_),
    .X(_08831_));
 sky130_fd_sc_hd__a21oi_1 _24735_ (.A1(_08688_),
    .A2(_08689_),
    .B1(_08687_),
    .Y(_08832_));
 sky130_fd_sc_hd__o21ba_1 _24736_ (.A1(_08702_),
    .A2(_08705_),
    .B1_N(_08704_),
    .X(_08833_));
 sky130_fd_sc_hd__o22a_1 _24737_ (.A1(_08049_),
    .A2(_07595_),
    .B1(_08518_),
    .B2(_07873_),
    .X(_08834_));
 sky130_fd_sc_hd__and4_1 _24738_ (.A(_13149_),
    .B(_13519_),
    .C(_13155_),
    .D(_13515_),
    .X(_08835_));
 sky130_fd_sc_hd__nor2_2 _24739_ (.A(_08834_),
    .B(_08835_),
    .Y(_08836_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _24740_ (.A(_07889_),
    .X(_08837_));
 sky130_fd_sc_hd__buf_1 _24741_ (.A(_08837_),
    .X(_08838_));
 sky130_fd_sc_hd__buf_2 _24742_ (.A(_08838_),
    .X(_08839_));
 sky130_fd_sc_hd__nor2_2 _24743_ (.A(_05425_),
    .B(_08839_),
    .Y(_08840_));
 sky130_fd_sc_hd__a2bb2o_1 _24744_ (.A1_N(_08836_),
    .A2_N(_08840_),
    .B1(_08836_),
    .B2(_08840_),
    .X(_08841_));
 sky130_fd_sc_hd__a2bb2o_1 _24745_ (.A1_N(_08833_),
    .A2_N(_08841_),
    .B1(_08833_),
    .B2(_08841_),
    .X(_08842_));
 sky130_fd_sc_hd__a2bb2o_1 _24746_ (.A1_N(_08832_),
    .A2_N(_08842_),
    .B1(_08832_),
    .B2(_08842_),
    .X(_08843_));
 sky130_fd_sc_hd__a2bb2o_1 _24747_ (.A1_N(_08831_),
    .A2_N(_08843_),
    .B1(_08831_),
    .B2(_08843_),
    .X(_08844_));
 sky130_fd_sc_hd__a2bb2o_1 _24748_ (.A1_N(_08830_),
    .A2_N(_08844_),
    .B1(_08830_),
    .B2(_08844_),
    .X(_08845_));
 sky130_fd_sc_hd__o22a_1 _24749_ (.A1(_08680_),
    .A2(_08692_),
    .B1(_08679_),
    .B2(_08693_),
    .X(_08846_));
 sky130_fd_sc_hd__a2bb2o_1 _24750_ (.A1_N(_08845_),
    .A2_N(_08846_),
    .B1(_08845_),
    .B2(_08846_),
    .X(_08847_));
 sky130_fd_sc_hd__a2bb2o_2 _24751_ (.A1_N(_08829_),
    .A2_N(_08847_),
    .B1(_08829_),
    .B2(_08847_),
    .X(_08848_));
 sky130_fd_sc_hd__a2bb2o_1 _24752_ (.A1_N(_08811_),
    .A2_N(_08848_),
    .B1(_08811_),
    .B2(_08848_),
    .X(_08849_));
 sky130_fd_sc_hd__a2bb2o_1 _24753_ (.A1_N(_08810_),
    .A2_N(_08849_),
    .B1(_08810_),
    .B2(_08849_),
    .X(_08850_));
 sky130_fd_sc_hd__o22a_1 _24754_ (.A1(_08726_),
    .A2(_08727_),
    .B1(_08715_),
    .B2(_08728_),
    .X(_08851_));
 sky130_fd_sc_hd__o22a_1 _24755_ (.A1(_08733_),
    .A2(_08753_),
    .B1(_08732_),
    .B2(_08754_),
    .X(_08852_));
 sky130_fd_sc_hd__or2_1 _24756_ (.A(_08535_),
    .B(_07733_),
    .X(_08853_));
 sky130_fd_sc_hd__o22a_1 _24757_ (.A1(_08537_),
    .A2(_07196_),
    .B1(_08538_),
    .B2(_08364_),
    .X(_08854_));
 sky130_fd_sc_hd__and4_1 _24758_ (.A(_13137_),
    .B(_13534_),
    .C(_13143_),
    .D(_07448_),
    .X(_08855_));
 sky130_fd_sc_hd__or2_1 _24759_ (.A(_08854_),
    .B(_08855_),
    .X(_08856_));
 sky130_fd_sc_hd__a2bb2o_1 _24760_ (.A1_N(_08853_),
    .A2_N(_08856_),
    .B1(_08853_),
    .B2(_08856_),
    .X(_08857_));
 sky130_fd_sc_hd__clkbuf_2 _24761_ (.A(_05794_),
    .X(_08858_));
 sky130_fd_sc_hd__or2_1 _24762_ (.A(_08858_),
    .B(_07458_),
    .X(_08859_));
 sky130_fd_sc_hd__o22a_1 _24763_ (.A1(_08544_),
    .A2(_07905_),
    .B1(_08545_),
    .B2(_08050_),
    .X(_08860_));
 sky130_fd_sc_hd__and4_1 _24764_ (.A(_08547_),
    .B(_07907_),
    .C(_08548_),
    .D(_07908_),
    .X(_08861_));
 sky130_fd_sc_hd__or2_1 _24765_ (.A(_08860_),
    .B(_08861_),
    .X(_08862_));
 sky130_fd_sc_hd__a2bb2o_1 _24766_ (.A1_N(_08859_),
    .A2_N(_08862_),
    .B1(_08859_),
    .B2(_08862_),
    .X(_08863_));
 sky130_fd_sc_hd__o21ba_1 _24767_ (.A1(_08707_),
    .A2(_08711_),
    .B1_N(_08710_),
    .X(_08864_));
 sky130_fd_sc_hd__a2bb2o_1 _24768_ (.A1_N(_08863_),
    .A2_N(_08864_),
    .B1(_08863_),
    .B2(_08864_),
    .X(_08865_));
 sky130_fd_sc_hd__a2bb2o_2 _24769_ (.A1_N(_08857_),
    .A2_N(_08865_),
    .B1(_08857_),
    .B2(_08865_),
    .X(_08866_));
 sky130_fd_sc_hd__o21ba_1 _24770_ (.A1(_08718_),
    .A2(_08723_),
    .B1_N(_08722_),
    .X(_08867_));
 sky130_fd_sc_hd__o21ba_1 _24771_ (.A1(_08735_),
    .A2(_08740_),
    .B1_N(_08739_),
    .X(_08868_));
 sky130_fd_sc_hd__clkbuf_2 _24772_ (.A(_07253_),
    .X(_08869_));
 sky130_fd_sc_hd__clkbuf_2 _24773_ (.A(_06093_),
    .X(_08870_));
 sky130_fd_sc_hd__o22a_1 _24774_ (.A1(_08869_),
    .A2(_06451_),
    .B1(_08870_),
    .B2(_07780_),
    .X(_08871_));
 sky130_fd_sc_hd__buf_1 _24775_ (.A(_07798_),
    .X(_08872_));
 sky130_fd_sc_hd__buf_1 _24776_ (.A(_07799_),
    .X(_08873_));
 sky130_fd_sc_hd__and4_2 _24777_ (.A(_08872_),
    .B(_06901_),
    .C(_08873_),
    .D(_07040_),
    .X(_08874_));
 sky130_fd_sc_hd__nor2_2 _24778_ (.A(_08871_),
    .B(_08874_),
    .Y(_08875_));
 sky130_fd_sc_hd__nor2_2 _24779_ (.A(_06000_),
    .B(_06755_),
    .Y(_08876_));
 sky130_fd_sc_hd__a2bb2o_2 _24780_ (.A1_N(_08875_),
    .A2_N(_08876_),
    .B1(_08875_),
    .B2(_08876_),
    .X(_08877_));
 sky130_fd_sc_hd__a2bb2o_1 _24781_ (.A1_N(_08868_),
    .A2_N(_08877_),
    .B1(_08868_),
    .B2(_08877_),
    .X(_08878_));
 sky130_fd_sc_hd__a2bb2o_1 _24782_ (.A1_N(_08867_),
    .A2_N(_08878_),
    .B1(_08867_),
    .B2(_08878_),
    .X(_08879_));
 sky130_fd_sc_hd__o22a_1 _24783_ (.A1(_08717_),
    .A2(_08724_),
    .B1(_08716_),
    .B2(_08725_),
    .X(_08880_));
 sky130_fd_sc_hd__a2bb2o_1 _24784_ (.A1_N(_08879_),
    .A2_N(_08880_),
    .B1(_08879_),
    .B2(_08880_),
    .X(_08881_));
 sky130_fd_sc_hd__a2bb2o_1 _24785_ (.A1_N(_08866_),
    .A2_N(_08881_),
    .B1(_08866_),
    .B2(_08881_),
    .X(_08882_));
 sky130_fd_sc_hd__a2bb2o_1 _24786_ (.A1_N(_08852_),
    .A2_N(_08882_),
    .B1(_08852_),
    .B2(_08882_),
    .X(_08883_));
 sky130_fd_sc_hd__a2bb2o_1 _24787_ (.A1_N(_08851_),
    .A2_N(_08883_),
    .B1(_08851_),
    .B2(_08883_),
    .X(_08884_));
 sky130_fd_sc_hd__o22a_1 _24788_ (.A1(_08750_),
    .A2(_08751_),
    .B1(_08741_),
    .B2(_08752_),
    .X(_08885_));
 sky130_fd_sc_hd__o22a_1 _24789_ (.A1(_08757_),
    .A2(_08764_),
    .B1(_08756_),
    .B2(_08765_),
    .X(_08886_));
 sky130_fd_sc_hd__clkbuf_2 _24790_ (.A(_08559_),
    .X(_08887_));
 sky130_fd_sc_hd__or2_1 _24791_ (.A(_08734_),
    .B(_08887_),
    .X(_08888_));
 sky130_fd_sc_hd__clkbuf_2 _24792_ (.A(_07081_),
    .X(_08889_));
 sky130_fd_sc_hd__buf_2 _24793_ (.A(_06328_),
    .X(_08890_));
 sky130_fd_sc_hd__o22a_1 _24794_ (.A1(_08889_),
    .A2(_06921_),
    .B1(_08736_),
    .B2(_08890_),
    .X(_08891_));
 sky130_fd_sc_hd__and4_1 _24795_ (.A(_13106_),
    .B(_08738_),
    .C(_13112_),
    .D(_13564_),
    .X(_08892_));
 sky130_fd_sc_hd__or2_1 _24796_ (.A(_08891_),
    .B(_08892_),
    .X(_08893_));
 sky130_fd_sc_hd__a2bb2o_1 _24797_ (.A1_N(_08888_),
    .A2_N(_08893_),
    .B1(_08888_),
    .B2(_08893_),
    .X(_08894_));
 sky130_fd_sc_hd__buf_2 _24798_ (.A(_07663_),
    .X(_08895_));
 sky130_fd_sc_hd__or2_1 _24799_ (.A(_08895_),
    .B(_06334_),
    .X(_08896_));
 sky130_fd_sc_hd__clkbuf_2 _24800_ (.A(_08261_),
    .X(_08897_));
 sky130_fd_sc_hd__o22a_1 _24801_ (.A1(_08897_),
    .A2(_05931_),
    .B1(_06806_),
    .B2(_08417_),
    .X(_08898_));
 sky130_fd_sc_hd__and4_1 _24802_ (.A(_08745_),
    .B(_08747_),
    .C(_08746_),
    .D(_08419_),
    .X(_08899_));
 sky130_fd_sc_hd__or2_1 _24803_ (.A(_08898_),
    .B(_08899_),
    .X(_08900_));
 sky130_fd_sc_hd__a2bb2o_1 _24804_ (.A1_N(_08896_),
    .A2_N(_08900_),
    .B1(_08896_),
    .B2(_08900_),
    .X(_08901_));
 sky130_fd_sc_hd__o21ba_1 _24805_ (.A1(_08742_),
    .A2(_08749_),
    .B1_N(_08748_),
    .X(_08902_));
 sky130_fd_sc_hd__a2bb2o_1 _24806_ (.A1_N(_08901_),
    .A2_N(_08902_),
    .B1(_08901_),
    .B2(_08902_),
    .X(_08903_));
 sky130_fd_sc_hd__a2bb2o_1 _24807_ (.A1_N(_08894_),
    .A2_N(_08903_),
    .B1(_08894_),
    .B2(_08903_),
    .X(_08904_));
 sky130_fd_sc_hd__a2bb2o_1 _24808_ (.A1_N(_08886_),
    .A2_N(_08904_),
    .B1(_08886_),
    .B2(_08904_),
    .X(_08905_));
 sky130_fd_sc_hd__a2bb2o_1 _24809_ (.A1_N(_08885_),
    .A2_N(_08905_),
    .B1(_08885_),
    .B2(_08905_),
    .X(_08906_));
 sky130_fd_sc_hd__o21ba_1 _24810_ (.A1(_08759_),
    .A2(_08763_),
    .B1_N(_08762_),
    .X(_08907_));
 sky130_fd_sc_hd__o21ba_1 _24811_ (.A1(_08767_),
    .A2(_08770_),
    .B1_N(_08769_),
    .X(_08908_));
 sky130_fd_sc_hd__or2_1 _24812_ (.A(_07273_),
    .B(_05821_),
    .X(_08909_));
 sky130_fd_sc_hd__o22a_1 _24813_ (.A1(_08600_),
    .A2(_05723_),
    .B1(_08601_),
    .B2(_05725_),
    .X(_08910_));
 sky130_fd_sc_hd__and4_1 _24814_ (.A(_08603_),
    .B(_13588_),
    .C(_13092_),
    .D(_13585_),
    .X(_08911_));
 sky130_fd_sc_hd__or2_1 _24815_ (.A(_08910_),
    .B(_08911_),
    .X(_08912_));
 sky130_fd_sc_hd__a2bb2o_1 _24816_ (.A1_N(_08909_),
    .A2_N(_08912_),
    .B1(_08909_),
    .B2(_08912_),
    .X(_08913_));
 sky130_fd_sc_hd__a2bb2o_1 _24817_ (.A1_N(_08908_),
    .A2_N(_08913_),
    .B1(_08908_),
    .B2(_08913_),
    .X(_08914_));
 sky130_fd_sc_hd__a2bb2o_1 _24818_ (.A1_N(_08907_),
    .A2_N(_08914_),
    .B1(_08907_),
    .B2(_08914_),
    .X(_08915_));
 sky130_fd_sc_hd__or2_1 _24819_ (.A(_07531_),
    .B(_05731_),
    .X(_08916_));
 sky130_fd_sc_hd__o22a_1 _24820_ (.A1(_08448_),
    .A2(_06099_),
    .B1(_08449_),
    .B2(_08439_),
    .X(_08917_));
 sky130_fd_sc_hd__and4_1 _24821_ (.A(_08451_),
    .B(_13599_),
    .C(_08614_),
    .D(_13595_),
    .X(_08918_));
 sky130_fd_sc_hd__or2_1 _24822_ (.A(_08917_),
    .B(_08918_),
    .X(_08919_));
 sky130_fd_sc_hd__a2bb2o_1 _24823_ (.A1_N(_08916_),
    .A2_N(_08919_),
    .B1(_08916_),
    .B2(_08919_),
    .X(_08920_));
 sky130_fd_sc_hd__buf_1 _24824_ (.A(_07970_),
    .X(_08921_));
 sky130_fd_sc_hd__or2_1 _24825_ (.A(_08921_),
    .B(_07079_),
    .X(_08922_));
 sky130_fd_sc_hd__buf_1 _24826_ (.A(_08457_),
    .X(_08923_));
 sky130_fd_sc_hd__and4_1 _24827_ (.A(_08774_),
    .B(_07082_),
    .C(_08923_),
    .D(_13608_),
    .X(_08924_));
 sky130_fd_sc_hd__buf_1 _24828_ (.A(_11716_),
    .X(_08925_));
 sky130_fd_sc_hd__clkbuf_2 _24829_ (.A(_08130_),
    .X(_08926_));
 sky130_fd_sc_hd__o22a_1 _24830_ (.A1(_08925_),
    .A2(_13613_),
    .B1(_08926_),
    .B2(_05866_),
    .X(_08927_));
 sky130_fd_sc_hd__or2_1 _24831_ (.A(_08924_),
    .B(_08927_),
    .X(_08928_));
 sky130_fd_sc_hd__a2bb2o_1 _24832_ (.A1_N(_08922_),
    .A2_N(_08928_),
    .B1(_08922_),
    .B2(_08928_),
    .X(_08929_));
 sky130_fd_sc_hd__o21ba_1 _24833_ (.A1(_08773_),
    .A2(_08780_),
    .B1_N(_08776_),
    .X(_08930_));
 sky130_fd_sc_hd__a2bb2o_1 _24834_ (.A1_N(_08929_),
    .A2_N(_08930_),
    .B1(_08929_),
    .B2(_08930_),
    .X(_08931_));
 sky130_fd_sc_hd__a2bb2o_1 _24835_ (.A1_N(_08920_),
    .A2_N(_08931_),
    .B1(_08920_),
    .B2(_08931_),
    .X(_08932_));
 sky130_fd_sc_hd__o22a_1 _24836_ (.A1(_08781_),
    .A2(_08782_),
    .B1(_08771_),
    .B2(_08783_),
    .X(_08933_));
 sky130_fd_sc_hd__a2bb2o_1 _24837_ (.A1_N(_08932_),
    .A2_N(_08933_),
    .B1(_08932_),
    .B2(_08933_),
    .X(_08934_));
 sky130_fd_sc_hd__a2bb2o_1 _24838_ (.A1_N(_08915_),
    .A2_N(_08934_),
    .B1(_08915_),
    .B2(_08934_),
    .X(_08935_));
 sky130_fd_sc_hd__o22a_1 _24839_ (.A1(_08784_),
    .A2(_08785_),
    .B1(_08766_),
    .B2(_08786_),
    .X(_08936_));
 sky130_fd_sc_hd__a2bb2o_1 _24840_ (.A1_N(_08935_),
    .A2_N(_08936_),
    .B1(_08935_),
    .B2(_08936_),
    .X(_08937_));
 sky130_fd_sc_hd__a2bb2o_1 _24841_ (.A1_N(_08906_),
    .A2_N(_08937_),
    .B1(_08906_),
    .B2(_08937_),
    .X(_08938_));
 sky130_fd_sc_hd__o22a_1 _24842_ (.A1(_08787_),
    .A2(_08788_),
    .B1(_08755_),
    .B2(_08789_),
    .X(_08939_));
 sky130_fd_sc_hd__a2bb2o_1 _24843_ (.A1_N(_08938_),
    .A2_N(_08939_),
    .B1(_08938_),
    .B2(_08939_),
    .X(_08940_));
 sky130_fd_sc_hd__a2bb2o_1 _24844_ (.A1_N(_08884_),
    .A2_N(_08940_),
    .B1(_08884_),
    .B2(_08940_),
    .X(_08941_));
 sky130_fd_sc_hd__o22a_1 _24845_ (.A1(_08790_),
    .A2(_08791_),
    .B1(_08731_),
    .B2(_08792_),
    .X(_08942_));
 sky130_fd_sc_hd__a2bb2o_1 _24846_ (.A1_N(_08941_),
    .A2_N(_08942_),
    .B1(_08941_),
    .B2(_08942_),
    .X(_08943_));
 sky130_fd_sc_hd__a2bb2o_1 _24847_ (.A1_N(_08850_),
    .A2_N(_08943_),
    .B1(_08850_),
    .B2(_08943_),
    .X(_08944_));
 sky130_fd_sc_hd__o22a_1 _24848_ (.A1(_08793_),
    .A2(_08794_),
    .B1(_08699_),
    .B2(_08795_),
    .X(_08945_));
 sky130_fd_sc_hd__a2bb2o_1 _24849_ (.A1_N(_08944_),
    .A2_N(_08945_),
    .B1(_08944_),
    .B2(_08945_),
    .X(_08946_));
 sky130_fd_sc_hd__a2bb2o_1 _24850_ (.A1_N(_08809_),
    .A2_N(_08946_),
    .B1(_08809_),
    .B2(_08946_),
    .X(_08947_));
 sky130_fd_sc_hd__o22a_1 _24851_ (.A1(_08796_),
    .A2(_08797_),
    .B1(_08656_),
    .B2(_08798_),
    .X(_08948_));
 sky130_fd_sc_hd__a2bb2o_1 _24852_ (.A1_N(_08947_),
    .A2_N(_08948_),
    .B1(_08947_),
    .B2(_08948_),
    .X(_08949_));
 sky130_fd_sc_hd__a2bb2o_1 _24853_ (.A1_N(_08655_),
    .A2_N(_08949_),
    .B1(_08655_),
    .B2(_08949_),
    .X(_08950_));
 sky130_fd_sc_hd__o22a_1 _24854_ (.A1(_08799_),
    .A2(_08800_),
    .B1(_08488_),
    .B2(_08801_),
    .X(_08951_));
 sky130_fd_sc_hd__or2_2 _24855_ (.A(_08950_),
    .B(_08951_),
    .X(_08952_));
 sky130_fd_sc_hd__a21bo_1 _24856_ (.A1(_08950_),
    .A2(_08951_),
    .B1_N(_08952_),
    .X(_08953_));
 sky130_fd_sc_hd__clkbuf_2 _24857_ (.A(_08953_),
    .X(_08954_));
 sky130_fd_sc_hd__or2_1 _24858_ (.A(_08648_),
    .B(_08804_),
    .X(_08955_));
 sky130_fd_sc_hd__or3_4 _24859_ (.A(_08321_),
    .B(_08485_),
    .C(_08955_),
    .X(_08956_));
 sky130_fd_sc_hd__o21ai_1 _24860_ (.A1(_08652_),
    .A2(_08803_),
    .B1(_08647_),
    .Y(_08957_));
 sky130_fd_sc_hd__o221a_1 _24861_ (.A1(_08651_),
    .A2(_08802_),
    .B1(_08649_),
    .B2(_08955_),
    .C1(_08957_),
    .X(_08958_));
 sky130_fd_sc_hd__o21ai_1 _24862_ (.A1(_08328_),
    .A2(_08956_),
    .B1(_08958_),
    .Y(_08959_));
 sky130_vsdinv _24863_ (.A(_08959_),
    .Y(_08960_));
 sky130_vsdinv _24864_ (.A(_08954_),
    .Y(_08961_));
 sky130_fd_sc_hd__o22a_4 _24865_ (.A1(_08954_),
    .A2(_08960_),
    .B1(_08961_),
    .B2(_08959_),
    .X(_02655_));
 sky130_fd_sc_hd__o22a_1 _24866_ (.A1(_08947_),
    .A2(_08948_),
    .B1(_08655_),
    .B2(_08949_),
    .X(_08962_));
 sky130_fd_sc_hd__o22a_1 _24867_ (.A1(_08811_),
    .A2(_08848_),
    .B1(_08810_),
    .B2(_08849_),
    .X(_08963_));
 sky130_fd_sc_hd__buf_1 _24868_ (.A(_08813_),
    .X(_08964_));
 sky130_fd_sc_hd__buf_1 _24869_ (.A(_08964_),
    .X(_08965_));
 sky130_fd_sc_hd__o22a_2 _24870_ (.A1(_08826_),
    .A2(_08827_),
    .B1(_08965_),
    .B2(_08828_),
    .X(_08966_));
 sky130_fd_sc_hd__or2_1 _24871_ (.A(_08963_),
    .B(_08966_),
    .X(_08967_));
 sky130_fd_sc_hd__a21bo_1 _24872_ (.A1(_08963_),
    .A2(_08966_),
    .B1_N(_08967_),
    .X(_08968_));
 sky130_fd_sc_hd__o22a_2 _24873_ (.A1(_08845_),
    .A2(_08846_),
    .B1(_08829_),
    .B2(_08847_),
    .X(_08969_));
 sky130_fd_sc_hd__o22a_1 _24874_ (.A1(_08852_),
    .A2(_08882_),
    .B1(_08851_),
    .B2(_08883_),
    .X(_08970_));
 sky130_fd_sc_hd__buf_1 _24875_ (.A(_08664_),
    .X(_08971_));
 sky130_fd_sc_hd__o22a_1 _24876_ (.A1(_08818_),
    .A2(_08824_),
    .B1(_08971_),
    .B2(_08825_),
    .X(_08972_));
 sky130_fd_sc_hd__or4_4 _24877_ (.A(_08661_),
    .B(_07184_),
    .C(_08661_),
    .D(_07182_),
    .X(_08973_));
 sky130_fd_sc_hd__buf_1 _24878_ (.A(_08815_),
    .X(_08974_));
 sky130_fd_sc_hd__a22o_1 _24879_ (.A1(_08974_),
    .A2(_13168_),
    .B1(_08974_),
    .B2(_13162_),
    .X(_08975_));
 sky130_fd_sc_hd__nand2_1 _24880_ (.A(_08973_),
    .B(_08975_),
    .Y(_08976_));
 sky130_fd_sc_hd__o22a_1 _24881_ (.A1(_08353_),
    .A2(_08821_),
    .B1(_05144_),
    .B2(_08819_),
    .X(_08977_));
 sky130_fd_sc_hd__a2bb2o_2 _24882_ (.A1_N(_08976_),
    .A2_N(_08977_),
    .B1(_08976_),
    .B2(_08977_),
    .X(_08978_));
 sky130_fd_sc_hd__nor2_1 _24883_ (.A(_08971_),
    .B(_08978_),
    .Y(_08979_));
 sky130_fd_sc_hd__a21oi_2 _24884_ (.A1(_08971_),
    .A2(_08978_),
    .B1(_08979_),
    .Y(_08980_));
 sky130_fd_sc_hd__o2bb2ai_1 _24885_ (.A1_N(_08972_),
    .A2_N(_08980_),
    .B1(_08972_),
    .B2(_08980_),
    .Y(_08981_));
 sky130_fd_sc_hd__a2bb2o_1 _24886_ (.A1_N(_08964_),
    .A2_N(_08981_),
    .B1(_08813_),
    .B2(_08981_),
    .X(_08982_));
 sky130_fd_sc_hd__o22a_1 _24887_ (.A1(_08833_),
    .A2(_08841_),
    .B1(_08832_),
    .B2(_08842_),
    .X(_08983_));
 sky130_fd_sc_hd__o22a_1 _24888_ (.A1(_08863_),
    .A2(_08864_),
    .B1(_08857_),
    .B2(_08865_),
    .X(_08984_));
 sky130_fd_sc_hd__a21oi_2 _24889_ (.A1(_08836_),
    .A2(_08840_),
    .B1(_08835_),
    .Y(_08985_));
 sky130_fd_sc_hd__o21ba_1 _24890_ (.A1(_08853_),
    .A2(_08856_),
    .B1_N(_08855_),
    .X(_08986_));
 sky130_fd_sc_hd__o22a_1 _24891_ (.A1(_08683_),
    .A2(_07873_),
    .B1(_08518_),
    .B2(_08838_),
    .X(_08987_));
 sky130_fd_sc_hd__and4_1 _24892_ (.A(_13149_),
    .B(_08023_),
    .C(_13155_),
    .D(_13510_),
    .X(_08988_));
 sky130_fd_sc_hd__nor2_2 _24893_ (.A(_08987_),
    .B(_08988_),
    .Y(_08989_));
 sky130_fd_sc_hd__nor2_2 _24894_ (.A(_05425_),
    .B(_08498_),
    .Y(_08990_));
 sky130_fd_sc_hd__a2bb2o_1 _24895_ (.A1_N(_08989_),
    .A2_N(_08990_),
    .B1(_08989_),
    .B2(_08990_),
    .X(_08991_));
 sky130_fd_sc_hd__a2bb2o_1 _24896_ (.A1_N(_08986_),
    .A2_N(_08991_),
    .B1(_08986_),
    .B2(_08991_),
    .X(_08992_));
 sky130_fd_sc_hd__a2bb2o_1 _24897_ (.A1_N(_08985_),
    .A2_N(_08992_),
    .B1(_08985_),
    .B2(_08992_),
    .X(_08993_));
 sky130_fd_sc_hd__a2bb2o_1 _24898_ (.A1_N(_08984_),
    .A2_N(_08993_),
    .B1(_08984_),
    .B2(_08993_),
    .X(_08994_));
 sky130_fd_sc_hd__a2bb2o_1 _24899_ (.A1_N(_08983_),
    .A2_N(_08994_),
    .B1(_08983_),
    .B2(_08994_),
    .X(_08995_));
 sky130_fd_sc_hd__o22a_1 _24900_ (.A1(_08831_),
    .A2(_08843_),
    .B1(_08830_),
    .B2(_08844_),
    .X(_08996_));
 sky130_fd_sc_hd__a2bb2o_1 _24901_ (.A1_N(_08995_),
    .A2_N(_08996_),
    .B1(_08995_),
    .B2(_08996_),
    .X(_08997_));
 sky130_fd_sc_hd__a2bb2o_2 _24902_ (.A1_N(_08982_),
    .A2_N(_08997_),
    .B1(_08982_),
    .B2(_08997_),
    .X(_08998_));
 sky130_fd_sc_hd__a2bb2o_1 _24903_ (.A1_N(_08970_),
    .A2_N(_08998_),
    .B1(_08970_),
    .B2(_08998_),
    .X(_08999_));
 sky130_fd_sc_hd__a2bb2o_1 _24904_ (.A1_N(_08969_),
    .A2_N(_08999_),
    .B1(_08969_),
    .B2(_08999_),
    .X(_09000_));
 sky130_fd_sc_hd__o22a_1 _24905_ (.A1(_08879_),
    .A2(_08880_),
    .B1(_08866_),
    .B2(_08881_),
    .X(_09001_));
 sky130_fd_sc_hd__o22a_1 _24906_ (.A1(_08886_),
    .A2(_08904_),
    .B1(_08885_),
    .B2(_08905_),
    .X(_09002_));
 sky130_fd_sc_hd__clkbuf_2 _24907_ (.A(_08217_),
    .X(_09003_));
 sky130_fd_sc_hd__o22a_1 _24908_ (.A1(_09003_),
    .A2(_07326_),
    .B1(_05589_),
    .B2(_08178_),
    .X(_09004_));
 sky130_fd_sc_hd__and4_1 _24909_ (.A(_13138_),
    .B(_13529_),
    .C(_13144_),
    .D(_08686_),
    .X(_09005_));
 sky130_fd_sc_hd__nor2_2 _24910_ (.A(_09004_),
    .B(_09005_),
    .Y(_09006_));
 sky130_fd_sc_hd__buf_2 _24911_ (.A(_08180_),
    .X(_09007_));
 sky130_fd_sc_hd__nor2_2 _24912_ (.A(_05538_),
    .B(_09007_),
    .Y(_09008_));
 sky130_fd_sc_hd__a2bb2o_1 _24913_ (.A1_N(_09006_),
    .A2_N(_09008_),
    .B1(_09006_),
    .B2(_09008_),
    .X(_09009_));
 sky130_fd_sc_hd__or2_1 _24914_ (.A(_08858_),
    .B(_07197_),
    .X(_09010_));
 sky130_fd_sc_hd__clkbuf_2 _24915_ (.A(_06710_),
    .X(_09011_));
 sky130_fd_sc_hd__o22a_1 _24916_ (.A1(_09011_),
    .A2(_08050_),
    .B1(_08545_),
    .B2(_07457_),
    .X(_09012_));
 sky130_fd_sc_hd__and4_1 _24917_ (.A(_13130_),
    .B(_07908_),
    .C(_13133_),
    .D(_08200_),
    .X(_09013_));
 sky130_fd_sc_hd__or2_1 _24918_ (.A(_09012_),
    .B(_09013_),
    .X(_09014_));
 sky130_fd_sc_hd__a2bb2o_1 _24919_ (.A1_N(_09010_),
    .A2_N(_09014_),
    .B1(_09010_),
    .B2(_09014_),
    .X(_09015_));
 sky130_fd_sc_hd__o21ba_1 _24920_ (.A1(_08859_),
    .A2(_08862_),
    .B1_N(_08861_),
    .X(_09016_));
 sky130_fd_sc_hd__a2bb2o_1 _24921_ (.A1_N(_09015_),
    .A2_N(_09016_),
    .B1(_09015_),
    .B2(_09016_),
    .X(_09017_));
 sky130_fd_sc_hd__a2bb2o_2 _24922_ (.A1_N(_09009_),
    .A2_N(_09017_),
    .B1(_09009_),
    .B2(_09017_),
    .X(_09018_));
 sky130_fd_sc_hd__a21oi_2 _24923_ (.A1(_08875_),
    .A2(_08876_),
    .B1(_08874_),
    .Y(_09019_));
 sky130_fd_sc_hd__o21ba_1 _24924_ (.A1(_08888_),
    .A2(_08893_),
    .B1_N(_08892_),
    .X(_09020_));
 sky130_fd_sc_hd__clkbuf_4 _24925_ (.A(_07383_),
    .X(_09021_));
 sky130_fd_sc_hd__o22a_1 _24926_ (.A1(_09021_),
    .A2(_06575_),
    .B1(_06090_),
    .B2(_06754_),
    .X(_09022_));
 sky130_fd_sc_hd__and4_2 _24927_ (.A(_13119_),
    .B(_13553_),
    .C(_13123_),
    .D(_07329_),
    .X(_09023_));
 sky130_fd_sc_hd__nor2_2 _24928_ (.A(_09022_),
    .B(_09023_),
    .Y(_09024_));
 sky130_fd_sc_hd__clkbuf_4 _24929_ (.A(_06881_),
    .X(_09025_));
 sky130_fd_sc_hd__nor2_2 _24930_ (.A(_06000_),
    .B(_09025_),
    .Y(_09026_));
 sky130_fd_sc_hd__a2bb2o_1 _24931_ (.A1_N(_09024_),
    .A2_N(_09026_),
    .B1(_09024_),
    .B2(_09026_),
    .X(_09027_));
 sky130_fd_sc_hd__a2bb2o_1 _24932_ (.A1_N(_09020_),
    .A2_N(_09027_),
    .B1(_09020_),
    .B2(_09027_),
    .X(_09028_));
 sky130_fd_sc_hd__a2bb2o_1 _24933_ (.A1_N(_09019_),
    .A2_N(_09028_),
    .B1(_09019_),
    .B2(_09028_),
    .X(_09029_));
 sky130_fd_sc_hd__o22a_1 _24934_ (.A1(_08868_),
    .A2(_08877_),
    .B1(_08867_),
    .B2(_08878_),
    .X(_09030_));
 sky130_fd_sc_hd__a2bb2o_1 _24935_ (.A1_N(_09029_),
    .A2_N(_09030_),
    .B1(_09029_),
    .B2(_09030_),
    .X(_09031_));
 sky130_fd_sc_hd__a2bb2o_1 _24936_ (.A1_N(_09018_),
    .A2_N(_09031_),
    .B1(_09018_),
    .B2(_09031_),
    .X(_09032_));
 sky130_fd_sc_hd__a2bb2o_1 _24937_ (.A1_N(_09002_),
    .A2_N(_09032_),
    .B1(_09002_),
    .B2(_09032_),
    .X(_09033_));
 sky130_fd_sc_hd__a2bb2o_2 _24938_ (.A1_N(_09001_),
    .A2_N(_09033_),
    .B1(_09001_),
    .B2(_09033_),
    .X(_09034_));
 sky130_fd_sc_hd__o22a_1 _24939_ (.A1(_08901_),
    .A2(_08902_),
    .B1(_08894_),
    .B2(_08903_),
    .X(_09035_));
 sky130_fd_sc_hd__o22a_1 _24940_ (.A1(_08908_),
    .A2(_08913_),
    .B1(_08907_),
    .B2(_08914_),
    .X(_09036_));
 sky130_fd_sc_hd__or2_1 _24941_ (.A(_06285_),
    .B(_08557_),
    .X(_09037_));
 sky130_fd_sc_hd__o22a_1 _24942_ (.A1(_08574_),
    .A2(_06916_),
    .B1(_08575_),
    .B2(_08559_),
    .X(_09038_));
 sky130_fd_sc_hd__and4_1 _24943_ (.A(_08577_),
    .B(_13564_),
    .C(_08578_),
    .D(_07212_),
    .X(_09039_));
 sky130_fd_sc_hd__or2_1 _24944_ (.A(_09038_),
    .B(_09039_),
    .X(_09040_));
 sky130_fd_sc_hd__a2bb2o_1 _24945_ (.A1_N(_09037_),
    .A2_N(_09040_),
    .B1(_09037_),
    .B2(_09040_),
    .X(_09041_));
 sky130_fd_sc_hd__or2_1 _24946_ (.A(_08895_),
    .B(_06327_),
    .X(_09042_));
 sky130_fd_sc_hd__o22a_1 _24947_ (.A1(_08743_),
    .A2(_06031_),
    .B1(_06806_),
    .B2(_08234_),
    .X(_09043_));
 sky130_fd_sc_hd__and4_1 _24948_ (.A(_08585_),
    .B(_08419_),
    .C(_08586_),
    .D(_08237_),
    .X(_09044_));
 sky130_fd_sc_hd__or2_1 _24949_ (.A(_09043_),
    .B(_09044_),
    .X(_09045_));
 sky130_fd_sc_hd__a2bb2o_1 _24950_ (.A1_N(_09042_),
    .A2_N(_09045_),
    .B1(_09042_),
    .B2(_09045_),
    .X(_09046_));
 sky130_fd_sc_hd__o21ba_1 _24951_ (.A1(_08896_),
    .A2(_08900_),
    .B1_N(_08899_),
    .X(_09047_));
 sky130_fd_sc_hd__a2bb2o_1 _24952_ (.A1_N(_09046_),
    .A2_N(_09047_),
    .B1(_09046_),
    .B2(_09047_),
    .X(_09048_));
 sky130_fd_sc_hd__a2bb2o_1 _24953_ (.A1_N(_09041_),
    .A2_N(_09048_),
    .B1(_09041_),
    .B2(_09048_),
    .X(_09049_));
 sky130_fd_sc_hd__a2bb2o_1 _24954_ (.A1_N(_09036_),
    .A2_N(_09049_),
    .B1(_09036_),
    .B2(_09049_),
    .X(_09050_));
 sky130_fd_sc_hd__a2bb2o_1 _24955_ (.A1_N(_09035_),
    .A2_N(_09050_),
    .B1(_09035_),
    .B2(_09050_),
    .X(_09051_));
 sky130_fd_sc_hd__o21ba_1 _24956_ (.A1(_08909_),
    .A2(_08912_),
    .B1_N(_08911_),
    .X(_09052_));
 sky130_fd_sc_hd__o21ba_1 _24957_ (.A1(_08916_),
    .A2(_08919_),
    .B1_N(_08918_),
    .X(_09053_));
 sky130_fd_sc_hd__or2_1 _24958_ (.A(_07273_),
    .B(_05932_),
    .X(_09054_));
 sky130_fd_sc_hd__o22a_1 _24959_ (.A1(_08600_),
    .A2(_08425_),
    .B1(_08601_),
    .B2(_05820_),
    .X(_09055_));
 sky130_fd_sc_hd__and4_1 _24960_ (.A(_08603_),
    .B(_08427_),
    .C(_08441_),
    .D(_08587_),
    .X(_09056_));
 sky130_fd_sc_hd__or2_1 _24961_ (.A(_09055_),
    .B(_09056_),
    .X(_09057_));
 sky130_fd_sc_hd__a2bb2o_1 _24962_ (.A1_N(_09054_),
    .A2_N(_09057_),
    .B1(_09054_),
    .B2(_09057_),
    .X(_09058_));
 sky130_fd_sc_hd__a2bb2o_1 _24963_ (.A1_N(_09053_),
    .A2_N(_09058_),
    .B1(_09053_),
    .B2(_09058_),
    .X(_09059_));
 sky130_fd_sc_hd__a2bb2o_1 _24964_ (.A1_N(_09052_),
    .A2_N(_09059_),
    .B1(_09052_),
    .B2(_09059_),
    .X(_09060_));
 sky130_fd_sc_hd__or2_1 _24965_ (.A(_08609_),
    .B(_05831_),
    .X(_09061_));
 sky130_fd_sc_hd__o22a_1 _24966_ (.A1(_08286_),
    .A2(_05663_),
    .B1(_08287_),
    .B2(_07126_),
    .X(_09062_));
 sky130_fd_sc_hd__and4_1 _24967_ (.A(_08451_),
    .B(_07249_),
    .C(_08452_),
    .D(_07251_),
    .X(_09063_));
 sky130_fd_sc_hd__or2_1 _24968_ (.A(_09062_),
    .B(_09063_),
    .X(_09064_));
 sky130_fd_sc_hd__a2bb2o_1 _24969_ (.A1_N(_09061_),
    .A2_N(_09064_),
    .B1(_09061_),
    .B2(_09064_),
    .X(_09065_));
 sky130_fd_sc_hd__or2_1 _24970_ (.A(_08921_),
    .B(_05862_),
    .X(_09066_));
 sky130_fd_sc_hd__buf_1 _24971_ (.A(_08294_),
    .X(_09067_));
 sky130_fd_sc_hd__and4_1 _24972_ (.A(_09067_),
    .B(_05866_),
    .C(_08923_),
    .D(_05872_),
    .X(_09068_));
 sky130_fd_sc_hd__clkbuf_2 _24973_ (.A(_08130_),
    .X(_09069_));
 sky130_fd_sc_hd__o22a_1 _24974_ (.A1(_08925_),
    .A2(_07086_),
    .B1(_09069_),
    .B2(_05868_),
    .X(_09070_));
 sky130_fd_sc_hd__or2_1 _24975_ (.A(_09068_),
    .B(_09070_),
    .X(_09071_));
 sky130_fd_sc_hd__a2bb2o_1 _24976_ (.A1_N(_09066_),
    .A2_N(_09071_),
    .B1(_09066_),
    .B2(_09071_),
    .X(_09072_));
 sky130_fd_sc_hd__o21ba_1 _24977_ (.A1(_08922_),
    .A2(_08928_),
    .B1_N(_08924_),
    .X(_09073_));
 sky130_fd_sc_hd__a2bb2o_1 _24978_ (.A1_N(_09072_),
    .A2_N(_09073_),
    .B1(_09072_),
    .B2(_09073_),
    .X(_09074_));
 sky130_fd_sc_hd__a2bb2o_1 _24979_ (.A1_N(_09065_),
    .A2_N(_09074_),
    .B1(_09065_),
    .B2(_09074_),
    .X(_09075_));
 sky130_fd_sc_hd__o22a_1 _24980_ (.A1(_08929_),
    .A2(_08930_),
    .B1(_08920_),
    .B2(_08931_),
    .X(_09076_));
 sky130_fd_sc_hd__a2bb2o_1 _24981_ (.A1_N(_09075_),
    .A2_N(_09076_),
    .B1(_09075_),
    .B2(_09076_),
    .X(_09077_));
 sky130_fd_sc_hd__a2bb2o_1 _24982_ (.A1_N(_09060_),
    .A2_N(_09077_),
    .B1(_09060_),
    .B2(_09077_),
    .X(_09078_));
 sky130_fd_sc_hd__o22a_1 _24983_ (.A1(_08932_),
    .A2(_08933_),
    .B1(_08915_),
    .B2(_08934_),
    .X(_09079_));
 sky130_fd_sc_hd__a2bb2o_1 _24984_ (.A1_N(_09078_),
    .A2_N(_09079_),
    .B1(_09078_),
    .B2(_09079_),
    .X(_09080_));
 sky130_fd_sc_hd__a2bb2o_1 _24985_ (.A1_N(_09051_),
    .A2_N(_09080_),
    .B1(_09051_),
    .B2(_09080_),
    .X(_09081_));
 sky130_fd_sc_hd__o22a_1 _24986_ (.A1(_08935_),
    .A2(_08936_),
    .B1(_08906_),
    .B2(_08937_),
    .X(_09082_));
 sky130_fd_sc_hd__a2bb2o_1 _24987_ (.A1_N(_09081_),
    .A2_N(_09082_),
    .B1(_09081_),
    .B2(_09082_),
    .X(_09083_));
 sky130_fd_sc_hd__a2bb2o_1 _24988_ (.A1_N(_09034_),
    .A2_N(_09083_),
    .B1(_09034_),
    .B2(_09083_),
    .X(_09084_));
 sky130_fd_sc_hd__o22a_1 _24989_ (.A1(_08938_),
    .A2(_08939_),
    .B1(_08884_),
    .B2(_08940_),
    .X(_09085_));
 sky130_fd_sc_hd__a2bb2o_1 _24990_ (.A1_N(_09084_),
    .A2_N(_09085_),
    .B1(_09084_),
    .B2(_09085_),
    .X(_09086_));
 sky130_fd_sc_hd__a2bb2o_1 _24991_ (.A1_N(_09000_),
    .A2_N(_09086_),
    .B1(_09000_),
    .B2(_09086_),
    .X(_09087_));
 sky130_fd_sc_hd__o22a_1 _24992_ (.A1(_08941_),
    .A2(_08942_),
    .B1(_08850_),
    .B2(_08943_),
    .X(_09088_));
 sky130_fd_sc_hd__a2bb2o_1 _24993_ (.A1_N(_09087_),
    .A2_N(_09088_),
    .B1(_09087_),
    .B2(_09088_),
    .X(_09089_));
 sky130_fd_sc_hd__a2bb2o_1 _24994_ (.A1_N(_08968_),
    .A2_N(_09089_),
    .B1(_08968_),
    .B2(_09089_),
    .X(_09090_));
 sky130_fd_sc_hd__o22a_1 _24995_ (.A1(_08944_),
    .A2(_08945_),
    .B1(_08809_),
    .B2(_08946_),
    .X(_09091_));
 sky130_fd_sc_hd__a2bb2o_1 _24996_ (.A1_N(_09090_),
    .A2_N(_09091_),
    .B1(_09090_),
    .B2(_09091_),
    .X(_09092_));
 sky130_fd_sc_hd__a2bb2o_1 _24997_ (.A1_N(_08808_),
    .A2_N(_09092_),
    .B1(_08808_),
    .B2(_09092_),
    .X(_09093_));
 sky130_fd_sc_hd__or2_1 _24998_ (.A(_08962_),
    .B(_09093_),
    .X(_09094_));
 sky130_fd_sc_hd__a21bo_1 _24999_ (.A1(_08962_),
    .A2(_09093_),
    .B1_N(_09094_),
    .X(_09095_));
 sky130_fd_sc_hd__o21ai_2 _25000_ (.A1(_08954_),
    .A2(_08960_),
    .B1(_08952_),
    .Y(_09096_));
 sky130_fd_sc_hd__a2bb2o_4 _25001_ (.A1_N(_09095_),
    .A2_N(_09096_),
    .B1(_09095_),
    .B2(_09096_),
    .X(_02656_));
 sky130_fd_sc_hd__o22a_1 _25002_ (.A1(_08970_),
    .A2(_08998_),
    .B1(_08969_),
    .B2(_08999_),
    .X(_09097_));
 sky130_fd_sc_hd__o22a_2 _25003_ (.A1(_08972_),
    .A2(_08980_),
    .B1(_08965_),
    .B2(_08981_),
    .X(_09098_));
 sky130_fd_sc_hd__or2_1 _25004_ (.A(_09097_),
    .B(_09098_),
    .X(_09099_));
 sky130_fd_sc_hd__a21bo_1 _25005_ (.A1(_09097_),
    .A2(_09098_),
    .B1_N(_09099_),
    .X(_09100_));
 sky130_fd_sc_hd__o22a_2 _25006_ (.A1(_08995_),
    .A2(_08996_),
    .B1(_08982_),
    .B2(_08997_),
    .X(_09101_));
 sky130_fd_sc_hd__o22a_1 _25007_ (.A1(_09002_),
    .A2(_09032_),
    .B1(_09001_),
    .B2(_09033_),
    .X(_09102_));
 sky130_fd_sc_hd__or2_1 _25008_ (.A(_08347_),
    .B(_08975_),
    .X(_09103_));
 sky130_vsdinv _25009_ (.A(_09103_),
    .Y(_09104_));
 sky130_fd_sc_hd__o32a_1 _25010_ (.A1(_08971_),
    .A2(_08978_),
    .A3(_09103_),
    .B1(_08979_),
    .B2(_09104_),
    .X(_09105_));
 sky130_fd_sc_hd__a2bb2o_1 _25011_ (.A1_N(_08964_),
    .A2_N(_09105_),
    .B1(_08964_),
    .B2(_09105_),
    .X(_09106_));
 sky130_fd_sc_hd__o22a_1 _25012_ (.A1(_08986_),
    .A2(_08991_),
    .B1(_08985_),
    .B2(_08992_),
    .X(_09107_));
 sky130_fd_sc_hd__o22a_1 _25013_ (.A1(_09015_),
    .A2(_09016_),
    .B1(_09009_),
    .B2(_09017_),
    .X(_09108_));
 sky130_fd_sc_hd__a21oi_2 _25014_ (.A1(_08989_),
    .A2(_08990_),
    .B1(_08988_),
    .Y(_09109_));
 sky130_fd_sc_hd__a21oi_2 _25015_ (.A1(_09006_),
    .A2(_09008_),
    .B1(_09005_),
    .Y(_09110_));
 sky130_fd_sc_hd__o22a_1 _25016_ (.A1(_07055_),
    .A2(_08837_),
    .B1(_07214_),
    .B2(_08034_),
    .X(_09111_));
 sky130_fd_sc_hd__and4_1 _25017_ (.A(_13148_),
    .B(_08667_),
    .C(_13154_),
    .D(_08668_),
    .X(_09112_));
 sky130_fd_sc_hd__or2_1 _25018_ (.A(_09111_),
    .B(_09112_),
    .X(_09113_));
 sky130_vsdinv _25019_ (.A(_09113_),
    .Y(_09114_));
 sky130_fd_sc_hd__or2_1 _25020_ (.A(_11701_),
    .B(_05421_),
    .X(_09115_));
 sky130_fd_sc_hd__buf_1 _25021_ (.A(_09115_),
    .X(_09116_));
 sky130_fd_sc_hd__a32o_1 _25022_ (.A1(_08816_),
    .A2(\pcpi_mul.rs2[6] ),
    .A3(_09114_),
    .B1(_09113_),
    .B2(_09116_),
    .X(_09117_));
 sky130_fd_sc_hd__a2bb2o_1 _25023_ (.A1_N(_09110_),
    .A2_N(_09117_),
    .B1(_09110_),
    .B2(_09117_),
    .X(_09118_));
 sky130_fd_sc_hd__a2bb2o_1 _25024_ (.A1_N(_09109_),
    .A2_N(_09118_),
    .B1(_09109_),
    .B2(_09118_),
    .X(_09119_));
 sky130_fd_sc_hd__a2bb2o_1 _25025_ (.A1_N(_09108_),
    .A2_N(_09119_),
    .B1(_09108_),
    .B2(_09119_),
    .X(_09120_));
 sky130_fd_sc_hd__a2bb2o_1 _25026_ (.A1_N(_09107_),
    .A2_N(_09120_),
    .B1(_09107_),
    .B2(_09120_),
    .X(_09121_));
 sky130_fd_sc_hd__o22a_1 _25027_ (.A1(_08984_),
    .A2(_08993_),
    .B1(_08983_),
    .B2(_08994_),
    .X(_09122_));
 sky130_fd_sc_hd__a2bb2o_1 _25028_ (.A1_N(_09121_),
    .A2_N(_09122_),
    .B1(_09121_),
    .B2(_09122_),
    .X(_09123_));
 sky130_fd_sc_hd__a2bb2o_2 _25029_ (.A1_N(_09106_),
    .A2_N(_09123_),
    .B1(_09106_),
    .B2(_09123_),
    .X(_09124_));
 sky130_fd_sc_hd__a2bb2o_1 _25030_ (.A1_N(_09102_),
    .A2_N(_09124_),
    .B1(_09102_),
    .B2(_09124_),
    .X(_09125_));
 sky130_fd_sc_hd__a2bb2o_1 _25031_ (.A1_N(_09101_),
    .A2_N(_09125_),
    .B1(_09101_),
    .B2(_09125_),
    .X(_09126_));
 sky130_fd_sc_hd__o22a_1 _25032_ (.A1(_09029_),
    .A2(_09030_),
    .B1(_09018_),
    .B2(_09031_),
    .X(_09127_));
 sky130_fd_sc_hd__o22a_1 _25033_ (.A1(_09036_),
    .A2(_09049_),
    .B1(_09035_),
    .B2(_09050_),
    .X(_09128_));
 sky130_fd_sc_hd__o22a_1 _25034_ (.A1(_09003_),
    .A2(_08684_),
    .B1(_05589_),
    .B2(_08180_),
    .X(_09129_));
 sky130_fd_sc_hd__and4_1 _25035_ (.A(_13138_),
    .B(_08686_),
    .C(_13144_),
    .D(_07877_),
    .X(_09130_));
 sky130_fd_sc_hd__nor2_2 _25036_ (.A(_09129_),
    .B(_09130_),
    .Y(_09131_));
 sky130_fd_sc_hd__nor2_2 _25037_ (.A(_08535_),
    .B(_07874_),
    .Y(_09132_));
 sky130_fd_sc_hd__a2bb2o_1 _25038_ (.A1_N(_09131_),
    .A2_N(_09132_),
    .B1(_09131_),
    .B2(_09132_),
    .X(_09133_));
 sky130_fd_sc_hd__or2_1 _25039_ (.A(_08858_),
    .B(_07736_),
    .X(_09134_));
 sky130_fd_sc_hd__o22a_1 _25040_ (.A1(_09011_),
    .A2(_07032_),
    .B1(_08545_),
    .B2(_08198_),
    .X(_09135_));
 sky130_fd_sc_hd__and4_1 _25041_ (.A(_08547_),
    .B(_08200_),
    .C(_08548_),
    .D(_13534_),
    .X(_09136_));
 sky130_fd_sc_hd__or2_1 _25042_ (.A(_09135_),
    .B(_09136_),
    .X(_09137_));
 sky130_fd_sc_hd__a2bb2o_1 _25043_ (.A1_N(_09134_),
    .A2_N(_09137_),
    .B1(_09134_),
    .B2(_09137_),
    .X(_09138_));
 sky130_fd_sc_hd__o21ba_1 _25044_ (.A1(_09010_),
    .A2(_09014_),
    .B1_N(_09013_),
    .X(_09139_));
 sky130_fd_sc_hd__a2bb2o_1 _25045_ (.A1_N(_09138_),
    .A2_N(_09139_),
    .B1(_09138_),
    .B2(_09139_),
    .X(_09140_));
 sky130_fd_sc_hd__a2bb2o_2 _25046_ (.A1_N(_09133_),
    .A2_N(_09140_),
    .B1(_09133_),
    .B2(_09140_),
    .X(_09141_));
 sky130_fd_sc_hd__a21oi_2 _25047_ (.A1(_09024_),
    .A2(_09026_),
    .B1(_09023_),
    .Y(_09142_));
 sky130_fd_sc_hd__o21ba_1 _25048_ (.A1(_09037_),
    .A2(_09040_),
    .B1_N(_09039_),
    .X(_09143_));
 sky130_fd_sc_hd__o22a_1 _25049_ (.A1(_08869_),
    .A2(_06650_),
    .B1(_08870_),
    .B2(_07332_),
    .X(_09144_));
 sky130_fd_sc_hd__and4_2 _25050_ (.A(_08872_),
    .B(_07329_),
    .C(_08873_),
    .D(_07764_),
    .X(_09145_));
 sky130_fd_sc_hd__nor2_2 _25051_ (.A(_09144_),
    .B(_09145_),
    .Y(_09146_));
 sky130_fd_sc_hd__buf_2 _25052_ (.A(_05999_),
    .X(_09147_));
 sky130_fd_sc_hd__nor2_2 _25053_ (.A(_09147_),
    .B(_06892_),
    .Y(_09148_));
 sky130_fd_sc_hd__a2bb2o_1 _25054_ (.A1_N(_09146_),
    .A2_N(_09148_),
    .B1(_09146_),
    .B2(_09148_),
    .X(_09149_));
 sky130_fd_sc_hd__a2bb2o_1 _25055_ (.A1_N(_09143_),
    .A2_N(_09149_),
    .B1(_09143_),
    .B2(_09149_),
    .X(_09150_));
 sky130_fd_sc_hd__a2bb2o_1 _25056_ (.A1_N(_09142_),
    .A2_N(_09150_),
    .B1(_09142_),
    .B2(_09150_),
    .X(_09151_));
 sky130_fd_sc_hd__o22a_1 _25057_ (.A1(_09020_),
    .A2(_09027_),
    .B1(_09019_),
    .B2(_09028_),
    .X(_09152_));
 sky130_fd_sc_hd__a2bb2o_1 _25058_ (.A1_N(_09151_),
    .A2_N(_09152_),
    .B1(_09151_),
    .B2(_09152_),
    .X(_09153_));
 sky130_fd_sc_hd__a2bb2o_1 _25059_ (.A1_N(_09141_),
    .A2_N(_09153_),
    .B1(_09141_),
    .B2(_09153_),
    .X(_09154_));
 sky130_fd_sc_hd__a2bb2o_1 _25060_ (.A1_N(_09128_),
    .A2_N(_09154_),
    .B1(_09128_),
    .B2(_09154_),
    .X(_09155_));
 sky130_fd_sc_hd__a2bb2o_1 _25061_ (.A1_N(_09127_),
    .A2_N(_09155_),
    .B1(_09127_),
    .B2(_09155_),
    .X(_09156_));
 sky130_fd_sc_hd__o22a_1 _25062_ (.A1(_09046_),
    .A2(_09047_),
    .B1(_09041_),
    .B2(_09048_),
    .X(_09157_));
 sky130_fd_sc_hd__o22a_1 _25063_ (.A1(_09053_),
    .A2(_09058_),
    .B1(_09052_),
    .B2(_09059_),
    .X(_09158_));
 sky130_fd_sc_hd__or2_1 _25064_ (.A(_06285_),
    .B(_06641_),
    .X(_09159_));
 sky130_fd_sc_hd__o22a_1 _25065_ (.A1(_08416_),
    .A2(_06437_),
    .B1(_08575_),
    .B2(_08719_),
    .X(_09160_));
 sky130_fd_sc_hd__and4_1 _25066_ (.A(_08577_),
    .B(_07212_),
    .C(_08578_),
    .D(_07485_),
    .X(_09161_));
 sky130_fd_sc_hd__or2_1 _25067_ (.A(_09160_),
    .B(_09161_),
    .X(_09162_));
 sky130_fd_sc_hd__a2bb2o_1 _25068_ (.A1_N(_09159_),
    .A2_N(_09162_),
    .B1(_09159_),
    .B2(_09162_),
    .X(_09163_));
 sky130_fd_sc_hd__or2_1 _25069_ (.A(_08582_),
    .B(_06917_),
    .X(_09164_));
 sky130_fd_sc_hd__o22a_1 _25070_ (.A1(_08743_),
    .A2(_06131_),
    .B1(_08424_),
    .B2(_06218_),
    .X(_09165_));
 sky130_fd_sc_hd__and4_1 _25071_ (.A(_08585_),
    .B(_13570_),
    .C(_08586_),
    .D(_08738_),
    .X(_09166_));
 sky130_fd_sc_hd__or2_1 _25072_ (.A(_09165_),
    .B(_09166_),
    .X(_09167_));
 sky130_fd_sc_hd__a2bb2o_1 _25073_ (.A1_N(_09164_),
    .A2_N(_09167_),
    .B1(_09164_),
    .B2(_09167_),
    .X(_09168_));
 sky130_fd_sc_hd__o21ba_1 _25074_ (.A1(_09042_),
    .A2(_09045_),
    .B1_N(_09044_),
    .X(_09169_));
 sky130_fd_sc_hd__a2bb2o_1 _25075_ (.A1_N(_09168_),
    .A2_N(_09169_),
    .B1(_09168_),
    .B2(_09169_),
    .X(_09170_));
 sky130_fd_sc_hd__a2bb2o_1 _25076_ (.A1_N(_09163_),
    .A2_N(_09170_),
    .B1(_09163_),
    .B2(_09170_),
    .X(_09171_));
 sky130_fd_sc_hd__a2bb2o_1 _25077_ (.A1_N(_09158_),
    .A2_N(_09171_),
    .B1(_09158_),
    .B2(_09171_),
    .X(_09172_));
 sky130_fd_sc_hd__a2bb2o_1 _25078_ (.A1_N(_09157_),
    .A2_N(_09172_),
    .B1(_09157_),
    .B2(_09172_),
    .X(_09173_));
 sky130_fd_sc_hd__o21ba_1 _25079_ (.A1(_09054_),
    .A2(_09057_),
    .B1_N(_09056_),
    .X(_09174_));
 sky130_fd_sc_hd__o21ba_1 _25080_ (.A1(_09061_),
    .A2(_09064_),
    .B1_N(_09063_),
    .X(_09175_));
 sky130_fd_sc_hd__or2_1 _25081_ (.A(_08118_),
    .B(_06130_),
    .X(_09176_));
 sky130_fd_sc_hd__o22a_1 _25082_ (.A1(_08120_),
    .A2(_06484_),
    .B1(_08121_),
    .B2(_05931_),
    .X(_09177_));
 sky130_fd_sc_hd__and4_1 _25083_ (.A(_08603_),
    .B(_08587_),
    .C(_08441_),
    .D(_13579_),
    .X(_09178_));
 sky130_fd_sc_hd__or2_1 _25084_ (.A(_09177_),
    .B(_09178_),
    .X(_09179_));
 sky130_fd_sc_hd__a2bb2o_1 _25085_ (.A1_N(_09176_),
    .A2_N(_09179_),
    .B1(_09176_),
    .B2(_09179_),
    .X(_09180_));
 sky130_fd_sc_hd__a2bb2o_1 _25086_ (.A1_N(_09175_),
    .A2_N(_09180_),
    .B1(_09175_),
    .B2(_09180_),
    .X(_09181_));
 sky130_fd_sc_hd__a2bb2o_1 _25087_ (.A1_N(_09174_),
    .A2_N(_09181_),
    .B1(_09174_),
    .B2(_09181_),
    .X(_09182_));
 sky130_fd_sc_hd__or2_1 _25088_ (.A(_08609_),
    .B(_05818_),
    .X(_09183_));
 sky130_fd_sc_hd__o22a_1 _25089_ (.A1(_08286_),
    .A2(_07255_),
    .B1(_08287_),
    .B2(_08263_),
    .X(_09184_));
 sky130_fd_sc_hd__and4_1 _25090_ (.A(_13073_),
    .B(_07251_),
    .C(_13078_),
    .D(_08265_),
    .X(_09185_));
 sky130_fd_sc_hd__or2_1 _25091_ (.A(_09184_),
    .B(_09185_),
    .X(_09186_));
 sky130_fd_sc_hd__a2bb2o_1 _25092_ (.A1_N(_09183_),
    .A2_N(_09186_),
    .B1(_09183_),
    .B2(_09186_),
    .X(_09187_));
 sky130_fd_sc_hd__buf_1 _25093_ (.A(_07970_),
    .X(_09188_));
 sky130_fd_sc_hd__or2_1 _25094_ (.A(_09188_),
    .B(_08439_),
    .X(_09189_));
 sky130_fd_sc_hd__buf_1 _25095_ (.A(_08294_),
    .X(_09190_));
 sky130_fd_sc_hd__buf_1 _25096_ (.A(_08457_),
    .X(_09191_));
 sky130_fd_sc_hd__and4_1 _25097_ (.A(_09190_),
    .B(_05868_),
    .C(_09191_),
    .D(_13598_),
    .X(_09192_));
 sky130_fd_sc_hd__o22a_1 _25098_ (.A1(_11718_),
    .A2(_07405_),
    .B1(_08132_),
    .B2(_06301_),
    .X(_09193_));
 sky130_fd_sc_hd__or2_1 _25099_ (.A(_09192_),
    .B(_09193_),
    .X(_09194_));
 sky130_fd_sc_hd__a2bb2o_1 _25100_ (.A1_N(_09189_),
    .A2_N(_09194_),
    .B1(_09189_),
    .B2(_09194_),
    .X(_09195_));
 sky130_fd_sc_hd__o21ba_1 _25101_ (.A1(_09066_),
    .A2(_09071_),
    .B1_N(_09068_),
    .X(_09196_));
 sky130_fd_sc_hd__a2bb2o_1 _25102_ (.A1_N(_09195_),
    .A2_N(_09196_),
    .B1(_09195_),
    .B2(_09196_),
    .X(_09197_));
 sky130_fd_sc_hd__a2bb2o_1 _25103_ (.A1_N(_09187_),
    .A2_N(_09197_),
    .B1(_09187_),
    .B2(_09197_),
    .X(_09198_));
 sky130_fd_sc_hd__o22a_1 _25104_ (.A1(_09072_),
    .A2(_09073_),
    .B1(_09065_),
    .B2(_09074_),
    .X(_09199_));
 sky130_fd_sc_hd__a2bb2o_1 _25105_ (.A1_N(_09198_),
    .A2_N(_09199_),
    .B1(_09198_),
    .B2(_09199_),
    .X(_09200_));
 sky130_fd_sc_hd__a2bb2o_1 _25106_ (.A1_N(_09182_),
    .A2_N(_09200_),
    .B1(_09182_),
    .B2(_09200_),
    .X(_09201_));
 sky130_fd_sc_hd__o22a_1 _25107_ (.A1(_09075_),
    .A2(_09076_),
    .B1(_09060_),
    .B2(_09077_),
    .X(_09202_));
 sky130_fd_sc_hd__a2bb2o_1 _25108_ (.A1_N(_09201_),
    .A2_N(_09202_),
    .B1(_09201_),
    .B2(_09202_),
    .X(_09203_));
 sky130_fd_sc_hd__a2bb2o_1 _25109_ (.A1_N(_09173_),
    .A2_N(_09203_),
    .B1(_09173_),
    .B2(_09203_),
    .X(_09204_));
 sky130_fd_sc_hd__o22a_1 _25110_ (.A1(_09078_),
    .A2(_09079_),
    .B1(_09051_),
    .B2(_09080_),
    .X(_09205_));
 sky130_fd_sc_hd__a2bb2o_1 _25111_ (.A1_N(_09204_),
    .A2_N(_09205_),
    .B1(_09204_),
    .B2(_09205_),
    .X(_09206_));
 sky130_fd_sc_hd__a2bb2o_1 _25112_ (.A1_N(_09156_),
    .A2_N(_09206_),
    .B1(_09156_),
    .B2(_09206_),
    .X(_09207_));
 sky130_fd_sc_hd__o22a_1 _25113_ (.A1(_09081_),
    .A2(_09082_),
    .B1(_09034_),
    .B2(_09083_),
    .X(_09208_));
 sky130_fd_sc_hd__a2bb2o_1 _25114_ (.A1_N(_09207_),
    .A2_N(_09208_),
    .B1(_09207_),
    .B2(_09208_),
    .X(_09209_));
 sky130_fd_sc_hd__a2bb2o_1 _25115_ (.A1_N(_09126_),
    .A2_N(_09209_),
    .B1(_09126_),
    .B2(_09209_),
    .X(_09210_));
 sky130_fd_sc_hd__o22a_1 _25116_ (.A1(_09084_),
    .A2(_09085_),
    .B1(_09000_),
    .B2(_09086_),
    .X(_09211_));
 sky130_fd_sc_hd__a2bb2o_1 _25117_ (.A1_N(_09210_),
    .A2_N(_09211_),
    .B1(_09210_),
    .B2(_09211_),
    .X(_09212_));
 sky130_fd_sc_hd__a2bb2o_1 _25118_ (.A1_N(_09100_),
    .A2_N(_09212_),
    .B1(_09100_),
    .B2(_09212_),
    .X(_09213_));
 sky130_fd_sc_hd__o22a_1 _25119_ (.A1(_09087_),
    .A2(_09088_),
    .B1(_08968_),
    .B2(_09089_),
    .X(_09214_));
 sky130_fd_sc_hd__a2bb2o_1 _25120_ (.A1_N(_09213_),
    .A2_N(_09214_),
    .B1(_09213_),
    .B2(_09214_),
    .X(_09215_));
 sky130_fd_sc_hd__a2bb2o_1 _25121_ (.A1_N(_08967_),
    .A2_N(_09215_),
    .B1(_08967_),
    .B2(_09215_),
    .X(_09216_));
 sky130_fd_sc_hd__o22a_1 _25122_ (.A1(_09090_),
    .A2(_09091_),
    .B1(_08808_),
    .B2(_09092_),
    .X(_09217_));
 sky130_fd_sc_hd__or2_1 _25123_ (.A(_09216_),
    .B(_09217_),
    .X(_09218_));
 sky130_fd_sc_hd__a21bo_2 _25124_ (.A1(_09216_),
    .A2(_09217_),
    .B1_N(_09218_),
    .X(_09219_));
 sky130_fd_sc_hd__a22o_1 _25125_ (.A1(_08962_),
    .A2(_09093_),
    .B1(_08952_),
    .B2(_09094_),
    .X(_09220_));
 sky130_fd_sc_hd__o31a_2 _25126_ (.A1(_08954_),
    .A2(_09095_),
    .A3(_08960_),
    .B1(_09220_),
    .X(_09221_));
 sky130_fd_sc_hd__a2bb2oi_4 _25127_ (.A1_N(_09219_),
    .A2_N(_09221_),
    .B1(_09219_),
    .B2(_09221_),
    .Y(_02657_));
 sky130_fd_sc_hd__o22a_1 _25128_ (.A1(_09213_),
    .A2(_09214_),
    .B1(_08967_),
    .B2(_09215_),
    .X(_09222_));
 sky130_fd_sc_hd__o22a_1 _25129_ (.A1(_09102_),
    .A2(_09124_),
    .B1(_09101_),
    .B2(_09125_),
    .X(_09223_));
 sky130_fd_sc_hd__or3_4 _25130_ (.A(_05143_),
    .B(_08973_),
    .C(_08663_),
    .X(_09224_));
 sky130_fd_sc_hd__o21a_1 _25131_ (.A1(_08965_),
    .A2(_09105_),
    .B1(_09224_),
    .X(_09225_));
 sky130_fd_sc_hd__or2_1 _25132_ (.A(_09223_),
    .B(_09225_),
    .X(_09226_));
 sky130_fd_sc_hd__a21bo_1 _25133_ (.A1(_09223_),
    .A2(_09225_),
    .B1_N(_09226_),
    .X(_09227_));
 sky130_fd_sc_hd__o22a_1 _25134_ (.A1(_09121_),
    .A2(_09122_),
    .B1(_09106_),
    .B2(_09123_),
    .X(_09228_));
 sky130_fd_sc_hd__o22a_1 _25135_ (.A1(_09128_),
    .A2(_09154_),
    .B1(_09127_),
    .B2(_09155_),
    .X(_09229_));
 sky130_fd_sc_hd__a21bo_1 _25136_ (.A1(_08664_),
    .A2(_09104_),
    .B1_N(_09224_),
    .X(_09230_));
 sky130_fd_sc_hd__a2bb2o_1 _25137_ (.A1_N(_08812_),
    .A2_N(_09230_),
    .B1(_08812_),
    .B2(_09230_),
    .X(_09231_));
 sky130_fd_sc_hd__buf_1 _25138_ (.A(_09231_),
    .X(_09232_));
 sky130_fd_sc_hd__buf_1 _25139_ (.A(_09232_),
    .X(_09233_));
 sky130_fd_sc_hd__o22a_1 _25140_ (.A1(_09110_),
    .A2(_09117_),
    .B1(_09109_),
    .B2(_09118_),
    .X(_09234_));
 sky130_fd_sc_hd__o22a_1 _25141_ (.A1(_09138_),
    .A2(_09139_),
    .B1(_09133_),
    .B2(_09140_),
    .X(_09235_));
 sky130_fd_sc_hd__buf_1 _25142_ (.A(_09116_),
    .X(_09236_));
 sky130_fd_sc_hd__o21ba_1 _25143_ (.A1(_09113_),
    .A2(_09236_),
    .B1_N(_09112_),
    .X(_09237_));
 sky130_fd_sc_hd__a21oi_2 _25144_ (.A1(_09131_),
    .A2(_09132_),
    .B1(_09130_),
    .Y(_09238_));
 sky130_fd_sc_hd__clkbuf_2 _25145_ (.A(_08497_),
    .X(_09239_));
 sky130_fd_sc_hd__nor2_1 _25146_ (.A(_08683_),
    .B(_09239_),
    .Y(_09240_));
 sky130_fd_sc_hd__clkbuf_1 _25147_ (.A(_11700_),
    .X(_09241_));
 sky130_fd_sc_hd__or2_2 _25148_ (.A(_09241_),
    .B(_05454_),
    .X(_09242_));
 sky130_vsdinv _25149_ (.A(_09242_),
    .Y(_09243_));
 sky130_fd_sc_hd__a2bb2o_1 _25150_ (.A1_N(_09240_),
    .A2_N(_09243_),
    .B1(_09240_),
    .B2(_09243_),
    .X(_09244_));
 sky130_fd_sc_hd__a2bb2o_1 _25151_ (.A1_N(_09236_),
    .A2_N(_09244_),
    .B1(_09236_),
    .B2(_09244_),
    .X(_09245_));
 sky130_fd_sc_hd__a2bb2o_1 _25152_ (.A1_N(_09238_),
    .A2_N(_09245_),
    .B1(_09238_),
    .B2(_09245_),
    .X(_09246_));
 sky130_fd_sc_hd__a2bb2o_1 _25153_ (.A1_N(_09237_),
    .A2_N(_09246_),
    .B1(_09237_),
    .B2(_09246_),
    .X(_09247_));
 sky130_fd_sc_hd__a2bb2o_1 _25154_ (.A1_N(_09235_),
    .A2_N(_09247_),
    .B1(_09235_),
    .B2(_09247_),
    .X(_09248_));
 sky130_fd_sc_hd__a2bb2o_1 _25155_ (.A1_N(_09234_),
    .A2_N(_09248_),
    .B1(_09234_),
    .B2(_09248_),
    .X(_09249_));
 sky130_fd_sc_hd__o22a_1 _25156_ (.A1(_09108_),
    .A2(_09119_),
    .B1(_09107_),
    .B2(_09120_),
    .X(_09250_));
 sky130_fd_sc_hd__a2bb2o_1 _25157_ (.A1_N(_09249_),
    .A2_N(_09250_),
    .B1(_09249_),
    .B2(_09250_),
    .X(_09251_));
 sky130_fd_sc_hd__buf_1 _25158_ (.A(_09232_),
    .X(_09252_));
 sky130_fd_sc_hd__a2bb2o_2 _25159_ (.A1_N(_09233_),
    .A2_N(_09251_),
    .B1(_09252_),
    .B2(_09251_),
    .X(_09253_));
 sky130_fd_sc_hd__a2bb2o_1 _25160_ (.A1_N(_09229_),
    .A2_N(_09253_),
    .B1(_09229_),
    .B2(_09253_),
    .X(_09254_));
 sky130_fd_sc_hd__a2bb2o_1 _25161_ (.A1_N(_09228_),
    .A2_N(_09254_),
    .B1(_09228_),
    .B2(_09254_),
    .X(_09255_));
 sky130_fd_sc_hd__o22a_1 _25162_ (.A1(_09151_),
    .A2(_09152_),
    .B1(_09141_),
    .B2(_09153_),
    .X(_09256_));
 sky130_fd_sc_hd__o22a_1 _25163_ (.A1(_09158_),
    .A2(_09171_),
    .B1(_09157_),
    .B2(_09172_),
    .X(_09257_));
 sky130_fd_sc_hd__clkbuf_2 _25164_ (.A(_07748_),
    .X(_09258_));
 sky130_fd_sc_hd__o22a_1 _25165_ (.A1(_09003_),
    .A2(_07870_),
    .B1(_05589_),
    .B2(_09258_),
    .X(_09259_));
 sky130_fd_sc_hd__and4_2 _25166_ (.A(_13138_),
    .B(_13520_),
    .C(_13144_),
    .D(_08023_),
    .X(_09260_));
 sky130_fd_sc_hd__nor2_2 _25167_ (.A(_09259_),
    .B(_09260_),
    .Y(_09261_));
 sky130_fd_sc_hd__nor2_2 _25168_ (.A(_05538_),
    .B(_08020_),
    .Y(_09262_));
 sky130_fd_sc_hd__a2bb2o_1 _25169_ (.A1_N(_09261_),
    .A2_N(_09262_),
    .B1(_09261_),
    .B2(_09262_),
    .X(_09263_));
 sky130_fd_sc_hd__or2_1 _25170_ (.A(_05791_),
    .B(_07463_),
    .X(_09264_));
 sky130_fd_sc_hd__o22a_1 _25171_ (.A1(_06830_),
    .A2(_07195_),
    .B1(_07238_),
    .B2(_07324_),
    .X(_09265_));
 sky130_fd_sc_hd__and4_1 _25172_ (.A(_07115_),
    .B(_07741_),
    .C(_07116_),
    .D(_07448_),
    .X(_09266_));
 sky130_fd_sc_hd__or2_1 _25173_ (.A(_09265_),
    .B(_09266_),
    .X(_09267_));
 sky130_fd_sc_hd__a2bb2o_1 _25174_ (.A1_N(_09264_),
    .A2_N(_09267_),
    .B1(_09264_),
    .B2(_09267_),
    .X(_09268_));
 sky130_fd_sc_hd__o21ba_1 _25175_ (.A1(_09134_),
    .A2(_09137_),
    .B1_N(_09136_),
    .X(_09269_));
 sky130_fd_sc_hd__a2bb2o_1 _25176_ (.A1_N(_09268_),
    .A2_N(_09269_),
    .B1(_09268_),
    .B2(_09269_),
    .X(_09270_));
 sky130_fd_sc_hd__a2bb2o_2 _25177_ (.A1_N(_09263_),
    .A2_N(_09270_),
    .B1(_09263_),
    .B2(_09270_),
    .X(_09271_));
 sky130_fd_sc_hd__a21oi_2 _25178_ (.A1(_09146_),
    .A2(_09148_),
    .B1(_09145_),
    .Y(_09272_));
 sky130_fd_sc_hd__o21ba_1 _25179_ (.A1(_09159_),
    .A2(_09162_),
    .B1_N(_09161_),
    .X(_09273_));
 sky130_fd_sc_hd__buf_1 _25180_ (.A(_06093_),
    .X(_09274_));
 sky130_fd_sc_hd__o22a_1 _25181_ (.A1(_08869_),
    .A2(_06762_),
    .B1(_09274_),
    .B2(_07468_),
    .X(_09275_));
 sky130_fd_sc_hd__and4_2 _25182_ (.A(_08872_),
    .B(_07764_),
    .C(_08873_),
    .D(_08053_),
    .X(_09276_));
 sky130_fd_sc_hd__nor2_2 _25183_ (.A(_09275_),
    .B(_09276_),
    .Y(_09277_));
 sky130_fd_sc_hd__nor2_2 _25184_ (.A(_09147_),
    .B(_07034_),
    .Y(_09278_));
 sky130_fd_sc_hd__a2bb2o_1 _25185_ (.A1_N(_09277_),
    .A2_N(_09278_),
    .B1(_09277_),
    .B2(_09278_),
    .X(_09279_));
 sky130_fd_sc_hd__a2bb2o_1 _25186_ (.A1_N(_09273_),
    .A2_N(_09279_),
    .B1(_09273_),
    .B2(_09279_),
    .X(_09280_));
 sky130_fd_sc_hd__a2bb2o_1 _25187_ (.A1_N(_09272_),
    .A2_N(_09280_),
    .B1(_09272_),
    .B2(_09280_),
    .X(_09281_));
 sky130_fd_sc_hd__o22a_1 _25188_ (.A1(_09143_),
    .A2(_09149_),
    .B1(_09142_),
    .B2(_09150_),
    .X(_09282_));
 sky130_fd_sc_hd__a2bb2o_1 _25189_ (.A1_N(_09281_),
    .A2_N(_09282_),
    .B1(_09281_),
    .B2(_09282_),
    .X(_09283_));
 sky130_fd_sc_hd__a2bb2o_1 _25190_ (.A1_N(_09271_),
    .A2_N(_09283_),
    .B1(_09271_),
    .B2(_09283_),
    .X(_09284_));
 sky130_fd_sc_hd__a2bb2o_1 _25191_ (.A1_N(_09257_),
    .A2_N(_09284_),
    .B1(_09257_),
    .B2(_09284_),
    .X(_09285_));
 sky130_fd_sc_hd__a2bb2o_1 _25192_ (.A1_N(_09256_),
    .A2_N(_09285_),
    .B1(_09256_),
    .B2(_09285_),
    .X(_09286_));
 sky130_fd_sc_hd__o22a_1 _25193_ (.A1(_09168_),
    .A2(_09169_),
    .B1(_09163_),
    .B2(_09170_),
    .X(_09287_));
 sky130_fd_sc_hd__o22a_1 _25194_ (.A1(_09175_),
    .A2(_09180_),
    .B1(_09174_),
    .B2(_09181_),
    .X(_09288_));
 sky130_fd_sc_hd__or2_1 _25195_ (.A(_08253_),
    .B(_06878_),
    .X(_09289_));
 sky130_fd_sc_hd__o22a_1 _25196_ (.A1(_08416_),
    .A2(_07348_),
    .B1(_08575_),
    .B2(_08388_),
    .X(_09290_));
 sky130_fd_sc_hd__and4_1 _25197_ (.A(_08256_),
    .B(_07485_),
    .C(_08578_),
    .D(_07187_),
    .X(_09291_));
 sky130_fd_sc_hd__or2_1 _25198_ (.A(_09290_),
    .B(_09291_),
    .X(_09292_));
 sky130_fd_sc_hd__a2bb2o_2 _25199_ (.A1_N(_09289_),
    .A2_N(_09292_),
    .B1(_09289_),
    .B2(_09292_),
    .X(_09293_));
 sky130_fd_sc_hd__or2_1 _25200_ (.A(_08582_),
    .B(_08887_),
    .X(_09294_));
 sky130_fd_sc_hd__o22a_1 _25201_ (.A1(_08743_),
    .A2(_06921_),
    .B1(_08424_),
    .B2(_06329_),
    .X(_09295_));
 sky130_fd_sc_hd__and4_1 _25202_ (.A(_08585_),
    .B(_08738_),
    .C(_08586_),
    .D(_07059_),
    .X(_09296_));
 sky130_fd_sc_hd__or2_1 _25203_ (.A(_09295_),
    .B(_09296_),
    .X(_09297_));
 sky130_fd_sc_hd__a2bb2o_1 _25204_ (.A1_N(_09294_),
    .A2_N(_09297_),
    .B1(_09294_),
    .B2(_09297_),
    .X(_09298_));
 sky130_fd_sc_hd__o21ba_1 _25205_ (.A1(_09164_),
    .A2(_09167_),
    .B1_N(_09166_),
    .X(_09299_));
 sky130_fd_sc_hd__a2bb2o_1 _25206_ (.A1_N(_09298_),
    .A2_N(_09299_),
    .B1(_09298_),
    .B2(_09299_),
    .X(_09300_));
 sky130_fd_sc_hd__a2bb2o_1 _25207_ (.A1_N(_09293_),
    .A2_N(_09300_),
    .B1(_09293_),
    .B2(_09300_),
    .X(_09301_));
 sky130_fd_sc_hd__a2bb2o_1 _25208_ (.A1_N(_09288_),
    .A2_N(_09301_),
    .B1(_09288_),
    .B2(_09301_),
    .X(_09302_));
 sky130_fd_sc_hd__a2bb2o_1 _25209_ (.A1_N(_09287_),
    .A2_N(_09302_),
    .B1(_09287_),
    .B2(_09302_),
    .X(_09303_));
 sky130_fd_sc_hd__o21ba_1 _25210_ (.A1(_09176_),
    .A2(_09179_),
    .B1_N(_09178_),
    .X(_09304_));
 sky130_fd_sc_hd__o21ba_1 _25211_ (.A1(_09183_),
    .A2(_09186_),
    .B1_N(_09185_),
    .X(_09305_));
 sky130_fd_sc_hd__buf_1 _25212_ (.A(_08599_),
    .X(_09306_));
 sky130_fd_sc_hd__buf_1 _25213_ (.A(_07267_),
    .X(_09307_));
 sky130_fd_sc_hd__o22a_1 _25214_ (.A1(_09306_),
    .A2(_05837_),
    .B1(_09307_),
    .B2(_05944_),
    .X(_09308_));
 sky130_fd_sc_hd__buf_1 _25215_ (.A(_08124_),
    .X(_09309_));
 sky130_fd_sc_hd__and4_2 _25216_ (.A(_08761_),
    .B(_08747_),
    .C(_09309_),
    .D(_06460_),
    .X(_09310_));
 sky130_fd_sc_hd__nor2_2 _25217_ (.A(_09308_),
    .B(_09310_),
    .Y(_09311_));
 sky130_fd_sc_hd__nor2_2 _25218_ (.A(_08758_),
    .B(_06334_),
    .Y(_09312_));
 sky130_fd_sc_hd__a2bb2o_1 _25219_ (.A1_N(_09311_),
    .A2_N(_09312_),
    .B1(_09311_),
    .B2(_09312_),
    .X(_09313_));
 sky130_fd_sc_hd__a2bb2o_1 _25220_ (.A1_N(_09305_),
    .A2_N(_09313_),
    .B1(_09305_),
    .B2(_09313_),
    .X(_09314_));
 sky130_fd_sc_hd__a2bb2o_1 _25221_ (.A1_N(_09304_),
    .A2_N(_09314_),
    .B1(_09304_),
    .B2(_09314_),
    .X(_09315_));
 sky130_fd_sc_hd__or2_1 _25222_ (.A(_07531_),
    .B(_05821_),
    .X(_09316_));
 sky130_fd_sc_hd__o22a_1 _25223_ (.A1(_08448_),
    .A2(_08263_),
    .B1(_08449_),
    .B2(_08425_),
    .X(_09317_));
 sky130_fd_sc_hd__and4_1 _25224_ (.A(_08613_),
    .B(_08265_),
    .C(_08614_),
    .D(_08427_),
    .X(_09318_));
 sky130_fd_sc_hd__or2_1 _25225_ (.A(_09317_),
    .B(_09318_),
    .X(_09319_));
 sky130_fd_sc_hd__a2bb2o_1 _25226_ (.A1_N(_09316_),
    .A2_N(_09319_),
    .B1(_09316_),
    .B2(_09319_),
    .X(_09320_));
 sky130_fd_sc_hd__or2_1 _25227_ (.A(_09188_),
    .B(_06298_),
    .X(_09321_));
 sky130_fd_sc_hd__and4_1 _25228_ (.A(_09190_),
    .B(_05861_),
    .C(_09191_),
    .D(_13594_),
    .X(_09322_));
 sky130_fd_sc_hd__o22a_1 _25229_ (.A1(_08777_),
    .A2(_07820_),
    .B1(_08778_),
    .B2(_06831_),
    .X(_09323_));
 sky130_fd_sc_hd__or2_1 _25230_ (.A(_09322_),
    .B(_09323_),
    .X(_09324_));
 sky130_fd_sc_hd__a2bb2o_1 _25231_ (.A1_N(_09321_),
    .A2_N(_09324_),
    .B1(_09321_),
    .B2(_09324_),
    .X(_09325_));
 sky130_fd_sc_hd__o21ba_1 _25232_ (.A1(_09189_),
    .A2(_09194_),
    .B1_N(_09192_),
    .X(_09326_));
 sky130_fd_sc_hd__a2bb2o_1 _25233_ (.A1_N(_09325_),
    .A2_N(_09326_),
    .B1(_09325_),
    .B2(_09326_),
    .X(_09327_));
 sky130_fd_sc_hd__a2bb2o_1 _25234_ (.A1_N(_09320_),
    .A2_N(_09327_),
    .B1(_09320_),
    .B2(_09327_),
    .X(_09328_));
 sky130_fd_sc_hd__o22a_1 _25235_ (.A1(_09195_),
    .A2(_09196_),
    .B1(_09187_),
    .B2(_09197_),
    .X(_09329_));
 sky130_fd_sc_hd__a2bb2o_1 _25236_ (.A1_N(_09328_),
    .A2_N(_09329_),
    .B1(_09328_),
    .B2(_09329_),
    .X(_09330_));
 sky130_fd_sc_hd__a2bb2o_1 _25237_ (.A1_N(_09315_),
    .A2_N(_09330_),
    .B1(_09315_),
    .B2(_09330_),
    .X(_09331_));
 sky130_fd_sc_hd__o22a_1 _25238_ (.A1(_09198_),
    .A2(_09199_),
    .B1(_09182_),
    .B2(_09200_),
    .X(_09332_));
 sky130_fd_sc_hd__a2bb2o_1 _25239_ (.A1_N(_09331_),
    .A2_N(_09332_),
    .B1(_09331_),
    .B2(_09332_),
    .X(_09333_));
 sky130_fd_sc_hd__a2bb2o_1 _25240_ (.A1_N(_09303_),
    .A2_N(_09333_),
    .B1(_09303_),
    .B2(_09333_),
    .X(_09334_));
 sky130_fd_sc_hd__o22a_1 _25241_ (.A1(_09201_),
    .A2(_09202_),
    .B1(_09173_),
    .B2(_09203_),
    .X(_09335_));
 sky130_fd_sc_hd__a2bb2o_1 _25242_ (.A1_N(_09334_),
    .A2_N(_09335_),
    .B1(_09334_),
    .B2(_09335_),
    .X(_09336_));
 sky130_fd_sc_hd__a2bb2o_1 _25243_ (.A1_N(_09286_),
    .A2_N(_09336_),
    .B1(_09286_),
    .B2(_09336_),
    .X(_09337_));
 sky130_fd_sc_hd__o22a_1 _25244_ (.A1(_09204_),
    .A2(_09205_),
    .B1(_09156_),
    .B2(_09206_),
    .X(_09338_));
 sky130_fd_sc_hd__a2bb2o_1 _25245_ (.A1_N(_09337_),
    .A2_N(_09338_),
    .B1(_09337_),
    .B2(_09338_),
    .X(_09339_));
 sky130_fd_sc_hd__a2bb2o_1 _25246_ (.A1_N(_09255_),
    .A2_N(_09339_),
    .B1(_09255_),
    .B2(_09339_),
    .X(_09340_));
 sky130_fd_sc_hd__o22a_1 _25247_ (.A1(_09207_),
    .A2(_09208_),
    .B1(_09126_),
    .B2(_09209_),
    .X(_09341_));
 sky130_fd_sc_hd__a2bb2o_1 _25248_ (.A1_N(_09340_),
    .A2_N(_09341_),
    .B1(_09340_),
    .B2(_09341_),
    .X(_09342_));
 sky130_fd_sc_hd__a2bb2o_1 _25249_ (.A1_N(_09227_),
    .A2_N(_09342_),
    .B1(_09227_),
    .B2(_09342_),
    .X(_09343_));
 sky130_fd_sc_hd__o22a_1 _25250_ (.A1(_09210_),
    .A2(_09211_),
    .B1(_09100_),
    .B2(_09212_),
    .X(_09344_));
 sky130_fd_sc_hd__a2bb2o_1 _25251_ (.A1_N(_09343_),
    .A2_N(_09344_),
    .B1(_09343_),
    .B2(_09344_),
    .X(_09345_));
 sky130_fd_sc_hd__a2bb2o_2 _25252_ (.A1_N(_09099_),
    .A2_N(_09345_),
    .B1(_09099_),
    .B2(_09345_),
    .X(_09346_));
 sky130_fd_sc_hd__a2bb2o_1 _25253_ (.A1_N(_09222_),
    .A2_N(_09346_),
    .B1(_09222_),
    .B2(_09346_),
    .X(_09347_));
 sky130_fd_sc_hd__o21ai_1 _25254_ (.A1(_09219_),
    .A2(_09221_),
    .B1(_09218_),
    .Y(_09348_));
 sky130_fd_sc_hd__a2bb2o_1 _25255_ (.A1_N(_09347_),
    .A2_N(_09348_),
    .B1(_09347_),
    .B2(_09348_),
    .X(_02658_));
 sky130_fd_sc_hd__o22a_1 _25256_ (.A1(_09229_),
    .A2(_09253_),
    .B1(_09228_),
    .B2(_09254_),
    .X(_09349_));
 sky130_fd_sc_hd__o21a_1 _25257_ (.A1(_08965_),
    .A2(_09230_),
    .B1(_09224_),
    .X(_09350_));
 sky130_fd_sc_hd__clkbuf_2 _25258_ (.A(_09350_),
    .X(_09351_));
 sky130_fd_sc_hd__buf_2 _25259_ (.A(_09351_),
    .X(_09352_));
 sky130_fd_sc_hd__clkbuf_2 _25260_ (.A(_09350_),
    .X(_09353_));
 sky130_fd_sc_hd__or2_1 _25261_ (.A(_09349_),
    .B(_09353_),
    .X(_09354_));
 sky130_fd_sc_hd__a21bo_1 _25262_ (.A1(_09349_),
    .A2(_09352_),
    .B1_N(_09354_),
    .X(_09355_));
 sky130_fd_sc_hd__buf_1 _25263_ (.A(_09231_),
    .X(_09356_));
 sky130_fd_sc_hd__buf_1 _25264_ (.A(_09356_),
    .X(_09357_));
 sky130_fd_sc_hd__o22a_1 _25265_ (.A1(_09249_),
    .A2(_09250_),
    .B1(_09357_),
    .B2(_09251_),
    .X(_09358_));
 sky130_fd_sc_hd__o22a_1 _25266_ (.A1(_09257_),
    .A2(_09284_),
    .B1(_09256_),
    .B2(_09285_),
    .X(_09359_));
 sky130_fd_sc_hd__o22a_1 _25267_ (.A1(_09238_),
    .A2(_09245_),
    .B1(_09237_),
    .B2(_09246_),
    .X(_09360_));
 sky130_fd_sc_hd__o22a_1 _25268_ (.A1(_09268_),
    .A2(_09269_),
    .B1(_09263_),
    .B2(_09270_),
    .X(_09361_));
 sky130_fd_sc_hd__o32a_2 _25269_ (.A1(_08683_),
    .A2(_08499_),
    .A3(_09242_),
    .B1(_09236_),
    .B2(_09244_),
    .X(_09362_));
 sky130_fd_sc_hd__a21oi_4 _25270_ (.A1(_09261_),
    .A2(_09262_),
    .B1(_09260_),
    .Y(_09363_));
 sky130_fd_sc_hd__or2_1 _25271_ (.A(_09241_),
    .B(_05682_),
    .X(_09364_));
 sky130_fd_sc_hd__a32o_1 _25272_ (.A1(_08814_),
    .A2(_13146_),
    .A3(_09243_),
    .B1(_09242_),
    .B2(_09364_),
    .X(_09365_));
 sky130_fd_sc_hd__a2bb2o_2 _25273_ (.A1_N(_09116_),
    .A2_N(_09365_),
    .B1(_09115_),
    .B2(_09365_),
    .X(_09366_));
 sky130_fd_sc_hd__buf_1 _25274_ (.A(_09366_),
    .X(_09367_));
 sky130_fd_sc_hd__buf_1 _25275_ (.A(_09367_),
    .X(_09368_));
 sky130_fd_sc_hd__a2bb2o_1 _25276_ (.A1_N(_09363_),
    .A2_N(_09368_),
    .B1(_09363_),
    .B2(_09368_),
    .X(_09369_));
 sky130_fd_sc_hd__a2bb2o_1 _25277_ (.A1_N(_09362_),
    .A2_N(_09369_),
    .B1(_09362_),
    .B2(_09369_),
    .X(_09370_));
 sky130_fd_sc_hd__a2bb2o_1 _25278_ (.A1_N(_09361_),
    .A2_N(_09370_),
    .B1(_09361_),
    .B2(_09370_),
    .X(_09371_));
 sky130_fd_sc_hd__a2bb2o_1 _25279_ (.A1_N(_09360_),
    .A2_N(_09371_),
    .B1(_09360_),
    .B2(_09371_),
    .X(_09372_));
 sky130_fd_sc_hd__o22a_1 _25280_ (.A1(_09235_),
    .A2(_09247_),
    .B1(_09234_),
    .B2(_09248_),
    .X(_09373_));
 sky130_fd_sc_hd__o2bb2ai_1 _25281_ (.A1_N(_09372_),
    .A2_N(_09373_),
    .B1(_09372_),
    .B2(_09373_),
    .Y(_09374_));
 sky130_fd_sc_hd__buf_1 _25282_ (.A(_09231_),
    .X(_09375_));
 sky130_fd_sc_hd__a2bb2o_1 _25283_ (.A1_N(_09252_),
    .A2_N(_09374_),
    .B1(_09375_),
    .B2(_09374_),
    .X(_09376_));
 sky130_fd_sc_hd__a2bb2o_1 _25284_ (.A1_N(_09359_),
    .A2_N(_09376_),
    .B1(_09359_),
    .B2(_09376_),
    .X(_09377_));
 sky130_fd_sc_hd__a2bb2o_2 _25285_ (.A1_N(_09358_),
    .A2_N(_09377_),
    .B1(_09358_),
    .B2(_09377_),
    .X(_09378_));
 sky130_fd_sc_hd__o22a_1 _25286_ (.A1(_09281_),
    .A2(_09282_),
    .B1(_09271_),
    .B2(_09283_),
    .X(_09379_));
 sky130_fd_sc_hd__o22a_1 _25287_ (.A1(_09288_),
    .A2(_09301_),
    .B1(_09287_),
    .B2(_09302_),
    .X(_09380_));
 sky130_fd_sc_hd__o22a_1 _25288_ (.A1(_08537_),
    .A2(_07748_),
    .B1(_08538_),
    .B2(_07890_),
    .X(_09381_));
 sky130_fd_sc_hd__and4_2 _25289_ (.A(_13137_),
    .B(_13515_),
    .C(_13143_),
    .D(_13509_),
    .X(_09382_));
 sky130_fd_sc_hd__nor2_2 _25290_ (.A(_09381_),
    .B(_09382_),
    .Y(_09383_));
 sky130_fd_sc_hd__nor2_2 _25291_ (.A(_08535_),
    .B(_09239_),
    .Y(_09384_));
 sky130_fd_sc_hd__a2bb2o_1 _25292_ (.A1_N(_09383_),
    .A2_N(_09384_),
    .B1(_09383_),
    .B2(_09384_),
    .X(_09385_));
 sky130_fd_sc_hd__o22a_1 _25293_ (.A1(_08223_),
    .A2(_07325_),
    .B1(_08708_),
    .B2(_07732_),
    .X(_09386_));
 sky130_fd_sc_hd__and4_1 _25294_ (.A(_08390_),
    .B(_07448_),
    .C(_08391_),
    .D(_13523_),
    .X(_09387_));
 sky130_fd_sc_hd__nor2_2 _25295_ (.A(_09386_),
    .B(_09387_),
    .Y(_09388_));
 sky130_fd_sc_hd__nor2_2 _25296_ (.A(_08386_),
    .B(_08180_),
    .Y(_09389_));
 sky130_fd_sc_hd__a2bb2o_1 _25297_ (.A1_N(_09388_),
    .A2_N(_09389_),
    .B1(_09388_),
    .B2(_09389_),
    .X(_09390_));
 sky130_fd_sc_hd__o21ba_1 _25298_ (.A1(_09264_),
    .A2(_09267_),
    .B1_N(_09266_),
    .X(_09391_));
 sky130_fd_sc_hd__a2bb2o_1 _25299_ (.A1_N(_09390_),
    .A2_N(_09391_),
    .B1(_09390_),
    .B2(_09391_),
    .X(_09392_));
 sky130_fd_sc_hd__a2bb2o_2 _25300_ (.A1_N(_09385_),
    .A2_N(_09392_),
    .B1(_09385_),
    .B2(_09392_),
    .X(_09393_));
 sky130_fd_sc_hd__a21oi_2 _25301_ (.A1(_09277_),
    .A2(_09278_),
    .B1(_09276_),
    .Y(_09394_));
 sky130_fd_sc_hd__o21ba_1 _25302_ (.A1(_09289_),
    .A2(_09292_),
    .B1_N(_09291_),
    .X(_09395_));
 sky130_fd_sc_hd__clkbuf_2 _25303_ (.A(_07128_),
    .X(_09396_));
 sky130_fd_sc_hd__o22a_1 _25304_ (.A1(_09396_),
    .A2(_06891_),
    .B1(_09274_),
    .B2(_07744_),
    .X(_09397_));
 sky130_fd_sc_hd__buf_1 _25305_ (.A(_07798_),
    .X(_09398_));
 sky130_fd_sc_hd__buf_1 _25306_ (.A(_07799_),
    .X(_09399_));
 sky130_fd_sc_hd__and4_2 _25307_ (.A(_09398_),
    .B(_08053_),
    .C(_09399_),
    .D(_07740_),
    .X(_09400_));
 sky130_fd_sc_hd__nor2_2 _25308_ (.A(_09397_),
    .B(_09400_),
    .Y(_09401_));
 sky130_fd_sc_hd__buf_2 _25309_ (.A(_05999_),
    .X(_09402_));
 sky130_fd_sc_hd__nor2_2 _25310_ (.A(_09402_),
    .B(_07453_),
    .Y(_09403_));
 sky130_fd_sc_hd__a2bb2o_1 _25311_ (.A1_N(_09401_),
    .A2_N(_09403_),
    .B1(_09401_),
    .B2(_09403_),
    .X(_09404_));
 sky130_fd_sc_hd__a2bb2o_1 _25312_ (.A1_N(_09395_),
    .A2_N(_09404_),
    .B1(_09395_),
    .B2(_09404_),
    .X(_09405_));
 sky130_fd_sc_hd__a2bb2o_1 _25313_ (.A1_N(_09394_),
    .A2_N(_09405_),
    .B1(_09394_),
    .B2(_09405_),
    .X(_09406_));
 sky130_fd_sc_hd__o22a_1 _25314_ (.A1(_09273_),
    .A2(_09279_),
    .B1(_09272_),
    .B2(_09280_),
    .X(_09407_));
 sky130_fd_sc_hd__a2bb2o_1 _25315_ (.A1_N(_09406_),
    .A2_N(_09407_),
    .B1(_09406_),
    .B2(_09407_),
    .X(_09408_));
 sky130_fd_sc_hd__a2bb2o_1 _25316_ (.A1_N(_09393_),
    .A2_N(_09408_),
    .B1(_09393_),
    .B2(_09408_),
    .X(_09409_));
 sky130_fd_sc_hd__a2bb2o_1 _25317_ (.A1_N(_09380_),
    .A2_N(_09409_),
    .B1(_09380_),
    .B2(_09409_),
    .X(_09410_));
 sky130_fd_sc_hd__a2bb2o_1 _25318_ (.A1_N(_09379_),
    .A2_N(_09410_),
    .B1(_09379_),
    .B2(_09410_),
    .X(_09411_));
 sky130_fd_sc_hd__o22a_1 _25319_ (.A1(_09298_),
    .A2(_09299_),
    .B1(_09293_),
    .B2(_09300_),
    .X(_09412_));
 sky130_fd_sc_hd__o22a_1 _25320_ (.A1(_09305_),
    .A2(_09313_),
    .B1(_09304_),
    .B2(_09314_),
    .X(_09413_));
 sky130_fd_sc_hd__buf_1 _25321_ (.A(_06390_),
    .X(_09414_));
 sky130_fd_sc_hd__o22a_1 _25322_ (.A1(_08889_),
    .A2(_07037_),
    .B1(_09414_),
    .B2(_07482_),
    .X(_09415_));
 sky130_fd_sc_hd__clkbuf_2 _25323_ (.A(_08102_),
    .X(_09416_));
 sky130_fd_sc_hd__and4_2 _25324_ (.A(_13106_),
    .B(_13553_),
    .C(_09416_),
    .D(_13550_),
    .X(_09417_));
 sky130_fd_sc_hd__nor2_2 _25325_ (.A(_09415_),
    .B(_09417_),
    .Y(_09418_));
 sky130_fd_sc_hd__clkbuf_2 _25326_ (.A(_08253_),
    .X(_09419_));
 sky130_fd_sc_hd__nor2_2 _25327_ (.A(_09419_),
    .B(_09025_),
    .Y(_09420_));
 sky130_fd_sc_hd__a2bb2o_1 _25328_ (.A1_N(_09418_),
    .A2_N(_09420_),
    .B1(_09418_),
    .B2(_09420_),
    .X(_09421_));
 sky130_fd_sc_hd__buf_1 _25329_ (.A(_06801_),
    .X(_09422_));
 sky130_fd_sc_hd__buf_1 _25330_ (.A(_06765_),
    .X(_09423_));
 sky130_fd_sc_hd__o22a_1 _25331_ (.A1(_08897_),
    .A2(_06434_),
    .B1(_09422_),
    .B2(_09423_),
    .X(_09424_));
 sky130_fd_sc_hd__and4_2 _25332_ (.A(_08745_),
    .B(_06654_),
    .C(_08746_),
    .D(_06769_),
    .X(_09425_));
 sky130_fd_sc_hd__nor2_2 _25333_ (.A(_09424_),
    .B(_09425_),
    .Y(_09426_));
 sky130_fd_sc_hd__nor2_2 _25334_ (.A(_08895_),
    .B(_06452_),
    .Y(_09427_));
 sky130_fd_sc_hd__a2bb2o_1 _25335_ (.A1_N(_09426_),
    .A2_N(_09427_),
    .B1(_09426_),
    .B2(_09427_),
    .X(_09428_));
 sky130_fd_sc_hd__o21ba_1 _25336_ (.A1(_09294_),
    .A2(_09297_),
    .B1_N(_09296_),
    .X(_09429_));
 sky130_fd_sc_hd__a2bb2o_1 _25337_ (.A1_N(_09428_),
    .A2_N(_09429_),
    .B1(_09428_),
    .B2(_09429_),
    .X(_09430_));
 sky130_fd_sc_hd__a2bb2o_1 _25338_ (.A1_N(_09421_),
    .A2_N(_09430_),
    .B1(_09421_),
    .B2(_09430_),
    .X(_09431_));
 sky130_fd_sc_hd__a2bb2o_1 _25339_ (.A1_N(_09413_),
    .A2_N(_09431_),
    .B1(_09413_),
    .B2(_09431_),
    .X(_09432_));
 sky130_fd_sc_hd__a2bb2o_1 _25340_ (.A1_N(_09412_),
    .A2_N(_09432_),
    .B1(_09412_),
    .B2(_09432_),
    .X(_09433_));
 sky130_fd_sc_hd__a21oi_2 _25341_ (.A1(_09311_),
    .A2(_09312_),
    .B1(_09310_),
    .Y(_09434_));
 sky130_fd_sc_hd__o21ba_1 _25342_ (.A1(_09316_),
    .A2(_09319_),
    .B1_N(_09318_),
    .X(_09435_));
 sky130_fd_sc_hd__clkbuf_2 _25343_ (.A(_08599_),
    .X(_09436_));
 sky130_fd_sc_hd__o22a_1 _25344_ (.A1(_09436_),
    .A2(_08417_),
    .B1(_07268_),
    .B2(_06457_),
    .X(_09437_));
 sky130_fd_sc_hd__and4_1 _25345_ (.A(_13088_),
    .B(_06460_),
    .C(_09309_),
    .D(_06463_),
    .X(_09438_));
 sky130_fd_sc_hd__nor2_2 _25346_ (.A(_09437_),
    .B(_09438_),
    .Y(_09439_));
 sky130_fd_sc_hd__nor2_2 _25347_ (.A(_07074_),
    .B(_06219_),
    .Y(_09440_));
 sky130_fd_sc_hd__a2bb2o_1 _25348_ (.A1_N(_09439_),
    .A2_N(_09440_),
    .B1(_09439_),
    .B2(_09440_),
    .X(_09441_));
 sky130_fd_sc_hd__a2bb2o_1 _25349_ (.A1_N(_09435_),
    .A2_N(_09441_),
    .B1(_09435_),
    .B2(_09441_),
    .X(_09442_));
 sky130_fd_sc_hd__a2bb2o_1 _25350_ (.A1_N(_09434_),
    .A2_N(_09442_),
    .B1(_09434_),
    .B2(_09442_),
    .X(_09443_));
 sky130_fd_sc_hd__or2_1 _25351_ (.A(_08609_),
    .B(_06029_),
    .X(_09444_));
 sky130_fd_sc_hd__o22a_1 _25352_ (.A1(_08448_),
    .A2(_05817_),
    .B1(_08449_),
    .B2(_06484_),
    .X(_09445_));
 sky130_fd_sc_hd__and4_1 _25353_ (.A(_08451_),
    .B(_06486_),
    .C(_08452_),
    .D(_13582_),
    .X(_09446_));
 sky130_fd_sc_hd__or2_1 _25354_ (.A(_09445_),
    .B(_09446_),
    .X(_09447_));
 sky130_fd_sc_hd__a2bb2o_1 _25355_ (.A1_N(_09444_),
    .A2_N(_09447_),
    .B1(_09444_),
    .B2(_09447_),
    .X(_09448_));
 sky130_fd_sc_hd__or2_1 _25356_ (.A(_09188_),
    .B(_05723_),
    .X(_09449_));
 sky130_fd_sc_hd__and4_1 _25357_ (.A(_09190_),
    .B(_06831_),
    .C(_09191_),
    .D(_13591_),
    .X(_09450_));
 sky130_fd_sc_hd__o22a_1 _25358_ (.A1(_08777_),
    .A2(_05846_),
    .B1(_08778_),
    .B2(_06251_),
    .X(_09451_));
 sky130_fd_sc_hd__or2_1 _25359_ (.A(_09450_),
    .B(_09451_),
    .X(_09452_));
 sky130_fd_sc_hd__a2bb2o_1 _25360_ (.A1_N(_09449_),
    .A2_N(_09452_),
    .B1(_09449_),
    .B2(_09452_),
    .X(_09453_));
 sky130_fd_sc_hd__o21ba_1 _25361_ (.A1(_09321_),
    .A2(_09324_),
    .B1_N(_09322_),
    .X(_09454_));
 sky130_fd_sc_hd__a2bb2o_1 _25362_ (.A1_N(_09453_),
    .A2_N(_09454_),
    .B1(_09453_),
    .B2(_09454_),
    .X(_09455_));
 sky130_fd_sc_hd__a2bb2o_1 _25363_ (.A1_N(_09448_),
    .A2_N(_09455_),
    .B1(_09448_),
    .B2(_09455_),
    .X(_09456_));
 sky130_fd_sc_hd__o22a_1 _25364_ (.A1(_09325_),
    .A2(_09326_),
    .B1(_09320_),
    .B2(_09327_),
    .X(_09457_));
 sky130_fd_sc_hd__a2bb2o_1 _25365_ (.A1_N(_09456_),
    .A2_N(_09457_),
    .B1(_09456_),
    .B2(_09457_),
    .X(_09458_));
 sky130_fd_sc_hd__a2bb2o_1 _25366_ (.A1_N(_09443_),
    .A2_N(_09458_),
    .B1(_09443_),
    .B2(_09458_),
    .X(_09459_));
 sky130_fd_sc_hd__o22a_1 _25367_ (.A1(_09328_),
    .A2(_09329_),
    .B1(_09315_),
    .B2(_09330_),
    .X(_09460_));
 sky130_fd_sc_hd__a2bb2o_1 _25368_ (.A1_N(_09459_),
    .A2_N(_09460_),
    .B1(_09459_),
    .B2(_09460_),
    .X(_09461_));
 sky130_fd_sc_hd__a2bb2o_1 _25369_ (.A1_N(_09433_),
    .A2_N(_09461_),
    .B1(_09433_),
    .B2(_09461_),
    .X(_09462_));
 sky130_fd_sc_hd__o22a_1 _25370_ (.A1(_09331_),
    .A2(_09332_),
    .B1(_09303_),
    .B2(_09333_),
    .X(_09463_));
 sky130_fd_sc_hd__a2bb2o_1 _25371_ (.A1_N(_09462_),
    .A2_N(_09463_),
    .B1(_09462_),
    .B2(_09463_),
    .X(_09464_));
 sky130_fd_sc_hd__a2bb2o_1 _25372_ (.A1_N(_09411_),
    .A2_N(_09464_),
    .B1(_09411_),
    .B2(_09464_),
    .X(_09465_));
 sky130_fd_sc_hd__o22a_1 _25373_ (.A1(_09334_),
    .A2(_09335_),
    .B1(_09286_),
    .B2(_09336_),
    .X(_09466_));
 sky130_fd_sc_hd__a2bb2o_1 _25374_ (.A1_N(_09465_),
    .A2_N(_09466_),
    .B1(_09465_),
    .B2(_09466_),
    .X(_09467_));
 sky130_fd_sc_hd__a2bb2o_1 _25375_ (.A1_N(_09378_),
    .A2_N(_09467_),
    .B1(_09378_),
    .B2(_09467_),
    .X(_09468_));
 sky130_fd_sc_hd__o22a_1 _25376_ (.A1(_09337_),
    .A2(_09338_),
    .B1(_09255_),
    .B2(_09339_),
    .X(_09469_));
 sky130_fd_sc_hd__a2bb2o_1 _25377_ (.A1_N(_09468_),
    .A2_N(_09469_),
    .B1(_09468_),
    .B2(_09469_),
    .X(_09470_));
 sky130_fd_sc_hd__a2bb2o_1 _25378_ (.A1_N(_09355_),
    .A2_N(_09470_),
    .B1(_09355_),
    .B2(_09470_),
    .X(_09471_));
 sky130_fd_sc_hd__o22a_1 _25379_ (.A1(_09340_),
    .A2(_09341_),
    .B1(_09227_),
    .B2(_09342_),
    .X(_09472_));
 sky130_fd_sc_hd__a2bb2o_1 _25380_ (.A1_N(_09471_),
    .A2_N(_09472_),
    .B1(_09471_),
    .B2(_09472_),
    .X(_09473_));
 sky130_fd_sc_hd__a2bb2o_1 _25381_ (.A1_N(_09226_),
    .A2_N(_09473_),
    .B1(_09226_),
    .B2(_09473_),
    .X(_09474_));
 sky130_fd_sc_hd__o22a_1 _25382_ (.A1(_09343_),
    .A2(_09344_),
    .B1(_09099_),
    .B2(_09345_),
    .X(_09475_));
 sky130_fd_sc_hd__or2_1 _25383_ (.A(_09474_),
    .B(_09475_),
    .X(_09476_));
 sky130_fd_sc_hd__a21bo_1 _25384_ (.A1(_09474_),
    .A2(_09475_),
    .B1_N(_09476_),
    .X(_09477_));
 sky130_fd_sc_hd__buf_1 _25385_ (.A(_09477_),
    .X(_09478_));
 sky130_fd_sc_hd__or2_1 _25386_ (.A(_09219_),
    .B(_09347_),
    .X(_09479_));
 sky130_fd_sc_hd__or3_1 _25387_ (.A(_08953_),
    .B(_09095_),
    .C(_09479_),
    .X(_09480_));
 sky130_fd_sc_hd__or2_4 _25388_ (.A(_08956_),
    .B(_09480_),
    .X(_09481_));
 sky130_fd_sc_hd__and2_1 _25389_ (.A(_09222_),
    .B(_09346_),
    .X(_09482_));
 sky130_fd_sc_hd__o22a_1 _25390_ (.A1(_09222_),
    .A2(_09346_),
    .B1(_09218_),
    .B2(_09482_),
    .X(_09483_));
 sky130_fd_sc_hd__o221a_2 _25391_ (.A1(_09220_),
    .A2(_09479_),
    .B1(_08958_),
    .B2(_09480_),
    .C1(_09483_),
    .X(_09484_));
 sky130_fd_sc_hd__o21ai_1 _25392_ (.A1(_08328_),
    .A2(_09481_),
    .B1(_09484_),
    .Y(_09485_));
 sky130_vsdinv _25393_ (.A(_09485_),
    .Y(_09486_));
 sky130_vsdinv _25394_ (.A(_09478_),
    .Y(_09487_));
 sky130_fd_sc_hd__o22a_4 _25395_ (.A1(_09478_),
    .A2(_09486_),
    .B1(_09487_),
    .B2(_09485_),
    .X(_02659_));
 sky130_fd_sc_hd__o22a_1 _25396_ (.A1(_09471_),
    .A2(_09472_),
    .B1(_09226_),
    .B2(_09473_),
    .X(_09488_));
 sky130_fd_sc_hd__buf_2 _25397_ (.A(_09353_),
    .X(_09489_));
 sky130_fd_sc_hd__o22a_1 _25398_ (.A1(_09359_),
    .A2(_09376_),
    .B1(_09358_),
    .B2(_09377_),
    .X(_09490_));
 sky130_fd_sc_hd__or2_1 _25399_ (.A(_09353_),
    .B(_09490_),
    .X(_09491_));
 sky130_fd_sc_hd__a21bo_1 _25400_ (.A1(_09489_),
    .A2(_09490_),
    .B1_N(_09491_),
    .X(_09492_));
 sky130_fd_sc_hd__o22a_1 _25401_ (.A1(_09372_),
    .A2(_09373_),
    .B1(_09357_),
    .B2(_09374_),
    .X(_09493_));
 sky130_fd_sc_hd__o22a_1 _25402_ (.A1(_09380_),
    .A2(_09409_),
    .B1(_09379_),
    .B2(_09410_),
    .X(_09494_));
 sky130_fd_sc_hd__buf_1 _25403_ (.A(_09368_),
    .X(_09495_));
 sky130_fd_sc_hd__o22a_1 _25404_ (.A1(_09363_),
    .A2(_09495_),
    .B1(_09362_),
    .B2(_09369_),
    .X(_09496_));
 sky130_fd_sc_hd__o22a_1 _25405_ (.A1(_09390_),
    .A2(_09391_),
    .B1(_09385_),
    .B2(_09392_),
    .X(_09497_));
 sky130_fd_sc_hd__o22a_2 _25406_ (.A1(_09242_),
    .A2(_09364_),
    .B1(_09116_),
    .B2(_09365_),
    .X(_09498_));
 sky130_fd_sc_hd__buf_1 _25407_ (.A(_09498_),
    .X(_09499_));
 sky130_fd_sc_hd__a21oi_4 _25408_ (.A1(_09383_),
    .A2(_09384_),
    .B1(_09382_),
    .Y(_09500_));
 sky130_fd_sc_hd__a2bb2o_1 _25409_ (.A1_N(_09367_),
    .A2_N(_09500_),
    .B1(_09367_),
    .B2(_09500_),
    .X(_09501_));
 sky130_fd_sc_hd__a2bb2o_1 _25410_ (.A1_N(_09499_),
    .A2_N(_09501_),
    .B1(_09499_),
    .B2(_09501_),
    .X(_09502_));
 sky130_fd_sc_hd__a2bb2o_1 _25411_ (.A1_N(_09497_),
    .A2_N(_09502_),
    .B1(_09497_),
    .B2(_09502_),
    .X(_09503_));
 sky130_fd_sc_hd__a2bb2o_1 _25412_ (.A1_N(_09496_),
    .A2_N(_09503_),
    .B1(_09496_),
    .B2(_09503_),
    .X(_09504_));
 sky130_fd_sc_hd__o22a_1 _25413_ (.A1(_09361_),
    .A2(_09370_),
    .B1(_09360_),
    .B2(_09371_),
    .X(_09505_));
 sky130_fd_sc_hd__o2bb2ai_1 _25414_ (.A1_N(_09504_),
    .A2_N(_09505_),
    .B1(_09504_),
    .B2(_09505_),
    .Y(_09506_));
 sky130_fd_sc_hd__buf_1 _25415_ (.A(_09231_),
    .X(_09507_));
 sky130_fd_sc_hd__a2bb2o_2 _25416_ (.A1_N(_09375_),
    .A2_N(_09506_),
    .B1(_09507_),
    .B2(_09506_),
    .X(_09508_));
 sky130_fd_sc_hd__a2bb2o_1 _25417_ (.A1_N(_09494_),
    .A2_N(_09508_),
    .B1(_09494_),
    .B2(_09508_),
    .X(_09509_));
 sky130_fd_sc_hd__a2bb2o_1 _25418_ (.A1_N(_09493_),
    .A2_N(_09509_),
    .B1(_09493_),
    .B2(_09509_),
    .X(_09510_));
 sky130_fd_sc_hd__o22a_1 _25419_ (.A1(_09406_),
    .A2(_09407_),
    .B1(_09393_),
    .B2(_09408_),
    .X(_09511_));
 sky130_fd_sc_hd__o22a_1 _25420_ (.A1(_09413_),
    .A2(_09431_),
    .B1(_09412_),
    .B2(_09432_),
    .X(_09512_));
 sky130_fd_sc_hd__o22a_1 _25421_ (.A1(_07107_),
    .A2(_08837_),
    .B1(_07108_),
    .B2(_08033_),
    .X(_09513_));
 sky130_fd_sc_hd__and4_1 _25422_ (.A(_06962_),
    .B(_08667_),
    .C(_06963_),
    .D(_08668_),
    .X(_09514_));
 sky130_fd_sc_hd__or2_1 _25423_ (.A(_09513_),
    .B(_09514_),
    .X(_09515_));
 sky130_vsdinv _25424_ (.A(_09515_),
    .Y(_09516_));
 sky130_fd_sc_hd__or2_1 _25425_ (.A(_11701_),
    .B(_05534_),
    .X(_09517_));
 sky130_fd_sc_hd__clkbuf_2 _25426_ (.A(_09517_),
    .X(_09518_));
 sky130_fd_sc_hd__buf_1 _25427_ (.A(_09518_),
    .X(_09519_));
 sky130_fd_sc_hd__a32o_1 _25428_ (.A1(_08816_),
    .A2(\pcpi_mul.rs2[9] ),
    .A3(_09516_),
    .B1(_09515_),
    .B2(_09519_),
    .X(_09520_));
 sky130_fd_sc_hd__o22a_1 _25429_ (.A1(_08223_),
    .A2(_07732_),
    .B1(_08708_),
    .B2(_08179_),
    .X(_09521_));
 sky130_fd_sc_hd__and4_1 _25430_ (.A(_08390_),
    .B(_13523_),
    .C(_08391_),
    .D(_07876_),
    .X(_09522_));
 sky130_fd_sc_hd__nor2_2 _25431_ (.A(_09521_),
    .B(_09522_),
    .Y(_09523_));
 sky130_fd_sc_hd__nor2_2 _25432_ (.A(_08858_),
    .B(_09258_),
    .Y(_09524_));
 sky130_fd_sc_hd__a2bb2o_1 _25433_ (.A1_N(_09523_),
    .A2_N(_09524_),
    .B1(_09523_),
    .B2(_09524_),
    .X(_09525_));
 sky130_fd_sc_hd__a21oi_2 _25434_ (.A1(_09388_),
    .A2(_09389_),
    .B1(_09387_),
    .Y(_09526_));
 sky130_fd_sc_hd__a2bb2o_1 _25435_ (.A1_N(_09525_),
    .A2_N(_09526_),
    .B1(_09525_),
    .B2(_09526_),
    .X(_09527_));
 sky130_fd_sc_hd__a2bb2o_2 _25436_ (.A1_N(_09520_),
    .A2_N(_09527_),
    .B1(_09520_),
    .B2(_09527_),
    .X(_09528_));
 sky130_fd_sc_hd__a21oi_2 _25437_ (.A1(_09401_),
    .A2(_09403_),
    .B1(_09400_),
    .Y(_09529_));
 sky130_fd_sc_hd__a21oi_2 _25438_ (.A1(_09418_),
    .A2(_09420_),
    .B1(_09417_),
    .Y(_09530_));
 sky130_fd_sc_hd__o22a_1 _25439_ (.A1(_09396_),
    .A2(_07744_),
    .B1(_06094_),
    .B2(_07452_),
    .X(_09531_));
 sky130_fd_sc_hd__and4_2 _25440_ (.A(_09398_),
    .B(_07740_),
    .C(_09399_),
    .D(_07742_),
    .X(_09532_));
 sky130_fd_sc_hd__nor2_2 _25441_ (.A(_09531_),
    .B(_09532_),
    .Y(_09533_));
 sky130_fd_sc_hd__nor2_2 _25442_ (.A(_09402_),
    .B(_07327_),
    .Y(_09534_));
 sky130_fd_sc_hd__a2bb2o_1 _25443_ (.A1_N(_09533_),
    .A2_N(_09534_),
    .B1(_09533_),
    .B2(_09534_),
    .X(_09535_));
 sky130_fd_sc_hd__a2bb2o_1 _25444_ (.A1_N(_09530_),
    .A2_N(_09535_),
    .B1(_09530_),
    .B2(_09535_),
    .X(_09536_));
 sky130_fd_sc_hd__a2bb2o_1 _25445_ (.A1_N(_09529_),
    .A2_N(_09536_),
    .B1(_09529_),
    .B2(_09536_),
    .X(_09537_));
 sky130_fd_sc_hd__o22a_1 _25446_ (.A1(_09395_),
    .A2(_09404_),
    .B1(_09394_),
    .B2(_09405_),
    .X(_09538_));
 sky130_fd_sc_hd__a2bb2o_1 _25447_ (.A1_N(_09537_),
    .A2_N(_09538_),
    .B1(_09537_),
    .B2(_09538_),
    .X(_09539_));
 sky130_fd_sc_hd__a2bb2o_1 _25448_ (.A1_N(_09528_),
    .A2_N(_09539_),
    .B1(_09528_),
    .B2(_09539_),
    .X(_09540_));
 sky130_fd_sc_hd__a2bb2o_1 _25449_ (.A1_N(_09512_),
    .A2_N(_09540_),
    .B1(_09512_),
    .B2(_09540_),
    .X(_09541_));
 sky130_fd_sc_hd__a2bb2o_1 _25450_ (.A1_N(_09511_),
    .A2_N(_09541_),
    .B1(_09511_),
    .B2(_09541_),
    .X(_09542_));
 sky130_fd_sc_hd__o22a_1 _25451_ (.A1(_09428_),
    .A2(_09429_),
    .B1(_09421_),
    .B2(_09430_),
    .X(_09543_));
 sky130_fd_sc_hd__o22a_1 _25452_ (.A1(_09435_),
    .A2(_09441_),
    .B1(_09434_),
    .B2(_09442_),
    .X(_09544_));
 sky130_fd_sc_hd__clkbuf_2 _25453_ (.A(_08416_),
    .X(_09545_));
 sky130_fd_sc_hd__o22a_1 _25454_ (.A1(_09545_),
    .A2(_07482_),
    .B1(_09414_),
    .B2(_06881_),
    .X(_09546_));
 sky130_fd_sc_hd__clkbuf_2 _25455_ (.A(_08256_),
    .X(_09547_));
 sky130_fd_sc_hd__and4_2 _25456_ (.A(_09547_),
    .B(_13550_),
    .C(_09416_),
    .D(_13546_),
    .X(_09548_));
 sky130_fd_sc_hd__nor2_2 _25457_ (.A(_09546_),
    .B(_09548_),
    .Y(_09549_));
 sky130_fd_sc_hd__nor2_2 _25458_ (.A(_09419_),
    .B(_07171_),
    .Y(_09550_));
 sky130_fd_sc_hd__a2bb2o_1 _25459_ (.A1_N(_09549_),
    .A2_N(_09550_),
    .B1(_09549_),
    .B2(_09550_),
    .X(_09551_));
 sky130_fd_sc_hd__clkbuf_2 _25460_ (.A(_08261_),
    .X(_09552_));
 sky130_fd_sc_hd__o22a_1 _25461_ (.A1(_09552_),
    .A2(_09423_),
    .B1(_06802_),
    .B2(_06451_),
    .X(_09553_));
 sky130_fd_sc_hd__buf_2 _25462_ (.A(_07667_),
    .X(_09554_));
 sky130_fd_sc_hd__buf_2 _25463_ (.A(_07668_),
    .X(_09555_));
 sky130_fd_sc_hd__and4_1 _25464_ (.A(_09554_),
    .B(_06769_),
    .C(_09555_),
    .D(_08721_),
    .X(_09556_));
 sky130_fd_sc_hd__nor2_2 _25465_ (.A(_09553_),
    .B(_09556_),
    .Y(_09557_));
 sky130_fd_sc_hd__buf_2 _25466_ (.A(_06688_),
    .X(_09558_));
 sky130_fd_sc_hd__nor2_2 _25467_ (.A(_09558_),
    .B(_06576_),
    .Y(_09559_));
 sky130_fd_sc_hd__a2bb2o_1 _25468_ (.A1_N(_09557_),
    .A2_N(_09559_),
    .B1(_09557_),
    .B2(_09559_),
    .X(_09560_));
 sky130_fd_sc_hd__a21oi_2 _25469_ (.A1(_09426_),
    .A2(_09427_),
    .B1(_09425_),
    .Y(_09561_));
 sky130_fd_sc_hd__a2bb2o_1 _25470_ (.A1_N(_09560_),
    .A2_N(_09561_),
    .B1(_09560_),
    .B2(_09561_),
    .X(_09562_));
 sky130_fd_sc_hd__a2bb2o_1 _25471_ (.A1_N(_09551_),
    .A2_N(_09562_),
    .B1(_09551_),
    .B2(_09562_),
    .X(_09563_));
 sky130_fd_sc_hd__a2bb2o_1 _25472_ (.A1_N(_09544_),
    .A2_N(_09563_),
    .B1(_09544_),
    .B2(_09563_),
    .X(_09564_));
 sky130_fd_sc_hd__a2bb2o_1 _25473_ (.A1_N(_09543_),
    .A2_N(_09564_),
    .B1(_09543_),
    .B2(_09564_),
    .X(_09565_));
 sky130_fd_sc_hd__a21oi_2 _25474_ (.A1(_09439_),
    .A2(_09440_),
    .B1(_09438_),
    .Y(_09566_));
 sky130_fd_sc_hd__o21ba_1 _25475_ (.A1(_09444_),
    .A2(_09447_),
    .B1_N(_09446_),
    .X(_09567_));
 sky130_fd_sc_hd__o22a_1 _25476_ (.A1(_09306_),
    .A2(_06040_),
    .B1(_09307_),
    .B2(_06140_),
    .X(_09568_));
 sky130_fd_sc_hd__and4_1 _25477_ (.A(_13088_),
    .B(_08237_),
    .C(_09309_),
    .D(_13567_),
    .X(_09569_));
 sky130_fd_sc_hd__nor2_2 _25478_ (.A(_09568_),
    .B(_09569_),
    .Y(_09570_));
 sky130_fd_sc_hd__nor2_2 _25479_ (.A(_07074_),
    .B(_06435_),
    .Y(_09571_));
 sky130_fd_sc_hd__a2bb2o_1 _25480_ (.A1_N(_09570_),
    .A2_N(_09571_),
    .B1(_09570_),
    .B2(_09571_),
    .X(_09572_));
 sky130_fd_sc_hd__a2bb2o_1 _25481_ (.A1_N(_09567_),
    .A2_N(_09572_),
    .B1(_09567_),
    .B2(_09572_),
    .X(_09573_));
 sky130_fd_sc_hd__a2bb2o_1 _25482_ (.A1_N(_09566_),
    .A2_N(_09573_),
    .B1(_09566_),
    .B2(_09573_),
    .X(_09574_));
 sky130_fd_sc_hd__clkbuf_2 _25483_ (.A(_08285_),
    .X(_09575_));
 sky130_fd_sc_hd__o22a_1 _25484_ (.A1(_09575_),
    .A2(_05928_),
    .B1(_07679_),
    .B2(_06029_),
    .X(_09576_));
 sky130_fd_sc_hd__clkbuf_2 _25485_ (.A(_13073_),
    .X(_09577_));
 sky130_fd_sc_hd__and4_2 _25486_ (.A(_09577_),
    .B(_13583_),
    .C(_13079_),
    .D(_13580_),
    .X(_09578_));
 sky130_fd_sc_hd__nor2_2 _25487_ (.A(_09576_),
    .B(_09578_),
    .Y(_09579_));
 sky130_fd_sc_hd__buf_2 _25488_ (.A(_07681_),
    .X(_09580_));
 sky130_fd_sc_hd__nor2_2 _25489_ (.A(_09580_),
    .B(_06032_),
    .Y(_09581_));
 sky130_fd_sc_hd__a2bb2o_1 _25490_ (.A1_N(_09579_),
    .A2_N(_09581_),
    .B1(_09579_),
    .B2(_09581_),
    .X(_09582_));
 sky130_fd_sc_hd__or2_1 _25491_ (.A(_08772_),
    .B(_05725_),
    .X(_09583_));
 sky130_fd_sc_hd__and4_1 _25492_ (.A(_08774_),
    .B(_06251_),
    .C(_08775_),
    .D(_05949_),
    .X(_09584_));
 sky130_fd_sc_hd__o22a_1 _25493_ (.A1(_08925_),
    .A2(_05848_),
    .B1(_08926_),
    .B2(_05722_),
    .X(_09585_));
 sky130_fd_sc_hd__or2_1 _25494_ (.A(_09584_),
    .B(_09585_),
    .X(_09586_));
 sky130_fd_sc_hd__a2bb2o_1 _25495_ (.A1_N(_09583_),
    .A2_N(_09586_),
    .B1(_09583_),
    .B2(_09586_),
    .X(_09587_));
 sky130_fd_sc_hd__o21ba_1 _25496_ (.A1(_09449_),
    .A2(_09452_),
    .B1_N(_09450_),
    .X(_09588_));
 sky130_fd_sc_hd__a2bb2o_1 _25497_ (.A1_N(_09587_),
    .A2_N(_09588_),
    .B1(_09587_),
    .B2(_09588_),
    .X(_09589_));
 sky130_fd_sc_hd__a2bb2o_1 _25498_ (.A1_N(_09582_),
    .A2_N(_09589_),
    .B1(_09582_),
    .B2(_09589_),
    .X(_09590_));
 sky130_fd_sc_hd__o22a_1 _25499_ (.A1(_09453_),
    .A2(_09454_),
    .B1(_09448_),
    .B2(_09455_),
    .X(_09591_));
 sky130_fd_sc_hd__a2bb2o_1 _25500_ (.A1_N(_09590_),
    .A2_N(_09591_),
    .B1(_09590_),
    .B2(_09591_),
    .X(_09592_));
 sky130_fd_sc_hd__a2bb2o_1 _25501_ (.A1_N(_09574_),
    .A2_N(_09592_),
    .B1(_09574_),
    .B2(_09592_),
    .X(_09593_));
 sky130_fd_sc_hd__o22a_1 _25502_ (.A1(_09456_),
    .A2(_09457_),
    .B1(_09443_),
    .B2(_09458_),
    .X(_09594_));
 sky130_fd_sc_hd__a2bb2o_1 _25503_ (.A1_N(_09593_),
    .A2_N(_09594_),
    .B1(_09593_),
    .B2(_09594_),
    .X(_09595_));
 sky130_fd_sc_hd__a2bb2o_1 _25504_ (.A1_N(_09565_),
    .A2_N(_09595_),
    .B1(_09565_),
    .B2(_09595_),
    .X(_09596_));
 sky130_fd_sc_hd__o22a_1 _25505_ (.A1(_09459_),
    .A2(_09460_),
    .B1(_09433_),
    .B2(_09461_),
    .X(_09597_));
 sky130_fd_sc_hd__a2bb2o_1 _25506_ (.A1_N(_09596_),
    .A2_N(_09597_),
    .B1(_09596_),
    .B2(_09597_),
    .X(_09598_));
 sky130_fd_sc_hd__a2bb2o_1 _25507_ (.A1_N(_09542_),
    .A2_N(_09598_),
    .B1(_09542_),
    .B2(_09598_),
    .X(_09599_));
 sky130_fd_sc_hd__o22a_1 _25508_ (.A1(_09462_),
    .A2(_09463_),
    .B1(_09411_),
    .B2(_09464_),
    .X(_09600_));
 sky130_fd_sc_hd__a2bb2o_1 _25509_ (.A1_N(_09599_),
    .A2_N(_09600_),
    .B1(_09599_),
    .B2(_09600_),
    .X(_09601_));
 sky130_fd_sc_hd__a2bb2o_1 _25510_ (.A1_N(_09510_),
    .A2_N(_09601_),
    .B1(_09510_),
    .B2(_09601_),
    .X(_09602_));
 sky130_fd_sc_hd__o22a_1 _25511_ (.A1(_09465_),
    .A2(_09466_),
    .B1(_09378_),
    .B2(_09467_),
    .X(_09603_));
 sky130_fd_sc_hd__a2bb2o_1 _25512_ (.A1_N(_09602_),
    .A2_N(_09603_),
    .B1(_09602_),
    .B2(_09603_),
    .X(_09604_));
 sky130_fd_sc_hd__a2bb2o_1 _25513_ (.A1_N(_09492_),
    .A2_N(_09604_),
    .B1(_09492_),
    .B2(_09604_),
    .X(_09605_));
 sky130_fd_sc_hd__o22a_1 _25514_ (.A1(_09468_),
    .A2(_09469_),
    .B1(_09355_),
    .B2(_09470_),
    .X(_09606_));
 sky130_fd_sc_hd__a2bb2o_1 _25515_ (.A1_N(_09605_),
    .A2_N(_09606_),
    .B1(_09605_),
    .B2(_09606_),
    .X(_09607_));
 sky130_fd_sc_hd__a2bb2o_1 _25516_ (.A1_N(_09354_),
    .A2_N(_09607_),
    .B1(_09354_),
    .B2(_09607_),
    .X(_09608_));
 sky130_fd_sc_hd__or2_1 _25517_ (.A(_09488_),
    .B(_09608_),
    .X(_09609_));
 sky130_fd_sc_hd__a21bo_1 _25518_ (.A1(_09488_),
    .A2(_09608_),
    .B1_N(_09609_),
    .X(_09610_));
 sky130_fd_sc_hd__o21ai_1 _25519_ (.A1(_09478_),
    .A2(_09486_),
    .B1(_09476_),
    .Y(_09611_));
 sky130_fd_sc_hd__a2bb2o_1 _25520_ (.A1_N(_09610_),
    .A2_N(_09611_),
    .B1(_09610_),
    .B2(_09611_),
    .X(_02660_));
 sky130_fd_sc_hd__o22a_1 _25521_ (.A1(_09494_),
    .A2(_09508_),
    .B1(_09493_),
    .B2(_09509_),
    .X(_09612_));
 sky130_fd_sc_hd__clkbuf_2 _25522_ (.A(_09350_),
    .X(_09613_));
 sky130_fd_sc_hd__or2_1 _25523_ (.A(_09613_),
    .B(_09612_),
    .X(_09614_));
 sky130_fd_sc_hd__a21bo_1 _25524_ (.A1(_09489_),
    .A2(_09612_),
    .B1_N(_09614_),
    .X(_09615_));
 sky130_fd_sc_hd__clkbuf_2 _25525_ (.A(_09232_),
    .X(_09616_));
 sky130_fd_sc_hd__o22a_1 _25526_ (.A1(_09504_),
    .A2(_09505_),
    .B1(_09616_),
    .B2(_09506_),
    .X(_09617_));
 sky130_fd_sc_hd__o22a_1 _25527_ (.A1(_09512_),
    .A2(_09540_),
    .B1(_09511_),
    .B2(_09541_),
    .X(_09618_));
 sky130_fd_sc_hd__o22a_2 _25528_ (.A1(_09525_),
    .A2(_09526_),
    .B1(_09520_),
    .B2(_09527_),
    .X(_09619_));
 sky130_fd_sc_hd__clkbuf_1 _25529_ (.A(_09498_),
    .X(_09620_));
 sky130_fd_sc_hd__clkbuf_1 _25530_ (.A(_09367_),
    .X(_09621_));
 sky130_fd_sc_hd__o21ba_2 _25531_ (.A1(_09515_),
    .A2(_09518_),
    .B1_N(_09514_),
    .X(_09622_));
 sky130_fd_sc_hd__a2bb2o_1 _25532_ (.A1_N(_09621_),
    .A2_N(_09622_),
    .B1(_09621_),
    .B2(_09622_),
    .X(_09623_));
 sky130_fd_sc_hd__a2bb2o_1 _25533_ (.A1_N(_09620_),
    .A2_N(_09623_),
    .B1(_09620_),
    .B2(_09623_),
    .X(_09624_));
 sky130_fd_sc_hd__o2bb2ai_1 _25534_ (.A1_N(_09619_),
    .A2_N(_09624_),
    .B1(_09619_),
    .B2(_09624_),
    .Y(_09625_));
 sky130_fd_sc_hd__buf_1 _25535_ (.A(_09499_),
    .X(_09626_));
 sky130_fd_sc_hd__o22a_1 _25536_ (.A1(_09368_),
    .A2(_09500_),
    .B1(_09626_),
    .B2(_09501_),
    .X(_09627_));
 sky130_fd_sc_hd__o2bb2a_1 _25537_ (.A1_N(_09625_),
    .A2_N(_09627_),
    .B1(_09625_),
    .B2(_09627_),
    .X(_09628_));
 sky130_vsdinv _25538_ (.A(_09628_),
    .Y(_09629_));
 sky130_fd_sc_hd__o22a_1 _25539_ (.A1(_09497_),
    .A2(_09502_),
    .B1(_09496_),
    .B2(_09503_),
    .X(_09630_));
 sky130_vsdinv _25540_ (.A(_09630_),
    .Y(_09631_));
 sky130_fd_sc_hd__a22o_1 _25541_ (.A1(_09629_),
    .A2(_09630_),
    .B1(_09628_),
    .B2(_09631_),
    .X(_09632_));
 sky130_fd_sc_hd__a2bb2o_1 _25542_ (.A1_N(_09507_),
    .A2_N(_09632_),
    .B1(_09356_),
    .B2(_09632_),
    .X(_09633_));
 sky130_fd_sc_hd__a2bb2o_1 _25543_ (.A1_N(_09618_),
    .A2_N(_09633_),
    .B1(_09618_),
    .B2(_09633_),
    .X(_09634_));
 sky130_fd_sc_hd__a2bb2o_1 _25544_ (.A1_N(_09617_),
    .A2_N(_09634_),
    .B1(_09617_),
    .B2(_09634_),
    .X(_09635_));
 sky130_fd_sc_hd__o22a_1 _25545_ (.A1(_09537_),
    .A2(_09538_),
    .B1(_09528_),
    .B2(_09539_),
    .X(_09636_));
 sky130_fd_sc_hd__o22a_1 _25546_ (.A1(_09544_),
    .A2(_09563_),
    .B1(_09543_),
    .B2(_09564_),
    .X(_09637_));
 sky130_fd_sc_hd__nor2_1 _25547_ (.A(_08537_),
    .B(_08497_),
    .Y(_09638_));
 sky130_fd_sc_hd__or2_2 _25548_ (.A(_09241_),
    .B(_05585_),
    .X(_09639_));
 sky130_vsdinv _25549_ (.A(_09639_),
    .Y(_09640_));
 sky130_fd_sc_hd__a2bb2o_1 _25550_ (.A1_N(_09638_),
    .A2_N(_09640_),
    .B1(_09638_),
    .B2(_09640_),
    .X(_09641_));
 sky130_fd_sc_hd__a2bb2o_1 _25551_ (.A1_N(_09519_),
    .A2_N(_09641_),
    .B1(_09519_),
    .B2(_09641_),
    .X(_09642_));
 sky130_fd_sc_hd__o22a_1 _25552_ (.A1(_08544_),
    .A2(_08179_),
    .B1(_08708_),
    .B2(_07872_),
    .X(_09643_));
 sky130_fd_sc_hd__and4_2 _25553_ (.A(_08547_),
    .B(_07876_),
    .C(_08548_),
    .D(_08022_),
    .X(_09644_));
 sky130_fd_sc_hd__nor2_2 _25554_ (.A(_09643_),
    .B(_09644_),
    .Y(_09645_));
 sky130_fd_sc_hd__nor2_2 _25555_ (.A(_05709_),
    .B(_07891_),
    .Y(_09646_));
 sky130_fd_sc_hd__a2bb2o_1 _25556_ (.A1_N(_09645_),
    .A2_N(_09646_),
    .B1(_09645_),
    .B2(_09646_),
    .X(_09647_));
 sky130_fd_sc_hd__a21oi_2 _25557_ (.A1(_09523_),
    .A2(_09524_),
    .B1(_09522_),
    .Y(_09648_));
 sky130_fd_sc_hd__a2bb2o_1 _25558_ (.A1_N(_09647_),
    .A2_N(_09648_),
    .B1(_09647_),
    .B2(_09648_),
    .X(_09649_));
 sky130_fd_sc_hd__a2bb2o_2 _25559_ (.A1_N(_09642_),
    .A2_N(_09649_),
    .B1(_09642_),
    .B2(_09649_),
    .X(_09650_));
 sky130_fd_sc_hd__a21oi_2 _25560_ (.A1(_09533_),
    .A2(_09534_),
    .B1(_09532_),
    .Y(_09651_));
 sky130_fd_sc_hd__a21oi_2 _25561_ (.A1(_09549_),
    .A2(_09550_),
    .B1(_09548_),
    .Y(_09652_));
 sky130_fd_sc_hd__o22a_1 _25562_ (.A1(_08869_),
    .A2(_07452_),
    .B1(_08870_),
    .B2(_07326_),
    .X(_09653_));
 sky130_fd_sc_hd__and4_2 _25563_ (.A(_08872_),
    .B(_07742_),
    .C(_08873_),
    .D(_07449_),
    .X(_09654_));
 sky130_fd_sc_hd__nor2_2 _25564_ (.A(_09653_),
    .B(_09654_),
    .Y(_09655_));
 sky130_fd_sc_hd__nor2_2 _25565_ (.A(_09147_),
    .B(_07464_),
    .Y(_09656_));
 sky130_fd_sc_hd__a2bb2o_1 _25566_ (.A1_N(_09655_),
    .A2_N(_09656_),
    .B1(_09655_),
    .B2(_09656_),
    .X(_09657_));
 sky130_fd_sc_hd__a2bb2o_1 _25567_ (.A1_N(_09652_),
    .A2_N(_09657_),
    .B1(_09652_),
    .B2(_09657_),
    .X(_09658_));
 sky130_fd_sc_hd__a2bb2o_1 _25568_ (.A1_N(_09651_),
    .A2_N(_09658_),
    .B1(_09651_),
    .B2(_09658_),
    .X(_09659_));
 sky130_fd_sc_hd__o22a_1 _25569_ (.A1(_09530_),
    .A2(_09535_),
    .B1(_09529_),
    .B2(_09536_),
    .X(_09660_));
 sky130_fd_sc_hd__a2bb2o_1 _25570_ (.A1_N(_09659_),
    .A2_N(_09660_),
    .B1(_09659_),
    .B2(_09660_),
    .X(_09661_));
 sky130_fd_sc_hd__a2bb2o_1 _25571_ (.A1_N(_09650_),
    .A2_N(_09661_),
    .B1(_09650_),
    .B2(_09661_),
    .X(_09662_));
 sky130_fd_sc_hd__a2bb2o_1 _25572_ (.A1_N(_09637_),
    .A2_N(_09662_),
    .B1(_09637_),
    .B2(_09662_),
    .X(_09663_));
 sky130_fd_sc_hd__a2bb2o_1 _25573_ (.A1_N(_09636_),
    .A2_N(_09663_),
    .B1(_09636_),
    .B2(_09663_),
    .X(_09664_));
 sky130_fd_sc_hd__o22a_1 _25574_ (.A1(_09560_),
    .A2(_09561_),
    .B1(_09551_),
    .B2(_09562_),
    .X(_09665_));
 sky130_fd_sc_hd__o22a_1 _25575_ (.A1(_09567_),
    .A2(_09572_),
    .B1(_09566_),
    .B2(_09573_),
    .X(_09666_));
 sky130_fd_sc_hd__o22a_1 _25576_ (.A1(_09545_),
    .A2(_07613_),
    .B1(_09414_),
    .B2(_07170_),
    .X(_09667_));
 sky130_fd_sc_hd__and4_2 _25577_ (.A(_09547_),
    .B(_13546_),
    .C(_09416_),
    .D(_13542_),
    .X(_09668_));
 sky130_fd_sc_hd__nor2_2 _25578_ (.A(_09667_),
    .B(_09668_),
    .Y(_09669_));
 sky130_fd_sc_hd__nor2_2 _25579_ (.A(_09419_),
    .B(_07034_),
    .Y(_09670_));
 sky130_fd_sc_hd__a2bb2o_1 _25580_ (.A1_N(_09669_),
    .A2_N(_09670_),
    .B1(_09669_),
    .B2(_09670_),
    .X(_09671_));
 sky130_fd_sc_hd__o22a_1 _25581_ (.A1(_09552_),
    .A2(_08719_),
    .B1(_09422_),
    .B2(_06575_),
    .X(_09672_));
 sky130_fd_sc_hd__and4_1 _25582_ (.A(_09554_),
    .B(_08721_),
    .C(_09555_),
    .D(_07040_),
    .X(_09673_));
 sky130_fd_sc_hd__nor2_2 _25583_ (.A(_09672_),
    .B(_09673_),
    .Y(_09674_));
 sky130_fd_sc_hd__nor2_2 _25584_ (.A(_09558_),
    .B(_06651_),
    .Y(_09675_));
 sky130_fd_sc_hd__a2bb2o_1 _25585_ (.A1_N(_09674_),
    .A2_N(_09675_),
    .B1(_09674_),
    .B2(_09675_),
    .X(_09676_));
 sky130_fd_sc_hd__a21oi_2 _25586_ (.A1(_09557_),
    .A2(_09559_),
    .B1(_09556_),
    .Y(_09677_));
 sky130_fd_sc_hd__a2bb2o_1 _25587_ (.A1_N(_09676_),
    .A2_N(_09677_),
    .B1(_09676_),
    .B2(_09677_),
    .X(_09678_));
 sky130_fd_sc_hd__a2bb2o_1 _25588_ (.A1_N(_09671_),
    .A2_N(_09678_),
    .B1(_09671_),
    .B2(_09678_),
    .X(_09679_));
 sky130_fd_sc_hd__a2bb2o_1 _25589_ (.A1_N(_09666_),
    .A2_N(_09679_),
    .B1(_09666_),
    .B2(_09679_),
    .X(_09680_));
 sky130_fd_sc_hd__a2bb2o_1 _25590_ (.A1_N(_09665_),
    .A2_N(_09680_),
    .B1(_09665_),
    .B2(_09680_),
    .X(_09681_));
 sky130_fd_sc_hd__a21oi_2 _25591_ (.A1(_09570_),
    .A2(_09571_),
    .B1(_09569_),
    .Y(_09682_));
 sky130_fd_sc_hd__a21oi_2 _25592_ (.A1(_09579_),
    .A2(_09581_),
    .B1(_09578_),
    .Y(_09683_));
 sky130_fd_sc_hd__o22a_1 _25593_ (.A1(_09306_),
    .A2(_06140_),
    .B1(_09307_),
    .B2(_06434_),
    .X(_09684_));
 sky130_fd_sc_hd__and4_1 _25594_ (.A(_08761_),
    .B(_13567_),
    .C(_09309_),
    .D(_06654_),
    .X(_09685_));
 sky130_fd_sc_hd__nor2_2 _25595_ (.A(_09684_),
    .B(_09685_),
    .Y(_09686_));
 sky130_fd_sc_hd__nor2_2 _25596_ (.A(_08758_),
    .B(_08887_),
    .Y(_09687_));
 sky130_fd_sc_hd__a2bb2o_1 _25597_ (.A1_N(_09686_),
    .A2_N(_09687_),
    .B1(_09686_),
    .B2(_09687_),
    .X(_09688_));
 sky130_fd_sc_hd__a2bb2o_1 _25598_ (.A1_N(_09683_),
    .A2_N(_09688_),
    .B1(_09683_),
    .B2(_09688_),
    .X(_09689_));
 sky130_fd_sc_hd__a2bb2o_1 _25599_ (.A1_N(_09682_),
    .A2_N(_09689_),
    .B1(_09682_),
    .B2(_09689_),
    .X(_09690_));
 sky130_fd_sc_hd__o22a_1 _25600_ (.A1(_08611_),
    .A2(_06479_),
    .B1(_07679_),
    .B2(_06599_),
    .X(_09691_));
 sky130_fd_sc_hd__and4_1 _25601_ (.A(_09577_),
    .B(_08747_),
    .C(_13079_),
    .D(_06460_),
    .X(_09692_));
 sky130_fd_sc_hd__nor2_2 _25602_ (.A(_09691_),
    .B(_09692_),
    .Y(_09693_));
 sky130_fd_sc_hd__nor2_2 _25603_ (.A(_09580_),
    .B(_06334_),
    .Y(_09694_));
 sky130_fd_sc_hd__a2bb2o_1 _25604_ (.A1_N(_09693_),
    .A2_N(_09694_),
    .B1(_09693_),
    .B2(_09694_),
    .X(_09695_));
 sky130_fd_sc_hd__or2_1 _25605_ (.A(_08921_),
    .B(_06702_),
    .X(_09696_));
 sky130_fd_sc_hd__and4_1 _25606_ (.A(_09067_),
    .B(_05722_),
    .C(_08923_),
    .D(_13584_),
    .X(_09697_));
 sky130_fd_sc_hd__o22a_1 _25607_ (.A1(_08620_),
    .A2(_05949_),
    .B1(_09069_),
    .B2(_06043_),
    .X(_09698_));
 sky130_fd_sc_hd__or2_1 _25608_ (.A(_09697_),
    .B(_09698_),
    .X(_09699_));
 sky130_fd_sc_hd__a2bb2o_1 _25609_ (.A1_N(_09696_),
    .A2_N(_09699_),
    .B1(_09696_),
    .B2(_09699_),
    .X(_09700_));
 sky130_fd_sc_hd__o21ba_1 _25610_ (.A1(_09583_),
    .A2(_09586_),
    .B1_N(_09584_),
    .X(_09701_));
 sky130_fd_sc_hd__a2bb2o_1 _25611_ (.A1_N(_09700_),
    .A2_N(_09701_),
    .B1(_09700_),
    .B2(_09701_),
    .X(_09702_));
 sky130_fd_sc_hd__a2bb2o_1 _25612_ (.A1_N(_09695_),
    .A2_N(_09702_),
    .B1(_09695_),
    .B2(_09702_),
    .X(_09703_));
 sky130_fd_sc_hd__o22a_1 _25613_ (.A1(_09587_),
    .A2(_09588_),
    .B1(_09582_),
    .B2(_09589_),
    .X(_09704_));
 sky130_fd_sc_hd__a2bb2o_1 _25614_ (.A1_N(_09703_),
    .A2_N(_09704_),
    .B1(_09703_),
    .B2(_09704_),
    .X(_09705_));
 sky130_fd_sc_hd__a2bb2o_1 _25615_ (.A1_N(_09690_),
    .A2_N(_09705_),
    .B1(_09690_),
    .B2(_09705_),
    .X(_09706_));
 sky130_fd_sc_hd__o22a_1 _25616_ (.A1(_09590_),
    .A2(_09591_),
    .B1(_09574_),
    .B2(_09592_),
    .X(_09707_));
 sky130_fd_sc_hd__a2bb2o_1 _25617_ (.A1_N(_09706_),
    .A2_N(_09707_),
    .B1(_09706_),
    .B2(_09707_),
    .X(_09708_));
 sky130_fd_sc_hd__a2bb2o_1 _25618_ (.A1_N(_09681_),
    .A2_N(_09708_),
    .B1(_09681_),
    .B2(_09708_),
    .X(_09709_));
 sky130_fd_sc_hd__o22a_1 _25619_ (.A1(_09593_),
    .A2(_09594_),
    .B1(_09565_),
    .B2(_09595_),
    .X(_09710_));
 sky130_fd_sc_hd__a2bb2o_1 _25620_ (.A1_N(_09709_),
    .A2_N(_09710_),
    .B1(_09709_),
    .B2(_09710_),
    .X(_09711_));
 sky130_fd_sc_hd__a2bb2o_1 _25621_ (.A1_N(_09664_),
    .A2_N(_09711_),
    .B1(_09664_),
    .B2(_09711_),
    .X(_09712_));
 sky130_fd_sc_hd__o22a_1 _25622_ (.A1(_09596_),
    .A2(_09597_),
    .B1(_09542_),
    .B2(_09598_),
    .X(_09713_));
 sky130_fd_sc_hd__a2bb2o_1 _25623_ (.A1_N(_09712_),
    .A2_N(_09713_),
    .B1(_09712_),
    .B2(_09713_),
    .X(_09714_));
 sky130_fd_sc_hd__a2bb2o_1 _25624_ (.A1_N(_09635_),
    .A2_N(_09714_),
    .B1(_09635_),
    .B2(_09714_),
    .X(_09715_));
 sky130_fd_sc_hd__o22a_1 _25625_ (.A1(_09599_),
    .A2(_09600_),
    .B1(_09510_),
    .B2(_09601_),
    .X(_09716_));
 sky130_fd_sc_hd__a2bb2o_1 _25626_ (.A1_N(_09715_),
    .A2_N(_09716_),
    .B1(_09715_),
    .B2(_09716_),
    .X(_09717_));
 sky130_fd_sc_hd__a2bb2o_1 _25627_ (.A1_N(_09615_),
    .A2_N(_09717_),
    .B1(_09615_),
    .B2(_09717_),
    .X(_09718_));
 sky130_fd_sc_hd__o22a_1 _25628_ (.A1(_09602_),
    .A2(_09603_),
    .B1(_09492_),
    .B2(_09604_),
    .X(_09719_));
 sky130_fd_sc_hd__a2bb2o_1 _25629_ (.A1_N(_09718_),
    .A2_N(_09719_),
    .B1(_09718_),
    .B2(_09719_),
    .X(_09720_));
 sky130_fd_sc_hd__a2bb2o_1 _25630_ (.A1_N(_09491_),
    .A2_N(_09720_),
    .B1(_09491_),
    .B2(_09720_),
    .X(_09721_));
 sky130_fd_sc_hd__o22a_1 _25631_ (.A1(_09605_),
    .A2(_09606_),
    .B1(_09354_),
    .B2(_09607_),
    .X(_09722_));
 sky130_fd_sc_hd__or2_1 _25632_ (.A(_09721_),
    .B(_09722_),
    .X(_09723_));
 sky130_fd_sc_hd__a21bo_1 _25633_ (.A1(_09721_),
    .A2(_09722_),
    .B1_N(_09723_),
    .X(_09724_));
 sky130_fd_sc_hd__a22o_1 _25634_ (.A1(_09488_),
    .A2(_09608_),
    .B1(_09476_),
    .B2(_09609_),
    .X(_09725_));
 sky130_fd_sc_hd__o31a_1 _25635_ (.A1(_09478_),
    .A2(_09610_),
    .A3(_09486_),
    .B1(_09725_),
    .X(_09726_));
 sky130_fd_sc_hd__a2bb2oi_1 _25636_ (.A1_N(_09724_),
    .A2_N(_09726_),
    .B1(_09724_),
    .B2(_09726_),
    .Y(_02661_));
 sky130_fd_sc_hd__o22a_1 _25637_ (.A1(_09718_),
    .A2(_09719_),
    .B1(_09491_),
    .B2(_09720_),
    .X(_09727_));
 sky130_fd_sc_hd__o22a_1 _25638_ (.A1(_09618_),
    .A2(_09633_),
    .B1(_09617_),
    .B2(_09634_),
    .X(_09728_));
 sky130_fd_sc_hd__or2_1 _25639_ (.A(_09613_),
    .B(_09728_),
    .X(_09729_));
 sky130_fd_sc_hd__a21bo_1 _25640_ (.A1(_09351_),
    .A2(_09728_),
    .B1_N(_09729_),
    .X(_09730_));
 sky130_fd_sc_hd__o22a_1 _25641_ (.A1(_09629_),
    .A2(_09630_),
    .B1(_09357_),
    .B2(_09632_),
    .X(_09731_));
 sky130_fd_sc_hd__o22a_1 _25642_ (.A1(_09637_),
    .A2(_09662_),
    .B1(_09636_),
    .B2(_09663_),
    .X(_09732_));
 sky130_fd_sc_hd__o22a_2 _25643_ (.A1(_09647_),
    .A2(_09648_),
    .B1(_09642_),
    .B2(_09649_),
    .X(_09733_));
 sky130_fd_sc_hd__o32a_4 _25644_ (.A1(_09003_),
    .A2(_08498_),
    .A3(_09639_),
    .B1(_09518_),
    .B2(_09641_),
    .X(_09734_));
 sky130_fd_sc_hd__a2bb2o_1 _25645_ (.A1_N(_09621_),
    .A2_N(_09734_),
    .B1(_09621_),
    .B2(_09734_),
    .X(_09735_));
 sky130_fd_sc_hd__a2bb2o_1 _25646_ (.A1_N(_09620_),
    .A2_N(_09735_),
    .B1(_09620_),
    .B2(_09735_),
    .X(_09736_));
 sky130_fd_sc_hd__o2bb2ai_1 _25647_ (.A1_N(_09733_),
    .A2_N(_09736_),
    .B1(_09733_),
    .B2(_09736_),
    .Y(_09737_));
 sky130_fd_sc_hd__buf_1 _25648_ (.A(_09499_),
    .X(_09738_));
 sky130_fd_sc_hd__o22a_1 _25649_ (.A1(_09495_),
    .A2(_09622_),
    .B1(_09738_),
    .B2(_09623_),
    .X(_09739_));
 sky130_fd_sc_hd__o2bb2a_1 _25650_ (.A1_N(_09737_),
    .A2_N(_09739_),
    .B1(_09737_),
    .B2(_09739_),
    .X(_09740_));
 sky130_vsdinv _25651_ (.A(_09740_),
    .Y(_09741_));
 sky130_fd_sc_hd__o22a_1 _25652_ (.A1(_09619_),
    .A2(_09624_),
    .B1(_09625_),
    .B2(_09627_),
    .X(_09742_));
 sky130_vsdinv _25653_ (.A(_09742_),
    .Y(_09743_));
 sky130_fd_sc_hd__a22o_1 _25654_ (.A1(_09741_),
    .A2(_09742_),
    .B1(_09740_),
    .B2(_09743_),
    .X(_09744_));
 sky130_fd_sc_hd__a2bb2o_1 _25655_ (.A1_N(_09252_),
    .A2_N(_09744_),
    .B1(_09252_),
    .B2(_09744_),
    .X(_09745_));
 sky130_fd_sc_hd__a2bb2o_1 _25656_ (.A1_N(_09732_),
    .A2_N(_09745_),
    .B1(_09732_),
    .B2(_09745_),
    .X(_09746_));
 sky130_fd_sc_hd__a2bb2o_1 _25657_ (.A1_N(_09731_),
    .A2_N(_09746_),
    .B1(_09731_),
    .B2(_09746_),
    .X(_09747_));
 sky130_fd_sc_hd__o22a_1 _25658_ (.A1(_09659_),
    .A2(_09660_),
    .B1(_09650_),
    .B2(_09661_),
    .X(_09748_));
 sky130_fd_sc_hd__o22a_2 _25659_ (.A1(_09666_),
    .A2(_09679_),
    .B1(_09665_),
    .B2(_09680_),
    .X(_09749_));
 sky130_fd_sc_hd__or2_1 _25660_ (.A(_09241_),
    .B(_05649_),
    .X(_09750_));
 sky130_fd_sc_hd__a32o_1 _25661_ (.A1(\pcpi_mul.rs1[32] ),
    .A2(_13135_),
    .A3(_09640_),
    .B1(_09639_),
    .B2(_09750_),
    .X(_09751_));
 sky130_fd_sc_hd__a2bb2o_2 _25662_ (.A1_N(_09519_),
    .A2_N(_09751_),
    .B1(_09518_),
    .B2(_09751_),
    .X(_09752_));
 sky130_fd_sc_hd__buf_1 _25663_ (.A(_09752_),
    .X(_09753_));
 sky130_fd_sc_hd__buf_1 _25664_ (.A(_09753_),
    .X(_09754_));
 sky130_fd_sc_hd__o22a_1 _25665_ (.A1(_06710_),
    .A2(_07747_),
    .B1(_06533_),
    .B2(_07889_),
    .X(_09755_));
 sky130_fd_sc_hd__and4_2 _25666_ (.A(_13129_),
    .B(\pcpi_mul.rs1[29] ),
    .C(_13132_),
    .D(\pcpi_mul.rs1[30] ),
    .X(_09756_));
 sky130_fd_sc_hd__nor2_2 _25667_ (.A(_09755_),
    .B(_09756_),
    .Y(_09757_));
 sky130_fd_sc_hd__nor2_1 _25668_ (.A(_05709_),
    .B(_09239_),
    .Y(_09758_));
 sky130_fd_sc_hd__a2bb2o_1 _25669_ (.A1_N(_09757_),
    .A2_N(_09758_),
    .B1(_09757_),
    .B2(_09758_),
    .X(_09759_));
 sky130_fd_sc_hd__a21oi_2 _25670_ (.A1(_09645_),
    .A2(_09646_),
    .B1(_09644_),
    .Y(_09760_));
 sky130_fd_sc_hd__a2bb2o_1 _25671_ (.A1_N(_09759_),
    .A2_N(_09760_),
    .B1(_09759_),
    .B2(_09760_),
    .X(_09761_));
 sky130_fd_sc_hd__a2bb2o_1 _25672_ (.A1_N(_09754_),
    .A2_N(_09761_),
    .B1(_09754_),
    .B2(_09761_),
    .X(_09762_));
 sky130_fd_sc_hd__a21oi_2 _25673_ (.A1(_09655_),
    .A2(_09656_),
    .B1(_09654_),
    .Y(_09763_));
 sky130_fd_sc_hd__a21oi_2 _25674_ (.A1(_09669_),
    .A2(_09670_),
    .B1(_09668_),
    .Y(_09764_));
 sky130_fd_sc_hd__o22a_1 _25675_ (.A1(_09396_),
    .A2(_08364_),
    .B1(_09274_),
    .B2(_08684_),
    .X(_09765_));
 sky130_fd_sc_hd__and4_2 _25676_ (.A(_09398_),
    .B(_13528_),
    .C(_09399_),
    .D(_07587_),
    .X(_09766_));
 sky130_fd_sc_hd__nor2_2 _25677_ (.A(_09765_),
    .B(_09766_),
    .Y(_09767_));
 sky130_fd_sc_hd__nor2_2 _25678_ (.A(_09147_),
    .B(_07871_),
    .Y(_09768_));
 sky130_fd_sc_hd__a2bb2o_1 _25679_ (.A1_N(_09767_),
    .A2_N(_09768_),
    .B1(_09767_),
    .B2(_09768_),
    .X(_09769_));
 sky130_fd_sc_hd__a2bb2o_1 _25680_ (.A1_N(_09764_),
    .A2_N(_09769_),
    .B1(_09764_),
    .B2(_09769_),
    .X(_09770_));
 sky130_fd_sc_hd__a2bb2o_1 _25681_ (.A1_N(_09763_),
    .A2_N(_09770_),
    .B1(_09763_),
    .B2(_09770_),
    .X(_09771_));
 sky130_fd_sc_hd__o22a_1 _25682_ (.A1(_09652_),
    .A2(_09657_),
    .B1(_09651_),
    .B2(_09658_),
    .X(_09772_));
 sky130_fd_sc_hd__a2bb2o_1 _25683_ (.A1_N(_09771_),
    .A2_N(_09772_),
    .B1(_09771_),
    .B2(_09772_),
    .X(_09773_));
 sky130_fd_sc_hd__a2bb2o_1 _25684_ (.A1_N(_09762_),
    .A2_N(_09773_),
    .B1(_09762_),
    .B2(_09773_),
    .X(_09774_));
 sky130_fd_sc_hd__a2bb2o_1 _25685_ (.A1_N(_09749_),
    .A2_N(_09774_),
    .B1(_09749_),
    .B2(_09774_),
    .X(_09775_));
 sky130_fd_sc_hd__a2bb2o_1 _25686_ (.A1_N(_09748_),
    .A2_N(_09775_),
    .B1(_09748_),
    .B2(_09775_),
    .X(_09776_));
 sky130_fd_sc_hd__o22a_1 _25687_ (.A1(_09676_),
    .A2(_09677_),
    .B1(_09671_),
    .B2(_09678_),
    .X(_09777_));
 sky130_fd_sc_hd__o22a_1 _25688_ (.A1(_09683_),
    .A2(_09688_),
    .B1(_09682_),
    .B2(_09689_),
    .X(_09778_));
 sky130_fd_sc_hd__o22a_1 _25689_ (.A1(_08889_),
    .A2(_07170_),
    .B1(_09414_),
    .B2(_07172_),
    .X(_09779_));
 sky130_fd_sc_hd__and4_2 _25690_ (.A(_09547_),
    .B(_07466_),
    .C(_09416_),
    .D(_13539_),
    .X(_09780_));
 sky130_fd_sc_hd__nor2_2 _25691_ (.A(_09779_),
    .B(_09780_),
    .Y(_09781_));
 sky130_fd_sc_hd__buf_1 _25692_ (.A(_07196_),
    .X(_09782_));
 sky130_fd_sc_hd__buf_2 _25693_ (.A(_09782_),
    .X(_09783_));
 sky130_fd_sc_hd__nor2_2 _25694_ (.A(_09419_),
    .B(_09783_),
    .Y(_09784_));
 sky130_fd_sc_hd__a2bb2o_1 _25695_ (.A1_N(_09781_),
    .A2_N(_09784_),
    .B1(_09781_),
    .B2(_09784_),
    .X(_09785_));
 sky130_fd_sc_hd__o22a_1 _25696_ (.A1(_08897_),
    .A2(_06575_),
    .B1(_09422_),
    .B2(_07762_),
    .X(_09786_));
 sky130_fd_sc_hd__and4_1 _25697_ (.A(_09554_),
    .B(_07187_),
    .C(_09555_),
    .D(_07191_),
    .X(_09787_));
 sky130_fd_sc_hd__nor2_2 _25698_ (.A(_09786_),
    .B(_09787_),
    .Y(_09788_));
 sky130_fd_sc_hd__nor2_2 _25699_ (.A(_09558_),
    .B(_06763_),
    .Y(_09789_));
 sky130_fd_sc_hd__a2bb2o_1 _25700_ (.A1_N(_09788_),
    .A2_N(_09789_),
    .B1(_09788_),
    .B2(_09789_),
    .X(_09790_));
 sky130_fd_sc_hd__a21oi_2 _25701_ (.A1(_09674_),
    .A2(_09675_),
    .B1(_09673_),
    .Y(_09791_));
 sky130_fd_sc_hd__a2bb2o_1 _25702_ (.A1_N(_09790_),
    .A2_N(_09791_),
    .B1(_09790_),
    .B2(_09791_),
    .X(_09792_));
 sky130_fd_sc_hd__a2bb2o_1 _25703_ (.A1_N(_09785_),
    .A2_N(_09792_),
    .B1(_09785_),
    .B2(_09792_),
    .X(_09793_));
 sky130_fd_sc_hd__a2bb2o_1 _25704_ (.A1_N(_09778_),
    .A2_N(_09793_),
    .B1(_09778_),
    .B2(_09793_),
    .X(_09794_));
 sky130_fd_sc_hd__a2bb2o_1 _25705_ (.A1_N(_09777_),
    .A2_N(_09794_),
    .B1(_09777_),
    .B2(_09794_),
    .X(_09795_));
 sky130_fd_sc_hd__a21oi_2 _25706_ (.A1(_09686_),
    .A2(_09687_),
    .B1(_09685_),
    .Y(_09796_));
 sky130_fd_sc_hd__a21oi_2 _25707_ (.A1(_09693_),
    .A2(_09694_),
    .B1(_09692_),
    .Y(_09797_));
 sky130_fd_sc_hd__o22a_1 _25708_ (.A1(_09306_),
    .A2(_08890_),
    .B1(_09307_),
    .B2(_09423_),
    .X(_09798_));
 sky130_fd_sc_hd__and4_1 _25709_ (.A(_08761_),
    .B(_06654_),
    .C(_13092_),
    .D(_06769_),
    .X(_09799_));
 sky130_fd_sc_hd__nor2_2 _25710_ (.A(_09798_),
    .B(_09799_),
    .Y(_09800_));
 sky130_fd_sc_hd__nor2_2 _25711_ (.A(_08758_),
    .B(_08557_),
    .Y(_09801_));
 sky130_fd_sc_hd__a2bb2o_1 _25712_ (.A1_N(_09800_),
    .A2_N(_09801_),
    .B1(_09800_),
    .B2(_09801_),
    .X(_09802_));
 sky130_fd_sc_hd__a2bb2o_1 _25713_ (.A1_N(_09797_),
    .A2_N(_09802_),
    .B1(_09797_),
    .B2(_09802_),
    .X(_09803_));
 sky130_fd_sc_hd__a2bb2o_1 _25714_ (.A1_N(_09796_),
    .A2_N(_09803_),
    .B1(_09796_),
    .B2(_09803_),
    .X(_09804_));
 sky130_fd_sc_hd__o22a_1 _25715_ (.A1(_09575_),
    .A2(_05944_),
    .B1(_07679_),
    .B2(_06132_),
    .X(_09805_));
 sky130_fd_sc_hd__buf_1 _25716_ (.A(_08452_),
    .X(_09806_));
 sky130_fd_sc_hd__and4_2 _25717_ (.A(_09577_),
    .B(_13576_),
    .C(_09806_),
    .D(_06463_),
    .X(_09807_));
 sky130_fd_sc_hd__nor2_2 _25718_ (.A(_09805_),
    .B(_09807_),
    .Y(_09808_));
 sky130_fd_sc_hd__nor2_2 _25719_ (.A(_09580_),
    .B(_06219_),
    .Y(_09809_));
 sky130_fd_sc_hd__a2bb2o_1 _25720_ (.A1_N(_09808_),
    .A2_N(_09809_),
    .B1(_09808_),
    .B2(_09809_),
    .X(_09810_));
 sky130_fd_sc_hd__or2_1 _25721_ (.A(_08921_),
    .B(_05837_),
    .X(_09811_));
 sky130_fd_sc_hd__and4_1 _25722_ (.A(_09067_),
    .B(_05724_),
    .C(_08923_),
    .D(_06145_),
    .X(_09812_));
 sky130_fd_sc_hd__o22a_1 _25723_ (.A1(_08620_),
    .A2(_06144_),
    .B1(_09069_),
    .B2(_05819_),
    .X(_09813_));
 sky130_fd_sc_hd__or2_1 _25724_ (.A(_09812_),
    .B(_09813_),
    .X(_09814_));
 sky130_fd_sc_hd__a2bb2o_1 _25725_ (.A1_N(_09811_),
    .A2_N(_09814_),
    .B1(_09811_),
    .B2(_09814_),
    .X(_09815_));
 sky130_fd_sc_hd__o21ba_1 _25726_ (.A1(_09696_),
    .A2(_09699_),
    .B1_N(_09697_),
    .X(_09816_));
 sky130_fd_sc_hd__a2bb2o_1 _25727_ (.A1_N(_09815_),
    .A2_N(_09816_),
    .B1(_09815_),
    .B2(_09816_),
    .X(_09817_));
 sky130_fd_sc_hd__a2bb2o_1 _25728_ (.A1_N(_09810_),
    .A2_N(_09817_),
    .B1(_09810_),
    .B2(_09817_),
    .X(_09818_));
 sky130_fd_sc_hd__o22a_1 _25729_ (.A1(_09700_),
    .A2(_09701_),
    .B1(_09695_),
    .B2(_09702_),
    .X(_09819_));
 sky130_fd_sc_hd__a2bb2o_1 _25730_ (.A1_N(_09818_),
    .A2_N(_09819_),
    .B1(_09818_),
    .B2(_09819_),
    .X(_09820_));
 sky130_fd_sc_hd__a2bb2o_1 _25731_ (.A1_N(_09804_),
    .A2_N(_09820_),
    .B1(_09804_),
    .B2(_09820_),
    .X(_09821_));
 sky130_fd_sc_hd__o22a_1 _25732_ (.A1(_09703_),
    .A2(_09704_),
    .B1(_09690_),
    .B2(_09705_),
    .X(_09822_));
 sky130_fd_sc_hd__a2bb2o_1 _25733_ (.A1_N(_09821_),
    .A2_N(_09822_),
    .B1(_09821_),
    .B2(_09822_),
    .X(_09823_));
 sky130_fd_sc_hd__a2bb2o_2 _25734_ (.A1_N(_09795_),
    .A2_N(_09823_),
    .B1(_09795_),
    .B2(_09823_),
    .X(_09824_));
 sky130_fd_sc_hd__o22a_2 _25735_ (.A1(_09706_),
    .A2(_09707_),
    .B1(_09681_),
    .B2(_09708_),
    .X(_09825_));
 sky130_fd_sc_hd__a2bb2o_1 _25736_ (.A1_N(_09824_),
    .A2_N(_09825_),
    .B1(_09824_),
    .B2(_09825_),
    .X(_09826_));
 sky130_fd_sc_hd__a2bb2o_1 _25737_ (.A1_N(_09776_),
    .A2_N(_09826_),
    .B1(_09776_),
    .B2(_09826_),
    .X(_09827_));
 sky130_fd_sc_hd__o22a_1 _25738_ (.A1(_09709_),
    .A2(_09710_),
    .B1(_09664_),
    .B2(_09711_),
    .X(_09828_));
 sky130_fd_sc_hd__a2bb2o_1 _25739_ (.A1_N(_09827_),
    .A2_N(_09828_),
    .B1(_09827_),
    .B2(_09828_),
    .X(_09829_));
 sky130_fd_sc_hd__a2bb2o_1 _25740_ (.A1_N(_09747_),
    .A2_N(_09829_),
    .B1(_09747_),
    .B2(_09829_),
    .X(_09830_));
 sky130_fd_sc_hd__o22a_1 _25741_ (.A1(_09712_),
    .A2(_09713_),
    .B1(_09635_),
    .B2(_09714_),
    .X(_09831_));
 sky130_fd_sc_hd__a2bb2o_1 _25742_ (.A1_N(_09830_),
    .A2_N(_09831_),
    .B1(_09830_),
    .B2(_09831_),
    .X(_09832_));
 sky130_fd_sc_hd__a2bb2o_1 _25743_ (.A1_N(_09730_),
    .A2_N(_09832_),
    .B1(_09730_),
    .B2(_09832_),
    .X(_09833_));
 sky130_fd_sc_hd__o22a_1 _25744_ (.A1(_09715_),
    .A2(_09716_),
    .B1(_09615_),
    .B2(_09717_),
    .X(_09834_));
 sky130_fd_sc_hd__a2bb2o_1 _25745_ (.A1_N(_09833_),
    .A2_N(_09834_),
    .B1(_09833_),
    .B2(_09834_),
    .X(_09835_));
 sky130_fd_sc_hd__a2bb2o_1 _25746_ (.A1_N(_09614_),
    .A2_N(_09835_),
    .B1(_09614_),
    .B2(_09835_),
    .X(_09836_));
 sky130_fd_sc_hd__and2_1 _25747_ (.A(_09727_),
    .B(_09836_),
    .X(_09837_));
 sky130_fd_sc_hd__or2_1 _25748_ (.A(_09727_),
    .B(_09836_),
    .X(_09838_));
 sky130_fd_sc_hd__or2b_1 _25749_ (.A(_09837_),
    .B_N(_09838_),
    .X(_09839_));
 sky130_fd_sc_hd__o21ai_1 _25750_ (.A1(_09724_),
    .A2(_09726_),
    .B1(_09723_),
    .Y(_09840_));
 sky130_fd_sc_hd__a2bb2o_1 _25751_ (.A1_N(_09839_),
    .A2_N(_09840_),
    .B1(_09839_),
    .B2(_09840_),
    .X(_02662_));
 sky130_fd_sc_hd__o22a_1 _25752_ (.A1(_09732_),
    .A2(_09745_),
    .B1(_09731_),
    .B2(_09746_),
    .X(_09841_));
 sky130_fd_sc_hd__or2_1 _25753_ (.A(_09353_),
    .B(_09841_),
    .X(_09842_));
 sky130_fd_sc_hd__a21bo_1 _25754_ (.A1(_09352_),
    .A2(_09841_),
    .B1_N(_09842_),
    .X(_09843_));
 sky130_fd_sc_hd__o22a_1 _25755_ (.A1(_09741_),
    .A2(_09742_),
    .B1(_09357_),
    .B2(_09744_),
    .X(_09844_));
 sky130_fd_sc_hd__o22a_1 _25756_ (.A1(_09749_),
    .A2(_09774_),
    .B1(_09748_),
    .B2(_09775_),
    .X(_09845_));
 sky130_fd_sc_hd__o22a_1 _25757_ (.A1(_09759_),
    .A2(_09760_),
    .B1(_09752_),
    .B2(_09761_),
    .X(_09846_));
 sky130_fd_sc_hd__o22a_2 _25758_ (.A1(_09639_),
    .A2(_09750_),
    .B1(_09517_),
    .B2(_09751_),
    .X(_09847_));
 sky130_fd_sc_hd__or2_1 _25759_ (.A(_09366_),
    .B(_09847_),
    .X(_09848_));
 sky130_fd_sc_hd__a21bo_1 _25760_ (.A1(_09366_),
    .A2(_09847_),
    .B1_N(_09848_),
    .X(_09849_));
 sky130_fd_sc_hd__a2bb2o_1 _25761_ (.A1_N(_09498_),
    .A2_N(_09849_),
    .B1(_09498_),
    .B2(_09849_),
    .X(_09850_));
 sky130_fd_sc_hd__buf_1 _25762_ (.A(_09850_),
    .X(_09851_));
 sky130_fd_sc_hd__o2bb2ai_1 _25763_ (.A1_N(_09846_),
    .A2_N(_09851_),
    .B1(_09846_),
    .B2(_09851_),
    .Y(_09852_));
 sky130_fd_sc_hd__o22a_1 _25764_ (.A1(_09495_),
    .A2(_09734_),
    .B1(_09626_),
    .B2(_09735_),
    .X(_09853_));
 sky130_fd_sc_hd__o2bb2a_1 _25765_ (.A1_N(_09852_),
    .A2_N(_09853_),
    .B1(_09852_),
    .B2(_09853_),
    .X(_09854_));
 sky130_vsdinv _25766_ (.A(_09854_),
    .Y(_09855_));
 sky130_fd_sc_hd__o22a_1 _25767_ (.A1(_09733_),
    .A2(_09736_),
    .B1(_09737_),
    .B2(_09739_),
    .X(_09856_));
 sky130_vsdinv _25768_ (.A(_09856_),
    .Y(_09857_));
 sky130_fd_sc_hd__a22o_1 _25769_ (.A1(_09855_),
    .A2(_09856_),
    .B1(_09854_),
    .B2(_09857_),
    .X(_09858_));
 sky130_fd_sc_hd__a2bb2o_1 _25770_ (.A1_N(_09375_),
    .A2_N(_09858_),
    .B1(_09375_),
    .B2(_09858_),
    .X(_09859_));
 sky130_fd_sc_hd__a2bb2o_1 _25771_ (.A1_N(_09845_),
    .A2_N(_09859_),
    .B1(_09845_),
    .B2(_09859_),
    .X(_09860_));
 sky130_fd_sc_hd__a2bb2o_1 _25772_ (.A1_N(_09844_),
    .A2_N(_09860_),
    .B1(_09844_),
    .B2(_09860_),
    .X(_09861_));
 sky130_fd_sc_hd__o22a_1 _25773_ (.A1(_09771_),
    .A2(_09772_),
    .B1(_09762_),
    .B2(_09773_),
    .X(_09862_));
 sky130_fd_sc_hd__o22a_2 _25774_ (.A1(_09778_),
    .A2(_09793_),
    .B1(_09777_),
    .B2(_09794_),
    .X(_09863_));
 sky130_fd_sc_hd__o22a_1 _25775_ (.A1(_06830_),
    .A2(_08837_),
    .B1(_05788_),
    .B2(_08033_),
    .X(_09864_));
 sky130_fd_sc_hd__and4_1 _25776_ (.A(_07115_),
    .B(_08667_),
    .C(_07116_),
    .D(_08668_),
    .X(_09865_));
 sky130_fd_sc_hd__nor2_4 _25777_ (.A(_09864_),
    .B(_09865_),
    .Y(_09866_));
 sky130_fd_sc_hd__clkbuf_2 _25778_ (.A(_08340_),
    .X(_09867_));
 sky130_fd_sc_hd__nor2_2 _25779_ (.A(_09867_),
    .B(_05708_),
    .Y(_09868_));
 sky130_fd_sc_hd__a2bb2o_1 _25780_ (.A1_N(_09866_),
    .A2_N(_09868_),
    .B1(_09866_),
    .B2(_09868_),
    .X(_09869_));
 sky130_fd_sc_hd__a31o_1 _25781_ (.A1(\pcpi_mul.rs2[12] ),
    .A2(_08820_),
    .A3(_09757_),
    .B1(_09756_),
    .X(_09870_));
 sky130_vsdinv _25782_ (.A(_09870_),
    .Y(_09871_));
 sky130_vsdinv _25783_ (.A(_09869_),
    .Y(_09872_));
 sky130_fd_sc_hd__a22o_1 _25784_ (.A1(_09869_),
    .A2(_09871_),
    .B1(_09872_),
    .B2(_09870_),
    .X(_09873_));
 sky130_fd_sc_hd__buf_1 _25785_ (.A(_09753_),
    .X(_09874_));
 sky130_fd_sc_hd__a2bb2o_1 _25786_ (.A1_N(_09754_),
    .A2_N(_09873_),
    .B1(_09874_),
    .B2(_09873_),
    .X(_09875_));
 sky130_fd_sc_hd__a21oi_2 _25787_ (.A1(_09767_),
    .A2(_09768_),
    .B1(_09766_),
    .Y(_09876_));
 sky130_fd_sc_hd__a21oi_4 _25788_ (.A1(_09781_),
    .A2(_09784_),
    .B1(_09780_),
    .Y(_09877_));
 sky130_fd_sc_hd__o22a_1 _25789_ (.A1(_09396_),
    .A2(_07463_),
    .B1(_09274_),
    .B2(_07595_),
    .X(_09878_));
 sky130_fd_sc_hd__and4_2 _25790_ (.A(_09398_),
    .B(_07587_),
    .C(_09399_),
    .D(_13519_),
    .X(_09879_));
 sky130_fd_sc_hd__nor2_2 _25791_ (.A(_09878_),
    .B(_09879_),
    .Y(_09880_));
 sky130_fd_sc_hd__nor2_2 _25792_ (.A(_09402_),
    .B(_07749_),
    .Y(_09881_));
 sky130_fd_sc_hd__a2bb2o_1 _25793_ (.A1_N(_09880_),
    .A2_N(_09881_),
    .B1(_09880_),
    .B2(_09881_),
    .X(_09882_));
 sky130_fd_sc_hd__a2bb2o_1 _25794_ (.A1_N(_09877_),
    .A2_N(_09882_),
    .B1(_09877_),
    .B2(_09882_),
    .X(_09883_));
 sky130_fd_sc_hd__a2bb2o_1 _25795_ (.A1_N(_09876_),
    .A2_N(_09883_),
    .B1(_09876_),
    .B2(_09883_),
    .X(_09884_));
 sky130_fd_sc_hd__o22a_1 _25796_ (.A1(_09764_),
    .A2(_09769_),
    .B1(_09763_),
    .B2(_09770_),
    .X(_09885_));
 sky130_fd_sc_hd__a2bb2o_1 _25797_ (.A1_N(_09884_),
    .A2_N(_09885_),
    .B1(_09884_),
    .B2(_09885_),
    .X(_09886_));
 sky130_fd_sc_hd__a2bb2o_1 _25798_ (.A1_N(_09875_),
    .A2_N(_09886_),
    .B1(_09875_),
    .B2(_09886_),
    .X(_09887_));
 sky130_fd_sc_hd__a2bb2o_1 _25799_ (.A1_N(_09863_),
    .A2_N(_09887_),
    .B1(_09863_),
    .B2(_09887_),
    .X(_09888_));
 sky130_fd_sc_hd__a2bb2o_1 _25800_ (.A1_N(_09862_),
    .A2_N(_09888_),
    .B1(_09862_),
    .B2(_09888_),
    .X(_09889_));
 sky130_fd_sc_hd__o22a_1 _25801_ (.A1(_09790_),
    .A2(_09791_),
    .B1(_09785_),
    .B2(_09792_),
    .X(_09890_));
 sky130_fd_sc_hd__o22a_1 _25802_ (.A1(_09797_),
    .A2(_09802_),
    .B1(_09796_),
    .B2(_09803_),
    .X(_09891_));
 sky130_fd_sc_hd__o22a_1 _25803_ (.A1(_08889_),
    .A2(_07172_),
    .B1(_08736_),
    .B2(_09782_),
    .X(_09892_));
 sky130_fd_sc_hd__and4_1 _25804_ (.A(_13106_),
    .B(_07598_),
    .C(_13112_),
    .D(_07886_),
    .X(_09893_));
 sky130_fd_sc_hd__nor2_2 _25805_ (.A(_09892_),
    .B(_09893_),
    .Y(_09894_));
 sky130_fd_sc_hd__clkbuf_2 _25806_ (.A(_07326_),
    .X(_09895_));
 sky130_fd_sc_hd__nor2_2 _25807_ (.A(_08734_),
    .B(_09895_),
    .Y(_09896_));
 sky130_fd_sc_hd__a2bb2o_2 _25808_ (.A1_N(_09894_),
    .A2_N(_09896_),
    .B1(_09894_),
    .B2(_09896_),
    .X(_09897_));
 sky130_fd_sc_hd__o22a_1 _25809_ (.A1(_08897_),
    .A2(_07762_),
    .B1(_09422_),
    .B2(_06762_),
    .X(_09898_));
 sky130_fd_sc_hd__and4_2 _25810_ (.A(_08745_),
    .B(_07191_),
    .C(_08746_),
    .D(_07764_),
    .X(_09899_));
 sky130_fd_sc_hd__nor2_2 _25811_ (.A(_09898_),
    .B(_09899_),
    .Y(_09900_));
 sky130_fd_sc_hd__nor2_4 _25812_ (.A(_08895_),
    .B(_06892_),
    .Y(_09901_));
 sky130_fd_sc_hd__a2bb2o_1 _25813_ (.A1_N(_09900_),
    .A2_N(_09901_),
    .B1(_09900_),
    .B2(_09901_),
    .X(_09902_));
 sky130_fd_sc_hd__a21oi_2 _25814_ (.A1(_09788_),
    .A2(_09789_),
    .B1(_09787_),
    .Y(_09903_));
 sky130_fd_sc_hd__a2bb2o_1 _25815_ (.A1_N(_09902_),
    .A2_N(_09903_),
    .B1(_09902_),
    .B2(_09903_),
    .X(_09904_));
 sky130_fd_sc_hd__a2bb2o_1 _25816_ (.A1_N(_09897_),
    .A2_N(_09904_),
    .B1(_09897_),
    .B2(_09904_),
    .X(_09905_));
 sky130_fd_sc_hd__a2bb2o_1 _25817_ (.A1_N(_09891_),
    .A2_N(_09905_),
    .B1(_09891_),
    .B2(_09905_),
    .X(_09906_));
 sky130_fd_sc_hd__a2bb2o_1 _25818_ (.A1_N(_09890_),
    .A2_N(_09906_),
    .B1(_09890_),
    .B2(_09906_),
    .X(_09907_));
 sky130_fd_sc_hd__a21oi_2 _25819_ (.A1(_09800_),
    .A2(_09801_),
    .B1(_09799_),
    .Y(_09908_));
 sky130_fd_sc_hd__a21oi_2 _25820_ (.A1(_09808_),
    .A2(_09809_),
    .B1(_09807_),
    .Y(_09909_));
 sky130_fd_sc_hd__o22a_1 _25821_ (.A1(_09436_),
    .A2(_06766_),
    .B1(_07268_),
    .B2(_07036_),
    .X(_09910_));
 sky130_fd_sc_hd__buf_1 _25822_ (.A(_08124_),
    .X(_09911_));
 sky130_fd_sc_hd__and4_1 _25823_ (.A(_13088_),
    .B(_06899_),
    .C(_09911_),
    .D(_06901_),
    .X(_09912_));
 sky130_fd_sc_hd__nor2_2 _25824_ (.A(_09910_),
    .B(_09912_),
    .Y(_09913_));
 sky130_fd_sc_hd__nor2_2 _25825_ (.A(_07074_),
    .B(_06576_),
    .Y(_09914_));
 sky130_fd_sc_hd__a2bb2o_1 _25826_ (.A1_N(_09913_),
    .A2_N(_09914_),
    .B1(_09913_),
    .B2(_09914_),
    .X(_09915_));
 sky130_fd_sc_hd__a2bb2o_1 _25827_ (.A1_N(_09909_),
    .A2_N(_09915_),
    .B1(_09909_),
    .B2(_09915_),
    .X(_09916_));
 sky130_fd_sc_hd__a2bb2o_1 _25828_ (.A1_N(_09908_),
    .A2_N(_09916_),
    .B1(_09908_),
    .B2(_09916_),
    .X(_09917_));
 sky130_fd_sc_hd__clkbuf_4 _25829_ (.A(_08286_),
    .X(_09918_));
 sky130_fd_sc_hd__clkbuf_4 _25830_ (.A(_08287_),
    .X(_09919_));
 sky130_fd_sc_hd__o22a_1 _25831_ (.A1(_09918_),
    .A2(_06669_),
    .B1(_09919_),
    .B2(_06327_),
    .X(_09920_));
 sky130_fd_sc_hd__and4_1 _25832_ (.A(_13074_),
    .B(_13571_),
    .C(_09806_),
    .D(_06584_),
    .X(_09921_));
 sky130_fd_sc_hd__nor2_2 _25833_ (.A(_09920_),
    .B(_09921_),
    .Y(_09922_));
 sky130_fd_sc_hd__nor2_2 _25834_ (.A(_07682_),
    .B(_06435_),
    .Y(_09923_));
 sky130_fd_sc_hd__a2bb2o_1 _25835_ (.A1_N(_09922_),
    .A2_N(_09923_),
    .B1(_09922_),
    .B2(_09923_),
    .X(_09924_));
 sky130_fd_sc_hd__or2_1 _25836_ (.A(_08772_),
    .B(_08417_),
    .X(_09925_));
 sky130_fd_sc_hd__and4_1 _25837_ (.A(_09190_),
    .B(_05926_),
    .C(_08775_),
    .D(_07371_),
    .X(_09926_));
 sky130_fd_sc_hd__o22a_1 _25838_ (.A1(_08777_),
    .A2(_06145_),
    .B1(_08778_),
    .B2(_05836_),
    .X(_09927_));
 sky130_fd_sc_hd__or2_1 _25839_ (.A(_09926_),
    .B(_09927_),
    .X(_09928_));
 sky130_fd_sc_hd__a2bb2o_1 _25840_ (.A1_N(_09925_),
    .A2_N(_09928_),
    .B1(_09925_),
    .B2(_09928_),
    .X(_09929_));
 sky130_fd_sc_hd__o21ba_1 _25841_ (.A1(_09811_),
    .A2(_09814_),
    .B1_N(_09812_),
    .X(_09930_));
 sky130_fd_sc_hd__a2bb2o_1 _25842_ (.A1_N(_09929_),
    .A2_N(_09930_),
    .B1(_09929_),
    .B2(_09930_),
    .X(_09931_));
 sky130_fd_sc_hd__a2bb2o_1 _25843_ (.A1_N(_09924_),
    .A2_N(_09931_),
    .B1(_09924_),
    .B2(_09931_),
    .X(_09932_));
 sky130_fd_sc_hd__o22a_1 _25844_ (.A1(_09815_),
    .A2(_09816_),
    .B1(_09810_),
    .B2(_09817_),
    .X(_09933_));
 sky130_fd_sc_hd__a2bb2o_1 _25845_ (.A1_N(_09932_),
    .A2_N(_09933_),
    .B1(_09932_),
    .B2(_09933_),
    .X(_09934_));
 sky130_fd_sc_hd__a2bb2o_1 _25846_ (.A1_N(_09917_),
    .A2_N(_09934_),
    .B1(_09917_),
    .B2(_09934_),
    .X(_09935_));
 sky130_fd_sc_hd__o22a_1 _25847_ (.A1(_09818_),
    .A2(_09819_),
    .B1(_09804_),
    .B2(_09820_),
    .X(_09936_));
 sky130_fd_sc_hd__a2bb2o_1 _25848_ (.A1_N(_09935_),
    .A2_N(_09936_),
    .B1(_09935_),
    .B2(_09936_),
    .X(_09937_));
 sky130_fd_sc_hd__a2bb2o_2 _25849_ (.A1_N(_09907_),
    .A2_N(_09937_),
    .B1(_09907_),
    .B2(_09937_),
    .X(_09938_));
 sky130_fd_sc_hd__o22a_2 _25850_ (.A1(_09821_),
    .A2(_09822_),
    .B1(_09795_),
    .B2(_09823_),
    .X(_09939_));
 sky130_fd_sc_hd__a2bb2o_1 _25851_ (.A1_N(_09938_),
    .A2_N(_09939_),
    .B1(_09938_),
    .B2(_09939_),
    .X(_09940_));
 sky130_fd_sc_hd__a2bb2o_1 _25852_ (.A1_N(_09889_),
    .A2_N(_09940_),
    .B1(_09889_),
    .B2(_09940_),
    .X(_09941_));
 sky130_fd_sc_hd__o22a_1 _25853_ (.A1(_09824_),
    .A2(_09825_),
    .B1(_09776_),
    .B2(_09826_),
    .X(_09942_));
 sky130_fd_sc_hd__a2bb2o_1 _25854_ (.A1_N(_09941_),
    .A2_N(_09942_),
    .B1(_09941_),
    .B2(_09942_),
    .X(_09943_));
 sky130_fd_sc_hd__a2bb2o_1 _25855_ (.A1_N(_09861_),
    .A2_N(_09943_),
    .B1(_09861_),
    .B2(_09943_),
    .X(_09944_));
 sky130_fd_sc_hd__o22a_1 _25856_ (.A1(_09827_),
    .A2(_09828_),
    .B1(_09747_),
    .B2(_09829_),
    .X(_09945_));
 sky130_fd_sc_hd__a2bb2o_1 _25857_ (.A1_N(_09944_),
    .A2_N(_09945_),
    .B1(_09944_),
    .B2(_09945_),
    .X(_09946_));
 sky130_fd_sc_hd__a2bb2o_1 _25858_ (.A1_N(_09843_),
    .A2_N(_09946_),
    .B1(_09843_),
    .B2(_09946_),
    .X(_09947_));
 sky130_fd_sc_hd__o22a_1 _25859_ (.A1(_09830_),
    .A2(_09831_),
    .B1(_09730_),
    .B2(_09832_),
    .X(_09948_));
 sky130_fd_sc_hd__a2bb2o_1 _25860_ (.A1_N(_09947_),
    .A2_N(_09948_),
    .B1(_09947_),
    .B2(_09948_),
    .X(_09949_));
 sky130_fd_sc_hd__a2bb2o_1 _25861_ (.A1_N(_09729_),
    .A2_N(_09949_),
    .B1(_09729_),
    .B2(_09949_),
    .X(_09950_));
 sky130_fd_sc_hd__o22a_1 _25862_ (.A1(_09833_),
    .A2(_09834_),
    .B1(_09614_),
    .B2(_09835_),
    .X(_09951_));
 sky130_fd_sc_hd__or2_1 _25863_ (.A(_09950_),
    .B(_09951_),
    .X(_09952_));
 sky130_fd_sc_hd__a21bo_1 _25864_ (.A1(_09950_),
    .A2(_09951_),
    .B1_N(_09952_),
    .X(_09953_));
 sky130_fd_sc_hd__buf_1 _25865_ (.A(_09953_),
    .X(_09954_));
 sky130_fd_sc_hd__or2_1 _25866_ (.A(_09724_),
    .B(_09839_),
    .X(_09955_));
 sky130_fd_sc_hd__or3_1 _25867_ (.A(_09477_),
    .B(_09610_),
    .C(_09955_),
    .X(_09956_));
 sky130_fd_sc_hd__o221a_1 _25868_ (.A1(_09723_),
    .A2(_09837_),
    .B1(_09725_),
    .B2(_09955_),
    .C1(_09838_),
    .X(_09957_));
 sky130_fd_sc_hd__o21ai_2 _25869_ (.A1(_09486_),
    .A2(_09956_),
    .B1(_09957_),
    .Y(_09958_));
 sky130_vsdinv _25870_ (.A(_09958_),
    .Y(_09959_));
 sky130_vsdinv _25871_ (.A(_09954_),
    .Y(_09960_));
 sky130_fd_sc_hd__o22a_1 _25872_ (.A1(_09954_),
    .A2(_09959_),
    .B1(_09960_),
    .B2(_09958_),
    .X(_02663_));
 sky130_fd_sc_hd__o22a_1 _25873_ (.A1(_09947_),
    .A2(_09948_),
    .B1(_09729_),
    .B2(_09949_),
    .X(_09961_));
 sky130_fd_sc_hd__o22a_1 _25874_ (.A1(_09845_),
    .A2(_09859_),
    .B1(_09844_),
    .B2(_09860_),
    .X(_09962_));
 sky130_fd_sc_hd__or2_1 _25875_ (.A(_09613_),
    .B(_09962_),
    .X(_09963_));
 sky130_fd_sc_hd__a21bo_1 _25876_ (.A1(_09489_),
    .A2(_09962_),
    .B1_N(_09963_),
    .X(_09964_));
 sky130_fd_sc_hd__o22a_1 _25877_ (.A1(_09855_),
    .A2(_09856_),
    .B1(_09616_),
    .B2(_09858_),
    .X(_09965_));
 sky130_fd_sc_hd__o22a_1 _25878_ (.A1(_09863_),
    .A2(_09887_),
    .B1(_09862_),
    .B2(_09888_),
    .X(_09966_));
 sky130_fd_sc_hd__o22a_1 _25879_ (.A1(_09869_),
    .A2(_09871_),
    .B1(_09752_),
    .B2(_09873_),
    .X(_09967_));
 sky130_fd_sc_hd__a2bb2o_1 _25880_ (.A1_N(_09851_),
    .A2_N(_09967_),
    .B1(_09850_),
    .B2(_09967_),
    .X(_09968_));
 sky130_fd_sc_hd__buf_1 _25881_ (.A(_09848_),
    .X(_09969_));
 sky130_fd_sc_hd__o21a_1 _25882_ (.A1(_09626_),
    .A2(_09849_),
    .B1(_09969_),
    .X(_09970_));
 sky130_fd_sc_hd__o2bb2a_1 _25883_ (.A1_N(_09968_),
    .A2_N(_09970_),
    .B1(_09968_),
    .B2(_09970_),
    .X(_09971_));
 sky130_vsdinv _25884_ (.A(_09971_),
    .Y(_09972_));
 sky130_fd_sc_hd__buf_1 _25885_ (.A(_09850_),
    .X(_09973_));
 sky130_fd_sc_hd__o22a_1 _25886_ (.A1(_09846_),
    .A2(_09973_),
    .B1(_09852_),
    .B2(_09853_),
    .X(_09974_));
 sky130_vsdinv _25887_ (.A(_09974_),
    .Y(_09975_));
 sky130_fd_sc_hd__a22o_1 _25888_ (.A1(_09972_),
    .A2(_09974_),
    .B1(_09971_),
    .B2(_09975_),
    .X(_09976_));
 sky130_fd_sc_hd__a2bb2o_1 _25889_ (.A1_N(_09507_),
    .A2_N(_09976_),
    .B1(_09507_),
    .B2(_09976_),
    .X(_09977_));
 sky130_fd_sc_hd__a2bb2o_1 _25890_ (.A1_N(_09966_),
    .A2_N(_09977_),
    .B1(_09966_),
    .B2(_09977_),
    .X(_09978_));
 sky130_fd_sc_hd__a2bb2o_1 _25891_ (.A1_N(_09965_),
    .A2_N(_09978_),
    .B1(_09965_),
    .B2(_09978_),
    .X(_09979_));
 sky130_fd_sc_hd__o22a_1 _25892_ (.A1(_09884_),
    .A2(_09885_),
    .B1(_09875_),
    .B2(_09886_),
    .X(_09980_));
 sky130_fd_sc_hd__o22a_2 _25893_ (.A1(_09891_),
    .A2(_09905_),
    .B1(_09890_),
    .B2(_09906_),
    .X(_09981_));
 sky130_fd_sc_hd__a31o_1 _25894_ (.A1(_08974_),
    .A2(\pcpi_mul.rs2[12] ),
    .A3(_09866_),
    .B1(_09865_),
    .X(_09982_));
 sky130_vsdinv _25895_ (.A(_09982_),
    .Y(_09983_));
 sky130_fd_sc_hd__buf_1 _25896_ (.A(_09868_),
    .X(_09984_));
 sky130_fd_sc_hd__o22a_1 _25897_ (.A1(_09011_),
    .A2(_08497_),
    .B1(_09867_),
    .B2(_05789_),
    .X(_09985_));
 sky130_fd_sc_hd__and4_1 _25898_ (.A(_13130_),
    .B(_13505_),
    .C(_08814_),
    .D(_13133_),
    .X(_09986_));
 sky130_fd_sc_hd__nor2_1 _25899_ (.A(_09985_),
    .B(_09986_),
    .Y(_09987_));
 sky130_fd_sc_hd__o2bb2a_1 _25900_ (.A1_N(_09984_),
    .A2_N(_09987_),
    .B1(_09984_),
    .B2(_09987_),
    .X(_09988_));
 sky130_vsdinv _25901_ (.A(_09988_),
    .Y(_09989_));
 sky130_fd_sc_hd__a22o_1 _25902_ (.A1(_09983_),
    .A2(_09989_),
    .B1(_09982_),
    .B2(_09988_),
    .X(_09990_));
 sky130_fd_sc_hd__a2bb2o_1 _25903_ (.A1_N(_09874_),
    .A2_N(_09990_),
    .B1(_09874_),
    .B2(_09990_),
    .X(_09991_));
 sky130_fd_sc_hd__a21oi_2 _25904_ (.A1(_09880_),
    .A2(_09881_),
    .B1(_09879_),
    .Y(_09992_));
 sky130_fd_sc_hd__a21oi_2 _25905_ (.A1(_09894_),
    .A2(_09896_),
    .B1(_09893_),
    .Y(_09993_));
 sky130_fd_sc_hd__o22a_1 _25906_ (.A1(_08233_),
    .A2(_07595_),
    .B1(_06094_),
    .B2(_07748_),
    .X(_09994_));
 sky130_fd_sc_hd__and4_2 _25907_ (.A(_08236_),
    .B(_13519_),
    .C(_08238_),
    .D(_13515_),
    .X(_09995_));
 sky130_fd_sc_hd__nor2_2 _25908_ (.A(_09994_),
    .B(_09995_),
    .Y(_09996_));
 sky130_fd_sc_hd__nor2_2 _25909_ (.A(_09402_),
    .B(_08839_),
    .Y(_09997_));
 sky130_fd_sc_hd__a2bb2o_1 _25910_ (.A1_N(_09996_),
    .A2_N(_09997_),
    .B1(_09996_),
    .B2(_09997_),
    .X(_09998_));
 sky130_fd_sc_hd__a2bb2o_1 _25911_ (.A1_N(_09993_),
    .A2_N(_09998_),
    .B1(_09993_),
    .B2(_09998_),
    .X(_09999_));
 sky130_fd_sc_hd__a2bb2o_1 _25912_ (.A1_N(_09992_),
    .A2_N(_09999_),
    .B1(_09992_),
    .B2(_09999_),
    .X(_10000_));
 sky130_fd_sc_hd__o22a_1 _25913_ (.A1(_09877_),
    .A2(_09882_),
    .B1(_09876_),
    .B2(_09883_),
    .X(_10001_));
 sky130_fd_sc_hd__a2bb2o_1 _25914_ (.A1_N(_10000_),
    .A2_N(_10001_),
    .B1(_10000_),
    .B2(_10001_),
    .X(_10002_));
 sky130_fd_sc_hd__a2bb2o_1 _25915_ (.A1_N(_09991_),
    .A2_N(_10002_),
    .B1(_09991_),
    .B2(_10002_),
    .X(_10003_));
 sky130_fd_sc_hd__a2bb2o_1 _25916_ (.A1_N(_09981_),
    .A2_N(_10003_),
    .B1(_09981_),
    .B2(_10003_),
    .X(_10004_));
 sky130_fd_sc_hd__a2bb2o_1 _25917_ (.A1_N(_09980_),
    .A2_N(_10004_),
    .B1(_09980_),
    .B2(_10004_),
    .X(_10005_));
 sky130_fd_sc_hd__o22a_2 _25918_ (.A1(_09902_),
    .A2(_09903_),
    .B1(_09897_),
    .B2(_09904_),
    .X(_10006_));
 sky130_fd_sc_hd__o22a_2 _25919_ (.A1(_09909_),
    .A2(_09915_),
    .B1(_09908_),
    .B2(_09916_),
    .X(_10007_));
 sky130_fd_sc_hd__buf_2 _25920_ (.A(_08574_),
    .X(_10008_));
 sky130_fd_sc_hd__o22a_1 _25921_ (.A1(_10008_),
    .A2(_09782_),
    .B1(_06391_),
    .B2(_07884_),
    .X(_10009_));
 sky130_fd_sc_hd__and4_1 _25922_ (.A(_13107_),
    .B(_07886_),
    .C(_13113_),
    .D(_07449_),
    .X(_10010_));
 sky130_fd_sc_hd__nor2_2 _25923_ (.A(_10009_),
    .B(_10010_),
    .Y(_10011_));
 sky130_fd_sc_hd__clkbuf_2 _25924_ (.A(_08178_),
    .X(_10012_));
 sky130_fd_sc_hd__nor2_2 _25925_ (.A(_06286_),
    .B(_10012_),
    .Y(_10013_));
 sky130_fd_sc_hd__a2bb2o_1 _25926_ (.A1_N(_10011_),
    .A2_N(_10013_),
    .B1(_10011_),
    .B2(_10013_),
    .X(_10014_));
 sky130_fd_sc_hd__o22a_1 _25927_ (.A1(_09552_),
    .A2(_07332_),
    .B1(_06802_),
    .B2(_07468_),
    .X(_10015_));
 sky130_fd_sc_hd__and4_2 _25928_ (.A(_13098_),
    .B(_07330_),
    .C(_13103_),
    .D(_08053_),
    .X(_10016_));
 sky130_fd_sc_hd__nor2_2 _25929_ (.A(_10015_),
    .B(_10016_),
    .Y(_10017_));
 sky130_fd_sc_hd__nor2_4 _25930_ (.A(_09558_),
    .B(_07034_),
    .Y(_10018_));
 sky130_fd_sc_hd__a2bb2o_2 _25931_ (.A1_N(_10017_),
    .A2_N(_10018_),
    .B1(_10017_),
    .B2(_10018_),
    .X(_10019_));
 sky130_fd_sc_hd__a21oi_4 _25932_ (.A1(_09900_),
    .A2(_09901_),
    .B1(_09899_),
    .Y(_10020_));
 sky130_fd_sc_hd__a2bb2o_1 _25933_ (.A1_N(_10019_),
    .A2_N(_10020_),
    .B1(_10019_),
    .B2(_10020_),
    .X(_10021_));
 sky130_fd_sc_hd__a2bb2o_1 _25934_ (.A1_N(_10014_),
    .A2_N(_10021_),
    .B1(_10014_),
    .B2(_10021_),
    .X(_10022_));
 sky130_fd_sc_hd__a2bb2o_1 _25935_ (.A1_N(_10007_),
    .A2_N(_10022_),
    .B1(_10007_),
    .B2(_10022_),
    .X(_10023_));
 sky130_fd_sc_hd__a2bb2o_1 _25936_ (.A1_N(_10006_),
    .A2_N(_10023_),
    .B1(_10006_),
    .B2(_10023_),
    .X(_10024_));
 sky130_fd_sc_hd__a21oi_2 _25937_ (.A1(_09913_),
    .A2(_09914_),
    .B1(_09912_),
    .Y(_10025_));
 sky130_fd_sc_hd__a21oi_2 _25938_ (.A1(_09922_),
    .A2(_09923_),
    .B1(_09921_),
    .Y(_10026_));
 sky130_fd_sc_hd__o22a_1 _25939_ (.A1(_09436_),
    .A2(_06451_),
    .B1(_07268_),
    .B2(_07037_),
    .X(_10027_));
 sky130_fd_sc_hd__clkbuf_2 _25940_ (.A(_08123_),
    .X(_10028_));
 sky130_fd_sc_hd__and4_1 _25941_ (.A(_10028_),
    .B(_13556_),
    .C(_09911_),
    .D(_07040_),
    .X(_10029_));
 sky130_fd_sc_hd__nor2_2 _25942_ (.A(_10027_),
    .B(_10029_),
    .Y(_10030_));
 sky130_fd_sc_hd__clkbuf_4 _25943_ (.A(_07073_),
    .X(_10031_));
 sky130_fd_sc_hd__nor2_2 _25944_ (.A(_10031_),
    .B(_06755_),
    .Y(_10032_));
 sky130_fd_sc_hd__a2bb2o_1 _25945_ (.A1_N(_10030_),
    .A2_N(_10032_),
    .B1(_10030_),
    .B2(_10032_),
    .X(_10033_));
 sky130_fd_sc_hd__a2bb2o_1 _25946_ (.A1_N(_10026_),
    .A2_N(_10033_),
    .B1(_10026_),
    .B2(_10033_),
    .X(_10034_));
 sky130_fd_sc_hd__a2bb2o_1 _25947_ (.A1_N(_10025_),
    .A2_N(_10034_),
    .B1(_10025_),
    .B2(_10034_),
    .X(_10035_));
 sky130_fd_sc_hd__o22a_1 _25948_ (.A1(_09575_),
    .A2(_06783_),
    .B1(_09919_),
    .B2(_06917_),
    .X(_10036_));
 sky130_fd_sc_hd__and4_1 _25949_ (.A(_13074_),
    .B(_06584_),
    .C(_09806_),
    .D(_06768_),
    .X(_10037_));
 sky130_fd_sc_hd__nor2_2 _25950_ (.A(_10036_),
    .B(_10037_),
    .Y(_10038_));
 sky130_fd_sc_hd__nor2_2 _25951_ (.A(_07682_),
    .B(_08887_),
    .Y(_10039_));
 sky130_fd_sc_hd__a2bb2o_1 _25952_ (.A1_N(_10038_),
    .A2_N(_10039_),
    .B1(_10038_),
    .B2(_10039_),
    .X(_10040_));
 sky130_fd_sc_hd__or2_1 _25953_ (.A(_08772_),
    .B(_06040_),
    .X(_10041_));
 sky130_fd_sc_hd__and4_1 _25954_ (.A(_08774_),
    .B(_05930_),
    .C(_08775_),
    .D(_13574_),
    .X(_10042_));
 sky130_fd_sc_hd__o22a_1 _25955_ (.A1(_08925_),
    .A2(_07371_),
    .B1(_08926_),
    .B2(_05943_),
    .X(_10043_));
 sky130_fd_sc_hd__or2_1 _25956_ (.A(_10042_),
    .B(_10043_),
    .X(_10044_));
 sky130_fd_sc_hd__a2bb2o_1 _25957_ (.A1_N(_10041_),
    .A2_N(_10044_),
    .B1(_10041_),
    .B2(_10044_),
    .X(_10045_));
 sky130_fd_sc_hd__o21ba_1 _25958_ (.A1(_09925_),
    .A2(_09928_),
    .B1_N(_09926_),
    .X(_10046_));
 sky130_fd_sc_hd__a2bb2o_1 _25959_ (.A1_N(_10045_),
    .A2_N(_10046_),
    .B1(_10045_),
    .B2(_10046_),
    .X(_10047_));
 sky130_fd_sc_hd__a2bb2o_1 _25960_ (.A1_N(_10040_),
    .A2_N(_10047_),
    .B1(_10040_),
    .B2(_10047_),
    .X(_10048_));
 sky130_fd_sc_hd__o22a_1 _25961_ (.A1(_09929_),
    .A2(_09930_),
    .B1(_09924_),
    .B2(_09931_),
    .X(_10049_));
 sky130_fd_sc_hd__a2bb2o_1 _25962_ (.A1_N(_10048_),
    .A2_N(_10049_),
    .B1(_10048_),
    .B2(_10049_),
    .X(_10050_));
 sky130_fd_sc_hd__a2bb2o_2 _25963_ (.A1_N(_10035_),
    .A2_N(_10050_),
    .B1(_10035_),
    .B2(_10050_),
    .X(_10051_));
 sky130_fd_sc_hd__o22a_2 _25964_ (.A1(_09932_),
    .A2(_09933_),
    .B1(_09917_),
    .B2(_09934_),
    .X(_10052_));
 sky130_fd_sc_hd__a2bb2o_1 _25965_ (.A1_N(_10051_),
    .A2_N(_10052_),
    .B1(_10051_),
    .B2(_10052_),
    .X(_10053_));
 sky130_fd_sc_hd__a2bb2o_1 _25966_ (.A1_N(_10024_),
    .A2_N(_10053_),
    .B1(_10024_),
    .B2(_10053_),
    .X(_10054_));
 sky130_fd_sc_hd__o22a_2 _25967_ (.A1(_09935_),
    .A2(_09936_),
    .B1(_09907_),
    .B2(_09937_),
    .X(_10055_));
 sky130_fd_sc_hd__a2bb2o_1 _25968_ (.A1_N(_10054_),
    .A2_N(_10055_),
    .B1(_10054_),
    .B2(_10055_),
    .X(_10056_));
 sky130_fd_sc_hd__a2bb2o_1 _25969_ (.A1_N(_10005_),
    .A2_N(_10056_),
    .B1(_10005_),
    .B2(_10056_),
    .X(_10057_));
 sky130_fd_sc_hd__o22a_1 _25970_ (.A1(_09938_),
    .A2(_09939_),
    .B1(_09889_),
    .B2(_09940_),
    .X(_10058_));
 sky130_fd_sc_hd__a2bb2o_1 _25971_ (.A1_N(_10057_),
    .A2_N(_10058_),
    .B1(_10057_),
    .B2(_10058_),
    .X(_10059_));
 sky130_fd_sc_hd__a2bb2o_1 _25972_ (.A1_N(_09979_),
    .A2_N(_10059_),
    .B1(_09979_),
    .B2(_10059_),
    .X(_10060_));
 sky130_fd_sc_hd__o22a_1 _25973_ (.A1(_09941_),
    .A2(_09942_),
    .B1(_09861_),
    .B2(_09943_),
    .X(_10061_));
 sky130_fd_sc_hd__a2bb2o_1 _25974_ (.A1_N(_10060_),
    .A2_N(_10061_),
    .B1(_10060_),
    .B2(_10061_),
    .X(_10062_));
 sky130_fd_sc_hd__a2bb2o_1 _25975_ (.A1_N(_09964_),
    .A2_N(_10062_),
    .B1(_09964_),
    .B2(_10062_),
    .X(_10063_));
 sky130_fd_sc_hd__o22a_1 _25976_ (.A1(_09944_),
    .A2(_09945_),
    .B1(_09843_),
    .B2(_09946_),
    .X(_10064_));
 sky130_fd_sc_hd__a2bb2o_1 _25977_ (.A1_N(_10063_),
    .A2_N(_10064_),
    .B1(_10063_),
    .B2(_10064_),
    .X(_10065_));
 sky130_fd_sc_hd__a2bb2o_1 _25978_ (.A1_N(_09842_),
    .A2_N(_10065_),
    .B1(_09842_),
    .B2(_10065_),
    .X(_10066_));
 sky130_fd_sc_hd__or2_1 _25979_ (.A(_09961_),
    .B(_10066_),
    .X(_10067_));
 sky130_fd_sc_hd__a21bo_1 _25980_ (.A1(_09961_),
    .A2(_10066_),
    .B1_N(_10067_),
    .X(_10068_));
 sky130_fd_sc_hd__o21ai_1 _25981_ (.A1(_09954_),
    .A2(_09959_),
    .B1(_09952_),
    .Y(_10069_));
 sky130_fd_sc_hd__a2bb2o_1 _25982_ (.A1_N(_10068_),
    .A2_N(_10069_),
    .B1(_10068_),
    .B2(_10069_),
    .X(_02664_));
 sky130_fd_sc_hd__o22a_1 _25983_ (.A1(_09966_),
    .A2(_09977_),
    .B1(_09965_),
    .B2(_09978_),
    .X(_10070_));
 sky130_fd_sc_hd__or2_1 _25984_ (.A(_09613_),
    .B(_10070_),
    .X(_10071_));
 sky130_fd_sc_hd__a21bo_1 _25985_ (.A1(_09351_),
    .A2(_10070_),
    .B1_N(_10071_),
    .X(_10072_));
 sky130_fd_sc_hd__o22a_1 _25986_ (.A1(_09972_),
    .A2(_09974_),
    .B1(_09616_),
    .B2(_09976_),
    .X(_10073_));
 sky130_fd_sc_hd__o22a_1 _25987_ (.A1(_09981_),
    .A2(_10003_),
    .B1(_09980_),
    .B2(_10004_),
    .X(_10074_));
 sky130_fd_sc_hd__buf_1 _25988_ (.A(_09970_),
    .X(_10075_));
 sky130_fd_sc_hd__o22a_1 _25989_ (.A1(_09983_),
    .A2(_09989_),
    .B1(_09753_),
    .B2(_09990_),
    .X(_10076_));
 sky130_fd_sc_hd__a2bb2o_1 _25990_ (.A1_N(_09973_),
    .A2_N(_10076_),
    .B1(_09851_),
    .B2(_10076_),
    .X(_10077_));
 sky130_fd_sc_hd__a2bb2o_1 _25991_ (.A1_N(_10075_),
    .A2_N(_10077_),
    .B1(_10075_),
    .B2(_10077_),
    .X(_10078_));
 sky130_fd_sc_hd__o22a_1 _25992_ (.A1(_09973_),
    .A2(_09967_),
    .B1(_09968_),
    .B2(_10075_),
    .X(_10079_));
 sky130_fd_sc_hd__o2bb2ai_1 _25993_ (.A1_N(_10078_),
    .A2_N(_10079_),
    .B1(_10078_),
    .B2(_10079_),
    .Y(_10080_));
 sky130_fd_sc_hd__a2bb2o_1 _25994_ (.A1_N(_09356_),
    .A2_N(_10080_),
    .B1(_09356_),
    .B2(_10080_),
    .X(_10081_));
 sky130_fd_sc_hd__a2bb2o_1 _25995_ (.A1_N(_10074_),
    .A2_N(_10081_),
    .B1(_10074_),
    .B2(_10081_),
    .X(_10082_));
 sky130_fd_sc_hd__a2bb2o_1 _25996_ (.A1_N(_10073_),
    .A2_N(_10082_),
    .B1(_10073_),
    .B2(_10082_),
    .X(_10083_));
 sky130_fd_sc_hd__o22a_1 _25997_ (.A1(_10000_),
    .A2(_10001_),
    .B1(_09991_),
    .B2(_10002_),
    .X(_10084_));
 sky130_fd_sc_hd__o22a_1 _25998_ (.A1(_10007_),
    .A2(_10022_),
    .B1(_10006_),
    .B2(_10023_),
    .X(_10085_));
 sky130_fd_sc_hd__clkbuf_2 _25999_ (.A(_09753_),
    .X(_10086_));
 sky130_fd_sc_hd__or4_4 _26000_ (.A(_11705_),
    .B(_05789_),
    .C(_11704_),
    .D(_09011_),
    .X(_10087_));
 sky130_fd_sc_hd__buf_1 _26001_ (.A(_08974_),
    .X(_10088_));
 sky130_fd_sc_hd__a22o_1 _26002_ (.A1(_10088_),
    .A2(_13133_),
    .B1(_10088_),
    .B2(_13130_),
    .X(_10089_));
 sky130_fd_sc_hd__nand2_2 _26003_ (.A(_10087_),
    .B(_10089_),
    .Y(_10090_));
 sky130_fd_sc_hd__clkbuf_2 _26004_ (.A(_05709_),
    .X(_10091_));
 sky130_fd_sc_hd__o22a_2 _26005_ (.A1(_09984_),
    .A2(_09986_),
    .B1(_10091_),
    .B2(_09985_),
    .X(_10092_));
 sky130_fd_sc_hd__a2bb2oi_4 _26006_ (.A1_N(_10090_),
    .A2_N(_10092_),
    .B1(_10090_),
    .B2(_10092_),
    .Y(_10093_));
 sky130_fd_sc_hd__a2bb2o_1 _26007_ (.A1_N(_10086_),
    .A2_N(_10093_),
    .B1(_10086_),
    .B2(_10093_),
    .X(_10094_));
 sky130_fd_sc_hd__a21oi_2 _26008_ (.A1(_09996_),
    .A2(_09997_),
    .B1(_09995_),
    .Y(_10095_));
 sky130_fd_sc_hd__a21oi_2 _26009_ (.A1(_10011_),
    .A2(_10013_),
    .B1(_10010_),
    .Y(_10096_));
 sky130_fd_sc_hd__o22a_1 _26010_ (.A1(_09021_),
    .A2(_07873_),
    .B1(_06090_),
    .B2(_08838_),
    .X(_10097_));
 sky130_fd_sc_hd__and4_1 _26011_ (.A(_13119_),
    .B(_08023_),
    .C(_13123_),
    .D(_13510_),
    .X(_10098_));
 sky130_fd_sc_hd__nor2_2 _26012_ (.A(_10097_),
    .B(_10098_),
    .Y(_10099_));
 sky130_fd_sc_hd__nor2_2 _26013_ (.A(_06000_),
    .B(_08036_),
    .Y(_10100_));
 sky130_fd_sc_hd__a2bb2o_1 _26014_ (.A1_N(_10099_),
    .A2_N(_10100_),
    .B1(_10099_),
    .B2(_10100_),
    .X(_10101_));
 sky130_fd_sc_hd__a2bb2o_1 _26015_ (.A1_N(_10096_),
    .A2_N(_10101_),
    .B1(_10096_),
    .B2(_10101_),
    .X(_10102_));
 sky130_fd_sc_hd__a2bb2o_1 _26016_ (.A1_N(_10095_),
    .A2_N(_10102_),
    .B1(_10095_),
    .B2(_10102_),
    .X(_10103_));
 sky130_fd_sc_hd__o22a_1 _26017_ (.A1(_09993_),
    .A2(_09998_),
    .B1(_09992_),
    .B2(_09999_),
    .X(_10104_));
 sky130_fd_sc_hd__a2bb2o_1 _26018_ (.A1_N(_10103_),
    .A2_N(_10104_),
    .B1(_10103_),
    .B2(_10104_),
    .X(_10105_));
 sky130_fd_sc_hd__a2bb2o_1 _26019_ (.A1_N(_10094_),
    .A2_N(_10105_),
    .B1(_10094_),
    .B2(_10105_),
    .X(_10106_));
 sky130_fd_sc_hd__a2bb2o_1 _26020_ (.A1_N(_10085_),
    .A2_N(_10106_),
    .B1(_10085_),
    .B2(_10106_),
    .X(_10107_));
 sky130_fd_sc_hd__a2bb2o_1 _26021_ (.A1_N(_10084_),
    .A2_N(_10107_),
    .B1(_10084_),
    .B2(_10107_),
    .X(_10108_));
 sky130_fd_sc_hd__o22a_1 _26022_ (.A1(_10019_),
    .A2(_10020_),
    .B1(_10014_),
    .B2(_10021_),
    .X(_10109_));
 sky130_fd_sc_hd__o22a_2 _26023_ (.A1(_10026_),
    .A2(_10033_),
    .B1(_10025_),
    .B2(_10034_),
    .X(_10110_));
 sky130_fd_sc_hd__o22a_1 _26024_ (.A1(_10008_),
    .A2(_07736_),
    .B1(_06391_),
    .B2(_08178_),
    .X(_10111_));
 sky130_fd_sc_hd__and4_1 _26025_ (.A(_13107_),
    .B(_13529_),
    .C(_13113_),
    .D(_13524_),
    .X(_10112_));
 sky130_fd_sc_hd__nor2_2 _26026_ (.A(_10111_),
    .B(_10112_),
    .Y(_10113_));
 sky130_fd_sc_hd__nor2_2 _26027_ (.A(_06286_),
    .B(_09007_),
    .Y(_10114_));
 sky130_fd_sc_hd__a2bb2o_1 _26028_ (.A1_N(_10113_),
    .A2_N(_10114_),
    .B1(_10113_),
    .B2(_10114_),
    .X(_10115_));
 sky130_fd_sc_hd__o22a_2 _26029_ (.A1(_09552_),
    .A2(_07468_),
    .B1(_06802_),
    .B2(_07033_),
    .X(_10116_));
 sky130_fd_sc_hd__and4_2 _26030_ (.A(_13098_),
    .B(_07466_),
    .C(_13103_),
    .D(_07598_),
    .X(_10117_));
 sky130_fd_sc_hd__nor2_2 _26031_ (.A(_10116_),
    .B(_10117_),
    .Y(_10118_));
 sky130_fd_sc_hd__nor2_2 _26032_ (.A(_06689_),
    .B(_09783_),
    .Y(_10119_));
 sky130_fd_sc_hd__a2bb2o_1 _26033_ (.A1_N(_10118_),
    .A2_N(_10119_),
    .B1(_10118_),
    .B2(_10119_),
    .X(_10120_));
 sky130_fd_sc_hd__a21oi_4 _26034_ (.A1(_10017_),
    .A2(_10018_),
    .B1(_10016_),
    .Y(_10121_));
 sky130_fd_sc_hd__a2bb2o_1 _26035_ (.A1_N(_10120_),
    .A2_N(_10121_),
    .B1(_10120_),
    .B2(_10121_),
    .X(_10122_));
 sky130_fd_sc_hd__a2bb2o_1 _26036_ (.A1_N(_10115_),
    .A2_N(_10122_),
    .B1(_10115_),
    .B2(_10122_),
    .X(_10123_));
 sky130_fd_sc_hd__a2bb2o_1 _26037_ (.A1_N(_10110_),
    .A2_N(_10123_),
    .B1(_10110_),
    .B2(_10123_),
    .X(_10124_));
 sky130_fd_sc_hd__a2bb2o_1 _26038_ (.A1_N(_10109_),
    .A2_N(_10124_),
    .B1(_10109_),
    .B2(_10124_),
    .X(_10125_));
 sky130_fd_sc_hd__a21oi_2 _26039_ (.A1(_10030_),
    .A2(_10032_),
    .B1(_10029_),
    .Y(_10126_));
 sky130_fd_sc_hd__a21oi_2 _26040_ (.A1(_10038_),
    .A2(_10039_),
    .B1(_10037_),
    .Y(_10127_));
 sky130_fd_sc_hd__o22a_1 _26041_ (.A1(_09436_),
    .A2(_07780_),
    .B1(_07272_),
    .B2(_06754_),
    .X(_10128_));
 sky130_fd_sc_hd__and4_1 _26042_ (.A(_10028_),
    .B(_13553_),
    .C(_09911_),
    .D(_07329_),
    .X(_10129_));
 sky130_fd_sc_hd__nor2_2 _26043_ (.A(_10128_),
    .B(_10129_),
    .Y(_10130_));
 sky130_fd_sc_hd__nor2_2 _26044_ (.A(_10031_),
    .B(_09025_),
    .Y(_10131_));
 sky130_fd_sc_hd__a2bb2o_1 _26045_ (.A1_N(_10130_),
    .A2_N(_10131_),
    .B1(_10130_),
    .B2(_10131_),
    .X(_10132_));
 sky130_fd_sc_hd__a2bb2o_1 _26046_ (.A1_N(_10127_),
    .A2_N(_10132_),
    .B1(_10127_),
    .B2(_10132_),
    .X(_10133_));
 sky130_fd_sc_hd__a2bb2o_1 _26047_ (.A1_N(_10126_),
    .A2_N(_10133_),
    .B1(_10126_),
    .B2(_10133_),
    .X(_10134_));
 sky130_fd_sc_hd__o22a_1 _26048_ (.A1(_09575_),
    .A2(_06227_),
    .B1(_09919_),
    .B2(_06339_),
    .X(_10135_));
 sky130_fd_sc_hd__and4_2 _26049_ (.A(_13074_),
    .B(_06768_),
    .C(_09806_),
    .D(_06899_),
    .X(_10136_));
 sky130_fd_sc_hd__nor2_2 _26050_ (.A(_10135_),
    .B(_10136_),
    .Y(_10137_));
 sky130_fd_sc_hd__nor2_4 _26051_ (.A(_07682_),
    .B(_06567_),
    .Y(_10138_));
 sky130_fd_sc_hd__a2bb2o_1 _26052_ (.A1_N(_10137_),
    .A2_N(_10138_),
    .B1(_10137_),
    .B2(_10138_),
    .X(_10139_));
 sky130_fd_sc_hd__buf_2 _26053_ (.A(_08295_),
    .X(_10140_));
 sky130_fd_sc_hd__and4_1 _26054_ (.A(_10140_),
    .B(_06030_),
    .C(_09191_),
    .D(_06462_),
    .X(_10141_));
 sky130_fd_sc_hd__o22a_1 _26055_ (.A1(_11718_),
    .A2(_13575_),
    .B1(_08132_),
    .B2(_06456_),
    .X(_10142_));
 sky130_fd_sc_hd__nor2_2 _26056_ (.A(_10141_),
    .B(_10142_),
    .Y(_10143_));
 sky130_fd_sc_hd__nor2_2 _26057_ (.A(_09188_),
    .B(_06140_),
    .Y(_10144_));
 sky130_fd_sc_hd__a2bb2o_1 _26058_ (.A1_N(_10143_),
    .A2_N(_10144_),
    .B1(_10143_),
    .B2(_10144_),
    .X(_10145_));
 sky130_fd_sc_hd__o21ba_1 _26059_ (.A1(_10041_),
    .A2(_10044_),
    .B1_N(_10042_),
    .X(_10146_));
 sky130_fd_sc_hd__a2bb2o_1 _26060_ (.A1_N(_10145_),
    .A2_N(_10146_),
    .B1(_10145_),
    .B2(_10146_),
    .X(_10147_));
 sky130_fd_sc_hd__a2bb2o_1 _26061_ (.A1_N(_10139_),
    .A2_N(_10147_),
    .B1(_10139_),
    .B2(_10147_),
    .X(_10148_));
 sky130_fd_sc_hd__o22a_1 _26062_ (.A1(_10045_),
    .A2(_10046_),
    .B1(_10040_),
    .B2(_10047_),
    .X(_10149_));
 sky130_fd_sc_hd__a2bb2o_1 _26063_ (.A1_N(_10148_),
    .A2_N(_10149_),
    .B1(_10148_),
    .B2(_10149_),
    .X(_10150_));
 sky130_fd_sc_hd__a2bb2o_2 _26064_ (.A1_N(_10134_),
    .A2_N(_10150_),
    .B1(_10134_),
    .B2(_10150_),
    .X(_10151_));
 sky130_fd_sc_hd__o22a_2 _26065_ (.A1(_10048_),
    .A2(_10049_),
    .B1(_10035_),
    .B2(_10050_),
    .X(_10152_));
 sky130_fd_sc_hd__a2bb2o_1 _26066_ (.A1_N(_10151_),
    .A2_N(_10152_),
    .B1(_10151_),
    .B2(_10152_),
    .X(_10153_));
 sky130_fd_sc_hd__a2bb2o_1 _26067_ (.A1_N(_10125_),
    .A2_N(_10153_),
    .B1(_10125_),
    .B2(_10153_),
    .X(_10154_));
 sky130_fd_sc_hd__o22a_1 _26068_ (.A1(_10051_),
    .A2(_10052_),
    .B1(_10024_),
    .B2(_10053_),
    .X(_10155_));
 sky130_fd_sc_hd__a2bb2o_1 _26069_ (.A1_N(_10154_),
    .A2_N(_10155_),
    .B1(_10154_),
    .B2(_10155_),
    .X(_10156_));
 sky130_fd_sc_hd__a2bb2o_1 _26070_ (.A1_N(_10108_),
    .A2_N(_10156_),
    .B1(_10108_),
    .B2(_10156_),
    .X(_10157_));
 sky130_fd_sc_hd__o22a_1 _26071_ (.A1(_10054_),
    .A2(_10055_),
    .B1(_10005_),
    .B2(_10056_),
    .X(_10158_));
 sky130_fd_sc_hd__a2bb2o_1 _26072_ (.A1_N(_10157_),
    .A2_N(_10158_),
    .B1(_10157_),
    .B2(_10158_),
    .X(_10159_));
 sky130_fd_sc_hd__a2bb2o_1 _26073_ (.A1_N(_10083_),
    .A2_N(_10159_),
    .B1(_10083_),
    .B2(_10159_),
    .X(_10160_));
 sky130_fd_sc_hd__o22a_1 _26074_ (.A1(_10057_),
    .A2(_10058_),
    .B1(_09979_),
    .B2(_10059_),
    .X(_10161_));
 sky130_fd_sc_hd__a2bb2o_1 _26075_ (.A1_N(_10160_),
    .A2_N(_10161_),
    .B1(_10160_),
    .B2(_10161_),
    .X(_10162_));
 sky130_fd_sc_hd__a2bb2o_1 _26076_ (.A1_N(_10072_),
    .A2_N(_10162_),
    .B1(_10072_),
    .B2(_10162_),
    .X(_10163_));
 sky130_fd_sc_hd__o22a_1 _26077_ (.A1(_10060_),
    .A2(_10061_),
    .B1(_09964_),
    .B2(_10062_),
    .X(_10164_));
 sky130_fd_sc_hd__a2bb2o_1 _26078_ (.A1_N(_10163_),
    .A2_N(_10164_),
    .B1(_10163_),
    .B2(_10164_),
    .X(_10165_));
 sky130_fd_sc_hd__a2bb2o_1 _26079_ (.A1_N(_09963_),
    .A2_N(_10165_),
    .B1(_09963_),
    .B2(_10165_),
    .X(_10166_));
 sky130_fd_sc_hd__o22a_1 _26080_ (.A1(_10063_),
    .A2(_10064_),
    .B1(_09842_),
    .B2(_10065_),
    .X(_10167_));
 sky130_fd_sc_hd__or2_1 _26081_ (.A(_10166_),
    .B(_10167_),
    .X(_10168_));
 sky130_fd_sc_hd__a21bo_1 _26082_ (.A1(_10166_),
    .A2(_10167_),
    .B1_N(_10168_),
    .X(_10169_));
 sky130_fd_sc_hd__a22o_1 _26083_ (.A1(_09961_),
    .A2(_10066_),
    .B1(_09952_),
    .B2(_10067_),
    .X(_10170_));
 sky130_fd_sc_hd__o31a_1 _26084_ (.A1(_09954_),
    .A2(_10068_),
    .A3(_09959_),
    .B1(_10170_),
    .X(_10171_));
 sky130_fd_sc_hd__a2bb2oi_1 _26085_ (.A1_N(_10169_),
    .A2_N(_10171_),
    .B1(_10169_),
    .B2(_10171_),
    .Y(_02665_));
 sky130_fd_sc_hd__o22a_1 _26086_ (.A1(_10163_),
    .A2(_10164_),
    .B1(_09963_),
    .B2(_10165_),
    .X(_10172_));
 sky130_fd_sc_hd__o22a_1 _26087_ (.A1(_10074_),
    .A2(_10081_),
    .B1(_10073_),
    .B2(_10082_),
    .X(_10173_));
 sky130_fd_sc_hd__or2_1 _26088_ (.A(_09350_),
    .B(_10173_),
    .X(_10174_));
 sky130_fd_sc_hd__a21bo_1 _26089_ (.A1(_09351_),
    .A2(_10173_),
    .B1_N(_10174_),
    .X(_10175_));
 sky130_fd_sc_hd__buf_1 _26090_ (.A(_09233_),
    .X(_10176_));
 sky130_fd_sc_hd__o22a_1 _26091_ (.A1(_10078_),
    .A2(_10079_),
    .B1(_10176_),
    .B2(_10080_),
    .X(_10177_));
 sky130_fd_sc_hd__o22a_1 _26092_ (.A1(_10085_),
    .A2(_10106_),
    .B1(_10084_),
    .B2(_10107_),
    .X(_10178_));
 sky130_fd_sc_hd__o22a_1 _26093_ (.A1(_09973_),
    .A2(_10076_),
    .B1(_10075_),
    .B2(_10077_),
    .X(_10179_));
 sky130_fd_sc_hd__o22ai_4 _26094_ (.A1(_10086_),
    .A2(_10093_),
    .B1(_10091_),
    .B2(_10087_),
    .Y(_10180_));
 sky130_fd_sc_hd__and3_1 _26095_ (.A(_09495_),
    .B(_09847_),
    .C(_09626_),
    .X(_10181_));
 sky130_fd_sc_hd__o21ba_1 _26096_ (.A1(_09738_),
    .A2(_09969_),
    .B1_N(_10181_),
    .X(_10182_));
 sky130_fd_sc_hd__a2bb2o_1 _26097_ (.A1_N(_10180_),
    .A2_N(_10182_),
    .B1(_10180_),
    .B2(_10182_),
    .X(_10183_));
 sky130_fd_sc_hd__o2bb2ai_1 _26098_ (.A1_N(_10179_),
    .A2_N(_10183_),
    .B1(_10179_),
    .B2(_10183_),
    .Y(_10184_));
 sky130_fd_sc_hd__a2bb2o_1 _26099_ (.A1_N(_09233_),
    .A2_N(_10184_),
    .B1(_09233_),
    .B2(_10184_),
    .X(_10185_));
 sky130_fd_sc_hd__a2bb2o_1 _26100_ (.A1_N(_10178_),
    .A2_N(_10185_),
    .B1(_10178_),
    .B2(_10185_),
    .X(_10186_));
 sky130_fd_sc_hd__a2bb2o_1 _26101_ (.A1_N(_10177_),
    .A2_N(_10186_),
    .B1(_10177_),
    .B2(_10186_),
    .X(_10187_));
 sky130_fd_sc_hd__o22a_1 _26102_ (.A1(_10103_),
    .A2(_10104_),
    .B1(_10094_),
    .B2(_10105_),
    .X(_10188_));
 sky130_fd_sc_hd__o22a_1 _26103_ (.A1(_10110_),
    .A2(_10123_),
    .B1(_10109_),
    .B2(_10124_),
    .X(_10189_));
 sky130_fd_sc_hd__o22ai_2 _26104_ (.A1(_10091_),
    .A2(_10087_),
    .B1(_09984_),
    .B2(_10089_),
    .Y(_10190_));
 sky130_fd_sc_hd__a2bb2o_2 _26105_ (.A1_N(_10086_),
    .A2_N(_10190_),
    .B1(_09754_),
    .B2(_10190_),
    .X(_10191_));
 sky130_fd_sc_hd__a21oi_2 _26106_ (.A1(_10099_),
    .A2(_10100_),
    .B1(_10098_),
    .Y(_10192_));
 sky130_fd_sc_hd__a21oi_2 _26107_ (.A1(_10113_),
    .A2(_10114_),
    .B1(_10112_),
    .Y(_10193_));
 sky130_fd_sc_hd__o22a_1 _26108_ (.A1(_09021_),
    .A2(_08838_),
    .B1(_06090_),
    .B2(_08035_),
    .X(_10194_));
 sky130_fd_sc_hd__and4_1 _26109_ (.A(_13119_),
    .B(_13510_),
    .C(_13123_),
    .D(_08820_),
    .X(_10195_));
 sky130_fd_sc_hd__nor2_1 _26110_ (.A(_10194_),
    .B(_10195_),
    .Y(_10196_));
 sky130_fd_sc_hd__or2_2 _26111_ (.A(_09867_),
    .B(_05998_),
    .X(_10197_));
 sky130_vsdinv _26112_ (.A(_10197_),
    .Y(_10198_));
 sky130_fd_sc_hd__buf_1 _26113_ (.A(_10198_),
    .X(_10199_));
 sky130_fd_sc_hd__a2bb2o_1 _26114_ (.A1_N(_10196_),
    .A2_N(_10199_),
    .B1(_10196_),
    .B2(_10198_),
    .X(_10200_));
 sky130_fd_sc_hd__a2bb2o_1 _26115_ (.A1_N(_10193_),
    .A2_N(_10200_),
    .B1(_10193_),
    .B2(_10200_),
    .X(_10201_));
 sky130_fd_sc_hd__a2bb2o_1 _26116_ (.A1_N(_10192_),
    .A2_N(_10201_),
    .B1(_10192_),
    .B2(_10201_),
    .X(_10202_));
 sky130_fd_sc_hd__o22a_1 _26117_ (.A1(_10096_),
    .A2(_10101_),
    .B1(_10095_),
    .B2(_10102_),
    .X(_10203_));
 sky130_fd_sc_hd__a2bb2o_1 _26118_ (.A1_N(_10202_),
    .A2_N(_10203_),
    .B1(_10202_),
    .B2(_10203_),
    .X(_10204_));
 sky130_fd_sc_hd__a2bb2o_1 _26119_ (.A1_N(_10191_),
    .A2_N(_10204_),
    .B1(_10191_),
    .B2(_10204_),
    .X(_10205_));
 sky130_fd_sc_hd__a2bb2o_1 _26120_ (.A1_N(_10189_),
    .A2_N(_10205_),
    .B1(_10189_),
    .B2(_10205_),
    .X(_10206_));
 sky130_fd_sc_hd__a2bb2o_1 _26121_ (.A1_N(_10188_),
    .A2_N(_10206_),
    .B1(_10188_),
    .B2(_10206_),
    .X(_10207_));
 sky130_fd_sc_hd__o22a_1 _26122_ (.A1(_10120_),
    .A2(_10121_),
    .B1(_10115_),
    .B2(_10122_),
    .X(_10208_));
 sky130_fd_sc_hd__o22a_2 _26123_ (.A1(_10127_),
    .A2(_10132_),
    .B1(_10126_),
    .B2(_10133_),
    .X(_10209_));
 sky130_fd_sc_hd__o22a_1 _26124_ (.A1(_09545_),
    .A2(_08684_),
    .B1(_06391_),
    .B2(_07870_),
    .X(_10210_));
 sky130_fd_sc_hd__and4_1 _26125_ (.A(_09547_),
    .B(_08686_),
    .C(_13113_),
    .D(_07877_),
    .X(_10211_));
 sky130_fd_sc_hd__nor2_2 _26126_ (.A(_10210_),
    .B(_10211_),
    .Y(_10212_));
 sky130_fd_sc_hd__nor2_1 _26127_ (.A(_06287_),
    .B(_08175_),
    .Y(_10213_));
 sky130_fd_sc_hd__a2bb2o_1 _26128_ (.A1_N(_10212_),
    .A2_N(_10213_),
    .B1(_10212_),
    .B2(_10213_),
    .X(_10214_));
 sky130_fd_sc_hd__buf_2 _26129_ (.A(_08262_),
    .X(_10215_));
 sky130_fd_sc_hd__clkbuf_4 _26130_ (.A(_07818_),
    .X(_10216_));
 sky130_fd_sc_hd__o22a_2 _26131_ (.A1(_10215_),
    .A2(_07033_),
    .B1(_10216_),
    .B2(_09782_),
    .X(_10217_));
 sky130_fd_sc_hd__and4_2 _26132_ (.A(_13098_),
    .B(_07598_),
    .C(_13103_),
    .D(_07886_),
    .X(_10218_));
 sky130_fd_sc_hd__nor2_2 _26133_ (.A(_10217_),
    .B(_10218_),
    .Y(_10219_));
 sky130_fd_sc_hd__nor2_2 _26134_ (.A(_06689_),
    .B(_09895_),
    .Y(_10220_));
 sky130_fd_sc_hd__a2bb2o_1 _26135_ (.A1_N(_10219_),
    .A2_N(_10220_),
    .B1(_10219_),
    .B2(_10220_),
    .X(_10221_));
 sky130_fd_sc_hd__a21oi_2 _26136_ (.A1(_10118_),
    .A2(_10119_),
    .B1(_10117_),
    .Y(_10222_));
 sky130_fd_sc_hd__a2bb2o_1 _26137_ (.A1_N(_10221_),
    .A2_N(_10222_),
    .B1(_10221_),
    .B2(_10222_),
    .X(_10223_));
 sky130_fd_sc_hd__a2bb2o_1 _26138_ (.A1_N(_10214_),
    .A2_N(_10223_),
    .B1(_10214_),
    .B2(_10223_),
    .X(_10224_));
 sky130_fd_sc_hd__a2bb2o_1 _26139_ (.A1_N(_10209_),
    .A2_N(_10224_),
    .B1(_10209_),
    .B2(_10224_),
    .X(_10225_));
 sky130_fd_sc_hd__a2bb2o_1 _26140_ (.A1_N(_10208_),
    .A2_N(_10225_),
    .B1(_10208_),
    .B2(_10225_),
    .X(_10226_));
 sky130_fd_sc_hd__a21oi_2 _26141_ (.A1(_10130_),
    .A2(_10131_),
    .B1(_10129_),
    .Y(_10227_));
 sky130_fd_sc_hd__a21oi_4 _26142_ (.A1(_10137_),
    .A2(_10138_),
    .B1(_10136_),
    .Y(_10228_));
 sky130_fd_sc_hd__buf_2 _26143_ (.A(_08599_),
    .X(_10229_));
 sky130_fd_sc_hd__o22a_1 _26144_ (.A1(_10229_),
    .A2(_06650_),
    .B1(_07272_),
    .B2(_07613_),
    .X(_10230_));
 sky130_fd_sc_hd__and4_2 _26145_ (.A(_10028_),
    .B(_13550_),
    .C(_09911_),
    .D(_07330_),
    .X(_10231_));
 sky130_fd_sc_hd__nor2_2 _26146_ (.A(_10230_),
    .B(_10231_),
    .Y(_10232_));
 sky130_fd_sc_hd__nor2_2 _26147_ (.A(_10031_),
    .B(_06892_),
    .Y(_10233_));
 sky130_fd_sc_hd__a2bb2o_1 _26148_ (.A1_N(_10232_),
    .A2_N(_10233_),
    .B1(_10232_),
    .B2(_10233_),
    .X(_10234_));
 sky130_fd_sc_hd__a2bb2o_1 _26149_ (.A1_N(_10228_),
    .A2_N(_10234_),
    .B1(_10228_),
    .B2(_10234_),
    .X(_10235_));
 sky130_fd_sc_hd__a2bb2o_2 _26150_ (.A1_N(_10227_),
    .A2_N(_10235_),
    .B1(_10227_),
    .B2(_10235_),
    .X(_10236_));
 sky130_fd_sc_hd__and4_2 _26151_ (.A(_09067_),
    .B(_06038_),
    .C(_13064_),
    .D(_13566_),
    .X(_10237_));
 sky130_fd_sc_hd__o22a_1 _26152_ (.A1(_08620_),
    .A2(_13569_),
    .B1(_09069_),
    .B2(_06139_),
    .X(_10238_));
 sky130_fd_sc_hd__nor2_2 _26153_ (.A(_10237_),
    .B(_10238_),
    .Y(_10239_));
 sky130_fd_sc_hd__nor2_4 _26154_ (.A(_08292_),
    .B(_08890_),
    .Y(_10240_));
 sky130_fd_sc_hd__a2bb2o_1 _26155_ (.A1_N(_10239_),
    .A2_N(_10240_),
    .B1(_10239_),
    .B2(_10240_),
    .X(_10241_));
 sky130_fd_sc_hd__a21oi_2 _26156_ (.A1(_10143_),
    .A2(_10144_),
    .B1(_10141_),
    .Y(_10242_));
 sky130_fd_sc_hd__o2bb2a_1 _26157_ (.A1_N(_10241_),
    .A2_N(_10242_),
    .B1(_10241_),
    .B2(_10242_),
    .X(_10243_));
 sky130_vsdinv _26158_ (.A(_10243_),
    .Y(_10244_));
 sky130_fd_sc_hd__o22a_1 _26159_ (.A1(_08611_),
    .A2(_09423_),
    .B1(_07684_),
    .B2(_08719_),
    .X(_10245_));
 sky130_fd_sc_hd__and4_2 _26160_ (.A(_08613_),
    .B(_13560_),
    .C(_13079_),
    .D(_08721_),
    .X(_10246_));
 sky130_fd_sc_hd__nor2_2 _26161_ (.A(_10245_),
    .B(_10246_),
    .Y(_10247_));
 sky130_fd_sc_hd__clkbuf_4 _26162_ (.A(_08388_),
    .X(_10248_));
 sky130_fd_sc_hd__nor2_2 _26163_ (.A(_09580_),
    .B(_10248_),
    .Y(_10249_));
 sky130_fd_sc_hd__a2bb2o_1 _26164_ (.A1_N(_10247_),
    .A2_N(_10249_),
    .B1(_10247_),
    .B2(_10249_),
    .X(_10250_));
 sky130_vsdinv _26165_ (.A(_10250_),
    .Y(_10251_));
 sky130_fd_sc_hd__a22o_2 _26166_ (.A1(_10244_),
    .A2(_10250_),
    .B1(_10243_),
    .B2(_10251_),
    .X(_10252_));
 sky130_fd_sc_hd__o22a_2 _26167_ (.A1(_10145_),
    .A2(_10146_),
    .B1(_10139_),
    .B2(_10147_),
    .X(_10253_));
 sky130_fd_sc_hd__a2bb2o_1 _26168_ (.A1_N(_10252_),
    .A2_N(_10253_),
    .B1(_10252_),
    .B2(_10253_),
    .X(_10254_));
 sky130_fd_sc_hd__a2bb2o_1 _26169_ (.A1_N(_10236_),
    .A2_N(_10254_),
    .B1(_10236_),
    .B2(_10254_),
    .X(_10255_));
 sky130_fd_sc_hd__o22a_2 _26170_ (.A1(_10148_),
    .A2(_10149_),
    .B1(_10134_),
    .B2(_10150_),
    .X(_10256_));
 sky130_fd_sc_hd__a2bb2o_1 _26171_ (.A1_N(_10255_),
    .A2_N(_10256_),
    .B1(_10255_),
    .B2(_10256_),
    .X(_10257_));
 sky130_fd_sc_hd__a2bb2o_1 _26172_ (.A1_N(_10226_),
    .A2_N(_10257_),
    .B1(_10226_),
    .B2(_10257_),
    .X(_10258_));
 sky130_fd_sc_hd__o22a_1 _26173_ (.A1(_10151_),
    .A2(_10152_),
    .B1(_10125_),
    .B2(_10153_),
    .X(_10259_));
 sky130_fd_sc_hd__a2bb2o_1 _26174_ (.A1_N(_10258_),
    .A2_N(_10259_),
    .B1(_10258_),
    .B2(_10259_),
    .X(_10260_));
 sky130_fd_sc_hd__a2bb2o_1 _26175_ (.A1_N(_10207_),
    .A2_N(_10260_),
    .B1(_10207_),
    .B2(_10260_),
    .X(_10261_));
 sky130_fd_sc_hd__o22a_1 _26176_ (.A1(_10154_),
    .A2(_10155_),
    .B1(_10108_),
    .B2(_10156_),
    .X(_10262_));
 sky130_fd_sc_hd__a2bb2o_1 _26177_ (.A1_N(_10261_),
    .A2_N(_10262_),
    .B1(_10261_),
    .B2(_10262_),
    .X(_10263_));
 sky130_fd_sc_hd__a2bb2o_1 _26178_ (.A1_N(_10187_),
    .A2_N(_10263_),
    .B1(_10187_),
    .B2(_10263_),
    .X(_10264_));
 sky130_fd_sc_hd__o22a_1 _26179_ (.A1(_10157_),
    .A2(_10158_),
    .B1(_10083_),
    .B2(_10159_),
    .X(_10265_));
 sky130_fd_sc_hd__a2bb2o_1 _26180_ (.A1_N(_10264_),
    .A2_N(_10265_),
    .B1(_10264_),
    .B2(_10265_),
    .X(_10266_));
 sky130_fd_sc_hd__a2bb2o_1 _26181_ (.A1_N(_10175_),
    .A2_N(_10266_),
    .B1(_10175_),
    .B2(_10266_),
    .X(_10267_));
 sky130_fd_sc_hd__o22a_1 _26182_ (.A1(_10160_),
    .A2(_10161_),
    .B1(_10072_),
    .B2(_10162_),
    .X(_10268_));
 sky130_fd_sc_hd__a2bb2o_1 _26183_ (.A1_N(_10267_),
    .A2_N(_10268_),
    .B1(_10267_),
    .B2(_10268_),
    .X(_10269_));
 sky130_fd_sc_hd__a2bb2o_1 _26184_ (.A1_N(_10071_),
    .A2_N(_10269_),
    .B1(_10071_),
    .B2(_10269_),
    .X(_10270_));
 sky130_fd_sc_hd__and2_1 _26185_ (.A(_10172_),
    .B(_10270_),
    .X(_10271_));
 sky130_fd_sc_hd__or2_1 _26186_ (.A(_10172_),
    .B(_10270_),
    .X(_10272_));
 sky130_fd_sc_hd__or2b_1 _26187_ (.A(_10271_),
    .B_N(_10272_),
    .X(_10273_));
 sky130_fd_sc_hd__o21ai_1 _26188_ (.A1(_10169_),
    .A2(_10171_),
    .B1(_10168_),
    .Y(_10274_));
 sky130_fd_sc_hd__a2bb2o_1 _26189_ (.A1_N(_10273_),
    .A2_N(_10274_),
    .B1(_10273_),
    .B2(_10274_),
    .X(_02666_));
 sky130_fd_sc_hd__buf_1 _26190_ (.A(_09352_),
    .X(_10275_));
 sky130_fd_sc_hd__clkbuf_2 _26191_ (.A(_10275_),
    .X(_10276_));
 sky130_fd_sc_hd__o22a_1 _26192_ (.A1(_10178_),
    .A2(_10185_),
    .B1(_10177_),
    .B2(_10186_),
    .X(_10277_));
 sky130_fd_sc_hd__clkbuf_2 _26193_ (.A(_09352_),
    .X(_10278_));
 sky130_fd_sc_hd__or2_1 _26194_ (.A(_10278_),
    .B(_10277_),
    .X(_10279_));
 sky130_fd_sc_hd__a21bo_1 _26195_ (.A1(_10276_),
    .A2(_10277_),
    .B1_N(_10279_),
    .X(_10280_));
 sky130_fd_sc_hd__buf_1 _26196_ (.A(_10176_),
    .X(_10281_));
 sky130_fd_sc_hd__o22a_1 _26197_ (.A1(_10179_),
    .A2(_10183_),
    .B1(_10281_),
    .B2(_10184_),
    .X(_10282_));
 sky130_fd_sc_hd__o22a_1 _26198_ (.A1(_10189_),
    .A2(_10205_),
    .B1(_10188_),
    .B2(_10206_),
    .X(_10283_));
 sky130_fd_sc_hd__o22a_1 _26199_ (.A1(_10091_),
    .A2(_10087_),
    .B1(_09874_),
    .B2(_10190_),
    .X(_10284_));
 sky130_fd_sc_hd__o22ai_1 _26200_ (.A1(_09738_),
    .A2(_09969_),
    .B1(_10180_),
    .B2(_10181_),
    .Y(_10285_));
 sky130_fd_sc_hd__o2bb2a_1 _26201_ (.A1_N(_10284_),
    .A2_N(_10285_),
    .B1(_10284_),
    .B2(_10285_),
    .X(_10286_));
 sky130_fd_sc_hd__a2bb2o_1 _26202_ (.A1_N(_10281_),
    .A2_N(_10286_),
    .B1(_10176_),
    .B2(_10286_),
    .X(_10287_));
 sky130_fd_sc_hd__a2bb2o_1 _26203_ (.A1_N(_10283_),
    .A2_N(_10287_),
    .B1(_10283_),
    .B2(_10287_),
    .X(_10288_));
 sky130_fd_sc_hd__a2bb2o_1 _26204_ (.A1_N(_10282_),
    .A2_N(_10288_),
    .B1(_10282_),
    .B2(_10288_),
    .X(_10289_));
 sky130_fd_sc_hd__buf_1 _26205_ (.A(_10191_),
    .X(_10290_));
 sky130_fd_sc_hd__clkbuf_2 _26206_ (.A(_10290_),
    .X(_10291_));
 sky130_fd_sc_hd__o22a_1 _26207_ (.A1(_10202_),
    .A2(_10203_),
    .B1(_10291_),
    .B2(_10204_),
    .X(_10292_));
 sky130_fd_sc_hd__o22a_1 _26208_ (.A1(_10209_),
    .A2(_10224_),
    .B1(_10208_),
    .B2(_10225_),
    .X(_10293_));
 sky130_fd_sc_hd__buf_1 _26209_ (.A(_10191_),
    .X(_10294_));
 sky130_fd_sc_hd__buf_1 _26210_ (.A(_10294_),
    .X(_10295_));
 sky130_fd_sc_hd__a31o_1 _26211_ (.A1(\pcpi_mul.rs2[18] ),
    .A2(_13517_),
    .A3(_10212_),
    .B1(_10211_),
    .X(_10296_));
 sky130_fd_sc_hd__o22a_1 _26212_ (.A1(_07941_),
    .A2(_08034_),
    .B1(_09867_),
    .B2(_08401_),
    .X(_10297_));
 sky130_fd_sc_hd__and4_1 _26213_ (.A(_13118_),
    .B(_13505_),
    .C(_08814_),
    .D(_13122_),
    .X(_10298_));
 sky130_fd_sc_hd__or2_1 _26214_ (.A(_10297_),
    .B(_10298_),
    .X(_10299_));
 sky130_vsdinv _26215_ (.A(_10299_),
    .Y(_10300_));
 sky130_fd_sc_hd__o22a_1 _26216_ (.A1(_10197_),
    .A2(_10299_),
    .B1(_10199_),
    .B2(_10300_),
    .X(_10301_));
 sky130_vsdinv _26217_ (.A(_10296_),
    .Y(_10302_));
 sky130_vsdinv _26218_ (.A(_10301_),
    .Y(_10303_));
 sky130_fd_sc_hd__o22a_1 _26219_ (.A1(_10296_),
    .A2(_10301_),
    .B1(_10302_),
    .B2(_10303_),
    .X(_10304_));
 sky130_fd_sc_hd__clkbuf_2 _26220_ (.A(_10088_),
    .X(_10305_));
 sky130_fd_sc_hd__a31o_1 _26221_ (.A1(_10305_),
    .A2(_13126_),
    .A3(_10196_),
    .B1(_10195_),
    .X(_10306_));
 sky130_vsdinv _26222_ (.A(_10304_),
    .Y(_10307_));
 sky130_vsdinv _26223_ (.A(_10306_),
    .Y(_10308_));
 sky130_fd_sc_hd__o22a_1 _26224_ (.A1(_10304_),
    .A2(_10306_),
    .B1(_10307_),
    .B2(_10308_),
    .X(_10309_));
 sky130_vsdinv _26225_ (.A(_10309_),
    .Y(_10310_));
 sky130_fd_sc_hd__o22a_1 _26226_ (.A1(_10193_),
    .A2(_10200_),
    .B1(_10192_),
    .B2(_10201_),
    .X(_10311_));
 sky130_vsdinv _26227_ (.A(_10311_),
    .Y(_10312_));
 sky130_fd_sc_hd__a22o_1 _26228_ (.A1(_10310_),
    .A2(_10311_),
    .B1(_10309_),
    .B2(_10312_),
    .X(_10313_));
 sky130_fd_sc_hd__buf_1 _26229_ (.A(_10294_),
    .X(_10314_));
 sky130_fd_sc_hd__a2bb2o_1 _26230_ (.A1_N(_10295_),
    .A2_N(_10313_),
    .B1(_10314_),
    .B2(_10313_),
    .X(_10315_));
 sky130_fd_sc_hd__a2bb2o_1 _26231_ (.A1_N(_10293_),
    .A2_N(_10315_),
    .B1(_10293_),
    .B2(_10315_),
    .X(_10316_));
 sky130_fd_sc_hd__a2bb2o_1 _26232_ (.A1_N(_10292_),
    .A2_N(_10316_),
    .B1(_10292_),
    .B2(_10316_),
    .X(_10317_));
 sky130_fd_sc_hd__o22a_1 _26233_ (.A1(_10221_),
    .A2(_10222_),
    .B1(_10214_),
    .B2(_10223_),
    .X(_10318_));
 sky130_fd_sc_hd__o22a_2 _26234_ (.A1(_10228_),
    .A2(_10234_),
    .B1(_10227_),
    .B2(_10235_),
    .X(_10319_));
 sky130_fd_sc_hd__o22a_1 _26235_ (.A1(_10008_),
    .A2(_07871_),
    .B1(_06392_),
    .B2(_07874_),
    .X(_10320_));
 sky130_fd_sc_hd__and4_2 _26236_ (.A(_13107_),
    .B(_07878_),
    .C(_13114_),
    .D(_13516_),
    .X(_10321_));
 sky130_fd_sc_hd__nor2_2 _26237_ (.A(_10320_),
    .B(_10321_),
    .Y(_10322_));
 sky130_fd_sc_hd__buf_2 _26238_ (.A(_08839_),
    .X(_10323_));
 sky130_fd_sc_hd__nor2_2 _26239_ (.A(_06286_),
    .B(_10323_),
    .Y(_10324_));
 sky130_fd_sc_hd__a2bb2o_1 _26240_ (.A1_N(_10322_),
    .A2_N(_10324_),
    .B1(_10322_),
    .B2(_10324_),
    .X(_10325_));
 sky130_fd_sc_hd__buf_1 _26241_ (.A(_10215_),
    .X(_10326_));
 sky130_fd_sc_hd__clkbuf_2 _26242_ (.A(_09783_),
    .X(_10327_));
 sky130_fd_sc_hd__buf_1 _26243_ (.A(_10216_),
    .X(_10328_));
 sky130_fd_sc_hd__clkbuf_2 _26244_ (.A(_09895_),
    .X(_10329_));
 sky130_fd_sc_hd__o22a_1 _26245_ (.A1(_10326_),
    .A2(_10327_),
    .B1(_10328_),
    .B2(_10329_),
    .X(_10330_));
 sky130_fd_sc_hd__and4_2 _26246_ (.A(_13099_),
    .B(_13536_),
    .C(_13104_),
    .D(_13530_),
    .X(_10331_));
 sky130_fd_sc_hd__nor2_2 _26247_ (.A(_10330_),
    .B(_10331_),
    .Y(_10332_));
 sky130_fd_sc_hd__clkbuf_2 _26248_ (.A(_06689_),
    .X(_10333_));
 sky130_fd_sc_hd__clkbuf_2 _26249_ (.A(_10012_),
    .X(_10334_));
 sky130_fd_sc_hd__nor2_2 _26250_ (.A(_10333_),
    .B(_10334_),
    .Y(_10335_));
 sky130_fd_sc_hd__a2bb2o_1 _26251_ (.A1_N(_10332_),
    .A2_N(_10335_),
    .B1(_10332_),
    .B2(_10335_),
    .X(_10336_));
 sky130_fd_sc_hd__a21oi_2 _26252_ (.A1(_10219_),
    .A2(_10220_),
    .B1(_10218_),
    .Y(_10337_));
 sky130_fd_sc_hd__a2bb2o_1 _26253_ (.A1_N(_10336_),
    .A2_N(_10337_),
    .B1(_10336_),
    .B2(_10337_),
    .X(_10338_));
 sky130_fd_sc_hd__a2bb2o_1 _26254_ (.A1_N(_10325_),
    .A2_N(_10338_),
    .B1(_10325_),
    .B2(_10338_),
    .X(_10339_));
 sky130_fd_sc_hd__a2bb2o_1 _26255_ (.A1_N(_10319_),
    .A2_N(_10339_),
    .B1(_10319_),
    .B2(_10339_),
    .X(_10340_));
 sky130_fd_sc_hd__a2bb2o_1 _26256_ (.A1_N(_10318_),
    .A2_N(_10340_),
    .B1(_10318_),
    .B2(_10340_),
    .X(_10341_));
 sky130_fd_sc_hd__clkbuf_2 _26257_ (.A(_10140_),
    .X(_10342_));
 sky130_fd_sc_hd__and4_4 _26258_ (.A(_10342_),
    .B(_06581_),
    .C(_13065_),
    .D(_06768_),
    .X(_10343_));
 sky130_fd_sc_hd__buf_1 _26259_ (.A(_11718_),
    .X(_10344_));
 sky130_fd_sc_hd__buf_1 _26260_ (.A(_08926_),
    .X(_10345_));
 sky130_fd_sc_hd__o22a_2 _26261_ (.A1(_10344_),
    .A2(_13568_),
    .B1(_10345_),
    .B2(_06330_),
    .X(_10346_));
 sky130_fd_sc_hd__nor2_2 _26262_ (.A(_10343_),
    .B(_10346_),
    .Y(_10347_));
 sky130_fd_sc_hd__clkbuf_4 _26263_ (.A(_07972_),
    .X(_10348_));
 sky130_fd_sc_hd__nor2_4 _26264_ (.A(_10348_),
    .B(_06439_),
    .Y(_10349_));
 sky130_fd_sc_hd__a2bb2o_2 _26265_ (.A1_N(_10347_),
    .A2_N(_10349_),
    .B1(_10347_),
    .B2(_10349_),
    .X(_10350_));
 sky130_fd_sc_hd__a21oi_4 _26266_ (.A1(_10239_),
    .A2(_10240_),
    .B1(_10237_),
    .Y(_10351_));
 sky130_fd_sc_hd__o2bb2ai_2 _26267_ (.A1_N(_10350_),
    .A2_N(_10351_),
    .B1(_10350_),
    .B2(_10351_),
    .Y(_10352_));
 sky130_fd_sc_hd__buf_1 _26268_ (.A(_09918_),
    .X(_10353_));
 sky130_fd_sc_hd__o22a_1 _26269_ (.A1(_10353_),
    .A2(_06452_),
    .B1(_07680_),
    .B2(_06642_),
    .X(_10354_));
 sky130_fd_sc_hd__clkbuf_2 _26270_ (.A(_09577_),
    .X(_10355_));
 sky130_fd_sc_hd__and4_2 _26271_ (.A(_10355_),
    .B(_13557_),
    .C(_13080_),
    .D(_13554_),
    .X(_10356_));
 sky130_fd_sc_hd__nor2_2 _26272_ (.A(_10354_),
    .B(_10356_),
    .Y(_10357_));
 sky130_fd_sc_hd__clkbuf_4 _26273_ (.A(_07532_),
    .X(_10358_));
 sky130_fd_sc_hd__nor2_2 _26274_ (.A(_10358_),
    .B(_06879_),
    .Y(_10359_));
 sky130_fd_sc_hd__a2bb2o_2 _26275_ (.A1_N(_10357_),
    .A2_N(_10359_),
    .B1(_10357_),
    .B2(_10359_),
    .X(_10360_));
 sky130_fd_sc_hd__o2bb2ai_2 _26276_ (.A1_N(_10352_),
    .A2_N(_10360_),
    .B1(_10352_),
    .B2(_10360_),
    .Y(_10361_));
 sky130_fd_sc_hd__o22a_2 _26277_ (.A1(_10241_),
    .A2(_10242_),
    .B1(_10244_),
    .B2(_10250_),
    .X(_10362_));
 sky130_fd_sc_hd__o2bb2a_1 _26278_ (.A1_N(_10361_),
    .A2_N(_10362_),
    .B1(_10361_),
    .B2(_10362_),
    .X(_10363_));
 sky130_vsdinv _26279_ (.A(_10363_),
    .Y(_10364_));
 sky130_fd_sc_hd__a21oi_4 _26280_ (.A1(_10232_),
    .A2(_10233_),
    .B1(_10231_),
    .Y(_10365_));
 sky130_fd_sc_hd__a21oi_4 _26281_ (.A1(_10247_),
    .A2(_10249_),
    .B1(_10246_),
    .Y(_10366_));
 sky130_fd_sc_hd__clkbuf_2 _26282_ (.A(_10229_),
    .X(_10367_));
 sky130_fd_sc_hd__buf_1 _26283_ (.A(_07272_),
    .X(_10368_));
 sky130_fd_sc_hd__o22a_1 _26284_ (.A1(_10367_),
    .A2(_07178_),
    .B1(_10368_),
    .B2(_07321_),
    .X(_10369_));
 sky130_fd_sc_hd__buf_1 _26285_ (.A(_10028_),
    .X(_10370_));
 sky130_fd_sc_hd__buf_1 _26286_ (.A(_13093_),
    .X(_10371_));
 sky130_fd_sc_hd__and4_1 _26287_ (.A(_10370_),
    .B(_13547_),
    .C(_10371_),
    .D(_13543_),
    .X(_10372_));
 sky130_fd_sc_hd__nor2_2 _26288_ (.A(_10369_),
    .B(_10372_),
    .Y(_10373_));
 sky130_fd_sc_hd__buf_2 _26289_ (.A(_10031_),
    .X(_10374_));
 sky130_fd_sc_hd__buf_2 _26290_ (.A(_07173_),
    .X(_10375_));
 sky130_fd_sc_hd__nor2_2 _26291_ (.A(_10374_),
    .B(_10375_),
    .Y(_10376_));
 sky130_fd_sc_hd__a2bb2o_2 _26292_ (.A1_N(_10373_),
    .A2_N(_10376_),
    .B1(_10373_),
    .B2(_10376_),
    .X(_10377_));
 sky130_fd_sc_hd__a2bb2o_1 _26293_ (.A1_N(_10366_),
    .A2_N(_10377_),
    .B1(_10366_),
    .B2(_10377_),
    .X(_10378_));
 sky130_fd_sc_hd__a2bb2o_1 _26294_ (.A1_N(_10365_),
    .A2_N(_10378_),
    .B1(_10365_),
    .B2(_10378_),
    .X(_10379_));
 sky130_vsdinv _26295_ (.A(_10379_),
    .Y(_10380_));
 sky130_fd_sc_hd__a22o_1 _26296_ (.A1(_10364_),
    .A2(_10379_),
    .B1(_10363_),
    .B2(_10380_),
    .X(_10381_));
 sky130_fd_sc_hd__o22a_1 _26297_ (.A1(_10252_),
    .A2(_10253_),
    .B1(_10236_),
    .B2(_10254_),
    .X(_10382_));
 sky130_fd_sc_hd__a2bb2o_1 _26298_ (.A1_N(_10381_),
    .A2_N(_10382_),
    .B1(_10381_),
    .B2(_10382_),
    .X(_10383_));
 sky130_fd_sc_hd__a2bb2o_1 _26299_ (.A1_N(_10341_),
    .A2_N(_10383_),
    .B1(_10341_),
    .B2(_10383_),
    .X(_10384_));
 sky130_fd_sc_hd__o22a_1 _26300_ (.A1(_10255_),
    .A2(_10256_),
    .B1(_10226_),
    .B2(_10257_),
    .X(_10385_));
 sky130_fd_sc_hd__a2bb2o_1 _26301_ (.A1_N(_10384_),
    .A2_N(_10385_),
    .B1(_10384_),
    .B2(_10385_),
    .X(_10386_));
 sky130_fd_sc_hd__a2bb2o_1 _26302_ (.A1_N(_10317_),
    .A2_N(_10386_),
    .B1(_10317_),
    .B2(_10386_),
    .X(_10387_));
 sky130_fd_sc_hd__o22a_1 _26303_ (.A1(_10258_),
    .A2(_10259_),
    .B1(_10207_),
    .B2(_10260_),
    .X(_10388_));
 sky130_fd_sc_hd__a2bb2o_1 _26304_ (.A1_N(_10387_),
    .A2_N(_10388_),
    .B1(_10387_),
    .B2(_10388_),
    .X(_10389_));
 sky130_fd_sc_hd__a2bb2o_1 _26305_ (.A1_N(_10289_),
    .A2_N(_10389_),
    .B1(_10289_),
    .B2(_10389_),
    .X(_10390_));
 sky130_fd_sc_hd__o22a_1 _26306_ (.A1(_10261_),
    .A2(_10262_),
    .B1(_10187_),
    .B2(_10263_),
    .X(_10391_));
 sky130_fd_sc_hd__a2bb2o_1 _26307_ (.A1_N(_10390_),
    .A2_N(_10391_),
    .B1(_10390_),
    .B2(_10391_),
    .X(_10392_));
 sky130_fd_sc_hd__a2bb2o_1 _26308_ (.A1_N(_10280_),
    .A2_N(_10392_),
    .B1(_10280_),
    .B2(_10392_),
    .X(_10393_));
 sky130_fd_sc_hd__o22a_1 _26309_ (.A1(_10264_),
    .A2(_10265_),
    .B1(_10175_),
    .B2(_10266_),
    .X(_10394_));
 sky130_fd_sc_hd__a2bb2o_1 _26310_ (.A1_N(_10393_),
    .A2_N(_10394_),
    .B1(_10393_),
    .B2(_10394_),
    .X(_10395_));
 sky130_fd_sc_hd__a2bb2o_1 _26311_ (.A1_N(_10174_),
    .A2_N(_10395_),
    .B1(_10174_),
    .B2(_10395_),
    .X(_10396_));
 sky130_fd_sc_hd__o22a_1 _26312_ (.A1(_10267_),
    .A2(_10268_),
    .B1(_10071_),
    .B2(_10269_),
    .X(_10397_));
 sky130_fd_sc_hd__or2_1 _26313_ (.A(_10396_),
    .B(_10397_),
    .X(_10398_));
 sky130_fd_sc_hd__a21bo_1 _26314_ (.A1(_10396_),
    .A2(_10397_),
    .B1_N(_10398_),
    .X(_10399_));
 sky130_fd_sc_hd__buf_1 _26315_ (.A(_10399_),
    .X(_10400_));
 sky130_fd_sc_hd__or2_1 _26316_ (.A(_10169_),
    .B(_10273_),
    .X(_10401_));
 sky130_fd_sc_hd__or3_4 _26317_ (.A(_09953_),
    .B(_10068_),
    .C(_10401_),
    .X(_10402_));
 sky130_fd_sc_hd__or2_1 _26318_ (.A(_09956_),
    .B(_10402_),
    .X(_10403_));
 sky130_fd_sc_hd__o221a_1 _26319_ (.A1(_10168_),
    .A2(_10271_),
    .B1(_10170_),
    .B2(_10401_),
    .C1(_10272_),
    .X(_10404_));
 sky130_fd_sc_hd__o221a_1 _26320_ (.A1(_09957_),
    .A2(_10402_),
    .B1(_09484_),
    .B2(_10403_),
    .C1(_10404_),
    .X(_10405_));
 sky130_fd_sc_hd__o31a_4 _26321_ (.A1(_09481_),
    .A2(_10403_),
    .A3(_08328_),
    .B1(_10405_),
    .X(_10406_));
 sky130_fd_sc_hd__buf_1 _26322_ (.A(_10406_),
    .X(_10407_));
 sky130_fd_sc_hd__a2bb2oi_1 _26323_ (.A1_N(_10400_),
    .A2_N(_10407_),
    .B1(_10400_),
    .B2(_10407_),
    .Y(_02667_));
 sky130_fd_sc_hd__o21ai_1 _26324_ (.A1(_10400_),
    .A2(_10407_),
    .B1(_10398_),
    .Y(_10408_));
 sky130_fd_sc_hd__o22a_1 _26325_ (.A1(_10283_),
    .A2(_10287_),
    .B1(_10282_),
    .B2(_10288_),
    .X(_10409_));
 sky130_fd_sc_hd__clkbuf_2 _26326_ (.A(_09489_),
    .X(_10410_));
 sky130_fd_sc_hd__or2_1 _26327_ (.A(_10410_),
    .B(_10409_),
    .X(_10411_));
 sky130_fd_sc_hd__a21bo_1 _26328_ (.A1(_10275_),
    .A2(_10409_),
    .B1_N(_10411_),
    .X(_10412_));
 sky130_fd_sc_hd__or3_1 _26329_ (.A(_09738_),
    .B(_09969_),
    .C(_10284_),
    .X(_10413_));
 sky130_fd_sc_hd__buf_1 _26330_ (.A(_10413_),
    .X(_10414_));
 sky130_fd_sc_hd__o21a_1 _26331_ (.A1(_10281_),
    .A2(_10286_),
    .B1(_10414_),
    .X(_10415_));
 sky130_fd_sc_hd__o22a_1 _26332_ (.A1(_10293_),
    .A2(_10315_),
    .B1(_10292_),
    .B2(_10316_),
    .X(_10416_));
 sky130_fd_sc_hd__nand2_1 _26333_ (.A(_10181_),
    .B(_10284_),
    .Y(_10417_));
 sky130_vsdinv _26334_ (.A(_09232_),
    .Y(_10418_));
 sky130_fd_sc_hd__nand2_1 _26335_ (.A(_10413_),
    .B(_10417_),
    .Y(_10419_));
 sky130_fd_sc_hd__a32o_1 _26336_ (.A1(_10414_),
    .A2(_10417_),
    .A3(_10418_),
    .B1(_09616_),
    .B2(_10419_),
    .X(_10420_));
 sky130_fd_sc_hd__buf_1 _26337_ (.A(_10420_),
    .X(_10421_));
 sky130_fd_sc_hd__a2bb2o_1 _26338_ (.A1_N(_10416_),
    .A2_N(_10421_),
    .B1(_10416_),
    .B2(_10421_),
    .X(_10422_));
 sky130_fd_sc_hd__a2bb2o_1 _26339_ (.A1_N(_10415_),
    .A2_N(_10422_),
    .B1(_10415_),
    .B2(_10422_),
    .X(_10423_));
 sky130_fd_sc_hd__buf_1 _26340_ (.A(_10295_),
    .X(_10424_));
 sky130_fd_sc_hd__o22a_1 _26341_ (.A1(_10310_),
    .A2(_10311_),
    .B1(_10424_),
    .B2(_10313_),
    .X(_10425_));
 sky130_fd_sc_hd__o22a_1 _26342_ (.A1(_10319_),
    .A2(_10339_),
    .B1(_10318_),
    .B2(_10340_),
    .X(_10426_));
 sky130_fd_sc_hd__buf_1 _26343_ (.A(_10290_),
    .X(_10427_));
 sky130_fd_sc_hd__a21oi_2 _26344_ (.A1(_10322_),
    .A2(_10324_),
    .B1(_10321_),
    .Y(_10428_));
 sky130_fd_sc_hd__or4_4 _26345_ (.A(_11702_),
    .B(_06093_),
    .C(_11702_),
    .D(_07253_),
    .X(_10429_));
 sky130_fd_sc_hd__buf_1 _26346_ (.A(_10429_),
    .X(_10430_));
 sky130_fd_sc_hd__o22a_2 _26347_ (.A1(_08660_),
    .A2(_08870_),
    .B1(_08660_),
    .B2(_09021_),
    .X(_10431_));
 sky130_vsdinv _26348_ (.A(_10431_),
    .Y(_10432_));
 sky130_vsdinv _26349_ (.A(_10429_),
    .Y(_10433_));
 sky130_fd_sc_hd__or2_1 _26350_ (.A(_10433_),
    .B(_10431_),
    .X(_10434_));
 sky130_fd_sc_hd__a32o_1 _26351_ (.A1(_10430_),
    .A2(_10432_),
    .A3(_10199_),
    .B1(_10197_),
    .B2(_10434_),
    .X(_10435_));
 sky130_fd_sc_hd__o2bb2a_1 _26352_ (.A1_N(_10428_),
    .A2_N(_10435_),
    .B1(_10428_),
    .B2(_10435_),
    .X(_10436_));
 sky130_fd_sc_hd__a31o_1 _26353_ (.A1(_10305_),
    .A2(_13126_),
    .A3(_10300_),
    .B1(_10298_),
    .X(_10437_));
 sky130_vsdinv _26354_ (.A(_10436_),
    .Y(_10438_));
 sky130_vsdinv _26355_ (.A(_10437_),
    .Y(_10439_));
 sky130_fd_sc_hd__o22a_1 _26356_ (.A1(_10436_),
    .A2(_10437_),
    .B1(_10438_),
    .B2(_10439_),
    .X(_10440_));
 sky130_vsdinv _26357_ (.A(_10440_),
    .Y(_10441_));
 sky130_fd_sc_hd__o22a_1 _26358_ (.A1(_10302_),
    .A2(_10303_),
    .B1(_10307_),
    .B2(_10308_),
    .X(_10442_));
 sky130_vsdinv _26359_ (.A(_10442_),
    .Y(_10443_));
 sky130_fd_sc_hd__a22o_1 _26360_ (.A1(_10441_),
    .A2(_10442_),
    .B1(_10440_),
    .B2(_10443_),
    .X(_10444_));
 sky130_fd_sc_hd__a2bb2o_1 _26361_ (.A1_N(_10427_),
    .A2_N(_10444_),
    .B1(_10427_),
    .B2(_10444_),
    .X(_10445_));
 sky130_fd_sc_hd__a2bb2o_1 _26362_ (.A1_N(_10426_),
    .A2_N(_10445_),
    .B1(_10426_),
    .B2(_10445_),
    .X(_10446_));
 sky130_fd_sc_hd__a2bb2o_1 _26363_ (.A1_N(_10425_),
    .A2_N(_10446_),
    .B1(_10425_),
    .B2(_10446_),
    .X(_10447_));
 sky130_fd_sc_hd__and4_2 _26364_ (.A(_10140_),
    .B(_08890_),
    .C(_13065_),
    .D(_06899_),
    .X(_10448_));
 sky130_fd_sc_hd__o22a_1 _26365_ (.A1(_10344_),
    .A2(_13565_),
    .B1(_10345_),
    .B2(_06438_),
    .X(_10449_));
 sky130_fd_sc_hd__nor2_2 _26366_ (.A(_10448_),
    .B(_10449_),
    .Y(_10450_));
 sky130_fd_sc_hd__nor2_4 _26367_ (.A(_07972_),
    .B(_06452_),
    .Y(_10451_));
 sky130_fd_sc_hd__a2bb2o_2 _26368_ (.A1_N(_10450_),
    .A2_N(_10451_),
    .B1(_10450_),
    .B2(_10451_),
    .X(_10452_));
 sky130_fd_sc_hd__a21oi_4 _26369_ (.A1(_10347_),
    .A2(_10349_),
    .B1(_10343_),
    .Y(_10453_));
 sky130_fd_sc_hd__o2bb2ai_2 _26370_ (.A1_N(_10452_),
    .A2_N(_10453_),
    .B1(_10452_),
    .B2(_10453_),
    .Y(_10454_));
 sky130_fd_sc_hd__o22a_1 _26371_ (.A1(_09918_),
    .A2(_10248_),
    .B1(_07680_),
    .B2(_06651_),
    .X(_10455_));
 sky130_fd_sc_hd__and4_1 _26372_ (.A(_10355_),
    .B(_07188_),
    .C(_13080_),
    .D(_07192_),
    .X(_10456_));
 sky130_fd_sc_hd__nor2_2 _26373_ (.A(_10455_),
    .B(_10456_),
    .Y(_10457_));
 sky130_fd_sc_hd__nor2_2 _26374_ (.A(_07532_),
    .B(_07178_),
    .Y(_10458_));
 sky130_fd_sc_hd__a2bb2o_2 _26375_ (.A1_N(_10457_),
    .A2_N(_10458_),
    .B1(_10457_),
    .B2(_10458_),
    .X(_10459_));
 sky130_fd_sc_hd__o2bb2ai_2 _26376_ (.A1_N(_10454_),
    .A2_N(_10459_),
    .B1(_10454_),
    .B2(_10459_),
    .Y(_10460_));
 sky130_fd_sc_hd__o22a_2 _26377_ (.A1(_10350_),
    .A2(_10351_),
    .B1(_10352_),
    .B2(_10360_),
    .X(_10461_));
 sky130_fd_sc_hd__o2bb2ai_2 _26378_ (.A1_N(_10460_),
    .A2_N(_10461_),
    .B1(_10460_),
    .B2(_10461_),
    .Y(_10462_));
 sky130_fd_sc_hd__a21oi_2 _26379_ (.A1(_10373_),
    .A2(_10376_),
    .B1(_10372_),
    .Y(_10463_));
 sky130_fd_sc_hd__a21oi_2 _26380_ (.A1(_10357_),
    .A2(_10359_),
    .B1(_10356_),
    .Y(_10464_));
 sky130_fd_sc_hd__buf_1 _26381_ (.A(_10229_),
    .X(_10465_));
 sky130_fd_sc_hd__o22a_1 _26382_ (.A1(_10465_),
    .A2(_07171_),
    .B1(_10368_),
    .B2(_07173_),
    .X(_10466_));
 sky130_fd_sc_hd__and4_2 _26383_ (.A(_10370_),
    .B(_07024_),
    .C(_10371_),
    .D(_07175_),
    .X(_10467_));
 sky130_fd_sc_hd__nor2_2 _26384_ (.A(_10466_),
    .B(_10467_),
    .Y(_10468_));
 sky130_fd_sc_hd__nor2_2 _26385_ (.A(_10374_),
    .B(_10327_),
    .Y(_10469_));
 sky130_fd_sc_hd__a2bb2o_1 _26386_ (.A1_N(_10468_),
    .A2_N(_10469_),
    .B1(_10468_),
    .B2(_10469_),
    .X(_10470_));
 sky130_fd_sc_hd__a2bb2o_1 _26387_ (.A1_N(_10464_),
    .A2_N(_10470_),
    .B1(_10464_),
    .B2(_10470_),
    .X(_10471_));
 sky130_fd_sc_hd__a2bb2o_2 _26388_ (.A1_N(_10463_),
    .A2_N(_10471_),
    .B1(_10463_),
    .B2(_10471_),
    .X(_10472_));
 sky130_fd_sc_hd__o2bb2ai_2 _26389_ (.A1_N(_10462_),
    .A2_N(_10472_),
    .B1(_10462_),
    .B2(_10472_),
    .Y(_10473_));
 sky130_fd_sc_hd__o22a_1 _26390_ (.A1(_10361_),
    .A2(_10362_),
    .B1(_10364_),
    .B2(_10379_),
    .X(_10474_));
 sky130_fd_sc_hd__o2bb2a_1 _26391_ (.A1_N(_10473_),
    .A2_N(_10474_),
    .B1(_10473_),
    .B2(_10474_),
    .X(_10475_));
 sky130_vsdinv _26392_ (.A(_10475_),
    .Y(_10476_));
 sky130_fd_sc_hd__o22a_1 _26393_ (.A1(_10336_),
    .A2(_10337_),
    .B1(_10325_),
    .B2(_10338_),
    .X(_10477_));
 sky130_fd_sc_hd__o22a_1 _26394_ (.A1(_10366_),
    .A2(_10377_),
    .B1(_10365_),
    .B2(_10378_),
    .X(_10478_));
 sky130_fd_sc_hd__buf_1 _26395_ (.A(_10008_),
    .X(_10479_));
 sky130_fd_sc_hd__buf_1 _26396_ (.A(_09258_),
    .X(_10480_));
 sky130_fd_sc_hd__o22a_1 _26397_ (.A1(_10479_),
    .A2(_10480_),
    .B1(_06392_),
    .B2(_07892_),
    .X(_10481_));
 sky130_fd_sc_hd__and4_2 _26398_ (.A(_13108_),
    .B(_08024_),
    .C(_13114_),
    .D(_13511_),
    .X(_10482_));
 sky130_fd_sc_hd__nor2_2 _26399_ (.A(_10481_),
    .B(_10482_),
    .Y(_10483_));
 sky130_fd_sc_hd__nor2_2 _26400_ (.A(_06287_),
    .B(_08500_),
    .Y(_10484_));
 sky130_fd_sc_hd__a2bb2o_1 _26401_ (.A1_N(_10483_),
    .A2_N(_10484_),
    .B1(_10483_),
    .B2(_10484_),
    .X(_10485_));
 sky130_fd_sc_hd__o22a_1 _26402_ (.A1(_10326_),
    .A2(_07737_),
    .B1(_10328_),
    .B2(_07881_),
    .X(_10486_));
 sky130_fd_sc_hd__and4_2 _26403_ (.A(_13099_),
    .B(_13530_),
    .C(_13104_),
    .D(_13525_),
    .X(_10487_));
 sky130_fd_sc_hd__nor2_2 _26404_ (.A(_10486_),
    .B(_10487_),
    .Y(_10488_));
 sky130_fd_sc_hd__buf_2 _26405_ (.A(_08027_),
    .X(_10489_));
 sky130_fd_sc_hd__nor2_2 _26406_ (.A(_10333_),
    .B(_10489_),
    .Y(_10490_));
 sky130_fd_sc_hd__a2bb2o_1 _26407_ (.A1_N(_10488_),
    .A2_N(_10490_),
    .B1(_10488_),
    .B2(_10490_),
    .X(_10491_));
 sky130_fd_sc_hd__a21oi_2 _26408_ (.A1(_10332_),
    .A2(_10335_),
    .B1(_10331_),
    .Y(_10492_));
 sky130_fd_sc_hd__a2bb2o_1 _26409_ (.A1_N(_10491_),
    .A2_N(_10492_),
    .B1(_10491_),
    .B2(_10492_),
    .X(_10493_));
 sky130_fd_sc_hd__a2bb2o_1 _26410_ (.A1_N(_10485_),
    .A2_N(_10493_),
    .B1(_10485_),
    .B2(_10493_),
    .X(_10494_));
 sky130_fd_sc_hd__a2bb2o_1 _26411_ (.A1_N(_10478_),
    .A2_N(_10494_),
    .B1(_10478_),
    .B2(_10494_),
    .X(_10495_));
 sky130_fd_sc_hd__a2bb2o_1 _26412_ (.A1_N(_10477_),
    .A2_N(_10495_),
    .B1(_10477_),
    .B2(_10495_),
    .X(_10496_));
 sky130_vsdinv _26413_ (.A(_10496_),
    .Y(_10497_));
 sky130_fd_sc_hd__a22o_1 _26414_ (.A1(_10476_),
    .A2(_10496_),
    .B1(_10475_),
    .B2(_10497_),
    .X(_10498_));
 sky130_fd_sc_hd__o22a_1 _26415_ (.A1(_10381_),
    .A2(_10382_),
    .B1(_10341_),
    .B2(_10383_),
    .X(_10499_));
 sky130_fd_sc_hd__a2bb2o_1 _26416_ (.A1_N(_10498_),
    .A2_N(_10499_),
    .B1(_10498_),
    .B2(_10499_),
    .X(_10500_));
 sky130_fd_sc_hd__a2bb2o_1 _26417_ (.A1_N(_10447_),
    .A2_N(_10500_),
    .B1(_10447_),
    .B2(_10500_),
    .X(_10501_));
 sky130_fd_sc_hd__o22a_1 _26418_ (.A1(_10384_),
    .A2(_10385_),
    .B1(_10317_),
    .B2(_10386_),
    .X(_10502_));
 sky130_fd_sc_hd__a2bb2o_1 _26419_ (.A1_N(_10501_),
    .A2_N(_10502_),
    .B1(_10501_),
    .B2(_10502_),
    .X(_10503_));
 sky130_fd_sc_hd__a2bb2o_1 _26420_ (.A1_N(_10423_),
    .A2_N(_10503_),
    .B1(_10423_),
    .B2(_10503_),
    .X(_10504_));
 sky130_fd_sc_hd__o22a_1 _26421_ (.A1(_10387_),
    .A2(_10388_),
    .B1(_10289_),
    .B2(_10389_),
    .X(_10505_));
 sky130_fd_sc_hd__a2bb2o_1 _26422_ (.A1_N(_10504_),
    .A2_N(_10505_),
    .B1(_10504_),
    .B2(_10505_),
    .X(_10506_));
 sky130_fd_sc_hd__a2bb2o_1 _26423_ (.A1_N(_10412_),
    .A2_N(_10506_),
    .B1(_10412_),
    .B2(_10506_),
    .X(_10507_));
 sky130_fd_sc_hd__o22a_1 _26424_ (.A1(_10390_),
    .A2(_10391_),
    .B1(_10280_),
    .B2(_10392_),
    .X(_10508_));
 sky130_fd_sc_hd__a2bb2o_1 _26425_ (.A1_N(_10507_),
    .A2_N(_10508_),
    .B1(_10507_),
    .B2(_10508_),
    .X(_10509_));
 sky130_fd_sc_hd__a2bb2o_1 _26426_ (.A1_N(_10279_),
    .A2_N(_10509_),
    .B1(_10279_),
    .B2(_10509_),
    .X(_10510_));
 sky130_fd_sc_hd__o22a_1 _26427_ (.A1(_10393_),
    .A2(_10394_),
    .B1(_10174_),
    .B2(_10395_),
    .X(_10511_));
 sky130_fd_sc_hd__or2_1 _26428_ (.A(_10510_),
    .B(_10511_),
    .X(_10512_));
 sky130_fd_sc_hd__a21bo_1 _26429_ (.A1(_10510_),
    .A2(_10511_),
    .B1_N(_10512_),
    .X(_10513_));
 sky130_fd_sc_hd__a2bb2o_1 _26430_ (.A1_N(_10408_),
    .A2_N(_10513_),
    .B1(_10408_),
    .B2(_10513_),
    .X(_02668_));
 sky130_fd_sc_hd__buf_1 _26431_ (.A(_10420_),
    .X(_10514_));
 sky130_fd_sc_hd__clkbuf_2 _26432_ (.A(_10514_),
    .X(_10515_));
 sky130_fd_sc_hd__o22a_1 _26433_ (.A1(_10416_),
    .A2(_10515_),
    .B1(_10415_),
    .B2(_10422_),
    .X(_10516_));
 sky130_fd_sc_hd__or2_1 _26434_ (.A(_10410_),
    .B(_10516_),
    .X(_10517_));
 sky130_fd_sc_hd__a21bo_1 _26435_ (.A1(_10275_),
    .A2(_10516_),
    .B1_N(_10517_),
    .X(_10518_));
 sky130_fd_sc_hd__o21a_1 _26436_ (.A1(_10176_),
    .A2(_10419_),
    .B1(_10414_),
    .X(_10519_));
 sky130_fd_sc_hd__buf_1 _26437_ (.A(_10519_),
    .X(_10520_));
 sky130_fd_sc_hd__buf_1 _26438_ (.A(_10420_),
    .X(_10521_));
 sky130_fd_sc_hd__o22a_1 _26439_ (.A1(_10426_),
    .A2(_10445_),
    .B1(_10425_),
    .B2(_10446_),
    .X(_10522_));
 sky130_fd_sc_hd__a2bb2o_1 _26440_ (.A1_N(_10521_),
    .A2_N(_10522_),
    .B1(_10521_),
    .B2(_10522_),
    .X(_10523_));
 sky130_fd_sc_hd__a2bb2o_1 _26441_ (.A1_N(_10520_),
    .A2_N(_10523_),
    .B1(_10520_),
    .B2(_10523_),
    .X(_10524_));
 sky130_fd_sc_hd__and4_4 _26442_ (.A(_10342_),
    .B(_06766_),
    .C(_13065_),
    .D(_13556_),
    .X(_10525_));
 sky130_fd_sc_hd__o22a_2 _26443_ (.A1(_10344_),
    .A2(_13561_),
    .B1(_10345_),
    .B2(_08557_),
    .X(_10526_));
 sky130_fd_sc_hd__nor2_2 _26444_ (.A(_10525_),
    .B(_10526_),
    .Y(_10527_));
 sky130_fd_sc_hd__nor2_4 _26445_ (.A(_10348_),
    .B(_06642_),
    .Y(_10528_));
 sky130_fd_sc_hd__a2bb2o_2 _26446_ (.A1_N(_10527_),
    .A2_N(_10528_),
    .B1(_10527_),
    .B2(_10528_),
    .X(_10529_));
 sky130_fd_sc_hd__a21oi_4 _26447_ (.A1(_10450_),
    .A2(_10451_),
    .B1(_10448_),
    .Y(_10530_));
 sky130_fd_sc_hd__o2bb2ai_1 _26448_ (.A1_N(_10529_),
    .A2_N(_10530_),
    .B1(_10529_),
    .B2(_10530_),
    .Y(_10531_));
 sky130_fd_sc_hd__o22a_1 _26449_ (.A1(_10353_),
    .A2(_06755_),
    .B1(_07680_),
    .B2(_06882_),
    .X(_10532_));
 sky130_fd_sc_hd__and4_2 _26450_ (.A(_10355_),
    .B(_07192_),
    .C(_13080_),
    .D(_06884_),
    .X(_10533_));
 sky130_fd_sc_hd__nor2_2 _26451_ (.A(_10532_),
    .B(_10533_),
    .Y(_10534_));
 sky130_fd_sc_hd__nor2_4 _26452_ (.A(_10358_),
    .B(_07321_),
    .Y(_10535_));
 sky130_fd_sc_hd__a2bb2o_2 _26453_ (.A1_N(_10534_),
    .A2_N(_10535_),
    .B1(_10534_),
    .B2(_10535_),
    .X(_10536_));
 sky130_fd_sc_hd__o2bb2ai_1 _26454_ (.A1_N(_10531_),
    .A2_N(_10536_),
    .B1(_10531_),
    .B2(_10536_),
    .Y(_10537_));
 sky130_fd_sc_hd__o22a_1 _26455_ (.A1(_10452_),
    .A2(_10453_),
    .B1(_10454_),
    .B2(_10459_),
    .X(_10538_));
 sky130_fd_sc_hd__o2bb2ai_1 _26456_ (.A1_N(_10537_),
    .A2_N(_10538_),
    .B1(_10537_),
    .B2(_10538_),
    .Y(_10539_));
 sky130_fd_sc_hd__a21oi_2 _26457_ (.A1(_10468_),
    .A2(_10469_),
    .B1(_10467_),
    .Y(_10540_));
 sky130_fd_sc_hd__a21oi_2 _26458_ (.A1(_10457_),
    .A2(_10458_),
    .B1(_10456_),
    .Y(_10541_));
 sky130_fd_sc_hd__o22a_1 _26459_ (.A1(_10229_),
    .A2(_07458_),
    .B1(_07269_),
    .B2(_07453_),
    .X(_10542_));
 sky130_fd_sc_hd__and4_1 _26460_ (.A(_13089_),
    .B(_13539_),
    .C(_13093_),
    .D(_13535_),
    .X(_10543_));
 sky130_fd_sc_hd__nor2_2 _26461_ (.A(_10542_),
    .B(_10543_),
    .Y(_10544_));
 sky130_fd_sc_hd__nor2_2 _26462_ (.A(_07075_),
    .B(_07737_),
    .Y(_10545_));
 sky130_fd_sc_hd__a2bb2o_1 _26463_ (.A1_N(_10544_),
    .A2_N(_10545_),
    .B1(_10544_),
    .B2(_10545_),
    .X(_10546_));
 sky130_fd_sc_hd__a2bb2o_1 _26464_ (.A1_N(_10541_),
    .A2_N(_10546_),
    .B1(_10541_),
    .B2(_10546_),
    .X(_10547_));
 sky130_fd_sc_hd__a2bb2o_1 _26465_ (.A1_N(_10540_),
    .A2_N(_10547_),
    .B1(_10540_),
    .B2(_10547_),
    .X(_10548_));
 sky130_fd_sc_hd__o2bb2ai_1 _26466_ (.A1_N(_10539_),
    .A2_N(_10548_),
    .B1(_10539_),
    .B2(_10548_),
    .Y(_10549_));
 sky130_fd_sc_hd__o22a_1 _26467_ (.A1(_10460_),
    .A2(_10461_),
    .B1(_10462_),
    .B2(_10472_),
    .X(_10550_));
 sky130_fd_sc_hd__o2bb2a_1 _26468_ (.A1_N(_10549_),
    .A2_N(_10550_),
    .B1(_10549_),
    .B2(_10550_),
    .X(_10551_));
 sky130_vsdinv _26469_ (.A(_10551_),
    .Y(_10552_));
 sky130_fd_sc_hd__o22a_1 _26470_ (.A1(_10491_),
    .A2(_10492_),
    .B1(_10485_),
    .B2(_10493_),
    .X(_10553_));
 sky130_fd_sc_hd__o22a_1 _26471_ (.A1(_10464_),
    .A2(_10470_),
    .B1(_10463_),
    .B2(_10471_),
    .X(_10554_));
 sky130_fd_sc_hd__o22a_1 _26472_ (.A1(_10479_),
    .A2(_08020_),
    .B1(_06392_),
    .B2(_08036_),
    .X(_10555_));
 sky130_fd_sc_hd__and4_1 _26473_ (.A(_13108_),
    .B(_08172_),
    .C(_13114_),
    .D(_13506_),
    .X(_10556_));
 sky130_fd_sc_hd__or2_1 _26474_ (.A(_10555_),
    .B(_10556_),
    .X(_10557_));
 sky130_vsdinv _26475_ (.A(_10557_),
    .Y(_10558_));
 sky130_fd_sc_hd__or2_1 _26476_ (.A(_11704_),
    .B(_08734_),
    .X(_10559_));
 sky130_fd_sc_hd__buf_1 _26477_ (.A(_10559_),
    .X(_10560_));
 sky130_fd_sc_hd__buf_1 _26478_ (.A(_10560_),
    .X(_10561_));
 sky130_fd_sc_hd__a32o_1 _26479_ (.A1(_10305_),
    .A2(\pcpi_mul.rs2[18] ),
    .A3(_10558_),
    .B1(_10557_),
    .B2(_10561_),
    .X(_10562_));
 sky130_fd_sc_hd__buf_1 _26480_ (.A(_10215_),
    .X(_10563_));
 sky130_fd_sc_hd__buf_1 _26481_ (.A(_10216_),
    .X(_10564_));
 sky130_fd_sc_hd__o22a_1 _26482_ (.A1(_10563_),
    .A2(_07881_),
    .B1(_10564_),
    .B2(_08027_),
    .X(_10565_));
 sky130_fd_sc_hd__and4_1 _26483_ (.A(_13099_),
    .B(_13525_),
    .C(_13104_),
    .D(_13521_),
    .X(_10566_));
 sky130_fd_sc_hd__nor2_2 _26484_ (.A(_10565_),
    .B(_10566_),
    .Y(_10567_));
 sky130_fd_sc_hd__clkbuf_2 _26485_ (.A(_10480_),
    .X(_10568_));
 sky130_fd_sc_hd__nor2_2 _26486_ (.A(_06690_),
    .B(_10568_),
    .Y(_10569_));
 sky130_fd_sc_hd__a2bb2o_1 _26487_ (.A1_N(_10567_),
    .A2_N(_10569_),
    .B1(_10567_),
    .B2(_10569_),
    .X(_10570_));
 sky130_fd_sc_hd__a21oi_2 _26488_ (.A1(_10488_),
    .A2(_10490_),
    .B1(_10487_),
    .Y(_10571_));
 sky130_fd_sc_hd__a2bb2o_1 _26489_ (.A1_N(_10570_),
    .A2_N(_10571_),
    .B1(_10570_),
    .B2(_10571_),
    .X(_10572_));
 sky130_fd_sc_hd__a2bb2o_1 _26490_ (.A1_N(_10562_),
    .A2_N(_10572_),
    .B1(_10562_),
    .B2(_10572_),
    .X(_10573_));
 sky130_fd_sc_hd__a2bb2o_1 _26491_ (.A1_N(_10554_),
    .A2_N(_10573_),
    .B1(_10554_),
    .B2(_10573_),
    .X(_10574_));
 sky130_fd_sc_hd__a2bb2o_1 _26492_ (.A1_N(_10553_),
    .A2_N(_10574_),
    .B1(_10553_),
    .B2(_10574_),
    .X(_10575_));
 sky130_vsdinv _26493_ (.A(_10575_),
    .Y(_10576_));
 sky130_fd_sc_hd__a22o_1 _26494_ (.A1(_10552_),
    .A2(_10575_),
    .B1(_10551_),
    .B2(_10576_),
    .X(_10577_));
 sky130_fd_sc_hd__o22a_1 _26495_ (.A1(_10473_),
    .A2(_10474_),
    .B1(_10476_),
    .B2(_10496_),
    .X(_10578_));
 sky130_fd_sc_hd__a2bb2o_1 _26496_ (.A1_N(_10577_),
    .A2_N(_10578_),
    .B1(_10577_),
    .B2(_10578_),
    .X(_10579_));
 sky130_fd_sc_hd__o22a_1 _26497_ (.A1(_10441_),
    .A2(_10442_),
    .B1(_10424_),
    .B2(_10444_),
    .X(_10580_));
 sky130_fd_sc_hd__o22a_1 _26498_ (.A1(_10478_),
    .A2(_10494_),
    .B1(_10477_),
    .B2(_10495_),
    .X(_10581_));
 sky130_fd_sc_hd__buf_1 _26499_ (.A(_10435_),
    .X(_10582_));
 sky130_fd_sc_hd__a21oi_4 _26500_ (.A1(_10483_),
    .A2(_10484_),
    .B1(_10482_),
    .Y(_10583_));
 sky130_fd_sc_hd__a2bb2o_1 _26501_ (.A1_N(_10582_),
    .A2_N(_10583_),
    .B1(_10582_),
    .B2(_10583_),
    .X(_10584_));
 sky130_fd_sc_hd__o21a_1 _26502_ (.A1(_10197_),
    .A2(_10434_),
    .B1(_10430_),
    .X(_10585_));
 sky130_fd_sc_hd__o2bb2a_1 _26503_ (.A1_N(_10584_),
    .A2_N(_10585_),
    .B1(_10584_),
    .B2(_10585_),
    .X(_10586_));
 sky130_vsdinv _26504_ (.A(_10586_),
    .Y(_10587_));
 sky130_fd_sc_hd__buf_1 _26505_ (.A(_10435_),
    .X(_10588_));
 sky130_fd_sc_hd__o22a_1 _26506_ (.A1(_10428_),
    .A2(_10588_),
    .B1(_10438_),
    .B2(_10439_),
    .X(_10589_));
 sky130_vsdinv _26507_ (.A(_10589_),
    .Y(_10590_));
 sky130_fd_sc_hd__a22o_1 _26508_ (.A1(_10587_),
    .A2(_10589_),
    .B1(_10586_),
    .B2(_10590_),
    .X(_10591_));
 sky130_fd_sc_hd__a2bb2o_1 _26509_ (.A1_N(_10427_),
    .A2_N(_10591_),
    .B1(_10427_),
    .B2(_10591_),
    .X(_10592_));
 sky130_fd_sc_hd__a2bb2o_1 _26510_ (.A1_N(_10581_),
    .A2_N(_10592_),
    .B1(_10581_),
    .B2(_10592_),
    .X(_10593_));
 sky130_fd_sc_hd__a2bb2o_1 _26511_ (.A1_N(_10580_),
    .A2_N(_10593_),
    .B1(_10580_),
    .B2(_10593_),
    .X(_10594_));
 sky130_fd_sc_hd__a2bb2o_1 _26512_ (.A1_N(_10579_),
    .A2_N(_10594_),
    .B1(_10579_),
    .B2(_10594_),
    .X(_10595_));
 sky130_fd_sc_hd__o22a_1 _26513_ (.A1(_10498_),
    .A2(_10499_),
    .B1(_10447_),
    .B2(_10500_),
    .X(_10596_));
 sky130_fd_sc_hd__a2bb2o_1 _26514_ (.A1_N(_10595_),
    .A2_N(_10596_),
    .B1(_10595_),
    .B2(_10596_),
    .X(_10597_));
 sky130_fd_sc_hd__a2bb2o_1 _26515_ (.A1_N(_10524_),
    .A2_N(_10597_),
    .B1(_10524_),
    .B2(_10597_),
    .X(_10598_));
 sky130_fd_sc_hd__o22a_1 _26516_ (.A1(_10501_),
    .A2(_10502_),
    .B1(_10423_),
    .B2(_10503_),
    .X(_10599_));
 sky130_fd_sc_hd__a2bb2o_1 _26517_ (.A1_N(_10598_),
    .A2_N(_10599_),
    .B1(_10598_),
    .B2(_10599_),
    .X(_10600_));
 sky130_fd_sc_hd__a2bb2o_1 _26518_ (.A1_N(_10518_),
    .A2_N(_10600_),
    .B1(_10518_),
    .B2(_10600_),
    .X(_10601_));
 sky130_fd_sc_hd__o22a_1 _26519_ (.A1(_10504_),
    .A2(_10505_),
    .B1(_10412_),
    .B2(_10506_),
    .X(_10602_));
 sky130_fd_sc_hd__a2bb2o_1 _26520_ (.A1_N(_10601_),
    .A2_N(_10602_),
    .B1(_10601_),
    .B2(_10602_),
    .X(_10603_));
 sky130_fd_sc_hd__a2bb2o_1 _26521_ (.A1_N(_10411_),
    .A2_N(_10603_),
    .B1(_10411_),
    .B2(_10603_),
    .X(_10604_));
 sky130_fd_sc_hd__o22a_1 _26522_ (.A1(_10507_),
    .A2(_10508_),
    .B1(_10279_),
    .B2(_10509_),
    .X(_10605_));
 sky130_fd_sc_hd__or2_1 _26523_ (.A(_10604_),
    .B(_10605_),
    .X(_10606_));
 sky130_fd_sc_hd__a21bo_1 _26524_ (.A1(_10604_),
    .A2(_10605_),
    .B1_N(_10606_),
    .X(_10607_));
 sky130_fd_sc_hd__a22o_1 _26525_ (.A1(_10510_),
    .A2(_10511_),
    .B1(_10398_),
    .B2(_10512_),
    .X(_10608_));
 sky130_fd_sc_hd__o31a_1 _26526_ (.A1(_10400_),
    .A2(_10513_),
    .A3(_10407_),
    .B1(_10608_),
    .X(_10609_));
 sky130_fd_sc_hd__a2bb2oi_1 _26527_ (.A1_N(_10607_),
    .A2_N(_10609_),
    .B1(_10607_),
    .B2(_10609_),
    .Y(_02669_));
 sky130_fd_sc_hd__buf_1 _26528_ (.A(_10521_),
    .X(_10610_));
 sky130_fd_sc_hd__buf_1 _26529_ (.A(_10519_),
    .X(_10611_));
 sky130_fd_sc_hd__o22a_1 _26530_ (.A1(_10610_),
    .A2(_10522_),
    .B1(_10611_),
    .B2(_10523_),
    .X(_10612_));
 sky130_fd_sc_hd__or2_1 _26531_ (.A(_10278_),
    .B(_10612_),
    .X(_10613_));
 sky130_fd_sc_hd__a21bo_1 _26532_ (.A1(_10276_),
    .A2(_10612_),
    .B1_N(_10613_),
    .X(_10614_));
 sky130_fd_sc_hd__and4_2 _26533_ (.A(_10342_),
    .B(_06566_),
    .C(_13066_),
    .D(_07188_),
    .X(_10615_));
 sky130_fd_sc_hd__clkbuf_2 _26534_ (.A(_10345_),
    .X(_10616_));
 sky130_fd_sc_hd__o22a_2 _26535_ (.A1(_10344_),
    .A2(_13556_),
    .B1(_10616_),
    .B2(_10248_),
    .X(_10617_));
 sky130_fd_sc_hd__nor2_2 _26536_ (.A(_10615_),
    .B(_10617_),
    .Y(_10618_));
 sky130_fd_sc_hd__nor2_4 _26537_ (.A(_10348_),
    .B(_06879_),
    .Y(_10619_));
 sky130_fd_sc_hd__a2bb2o_2 _26538_ (.A1_N(_10618_),
    .A2_N(_10619_),
    .B1(_10618_),
    .B2(_10619_),
    .X(_10620_));
 sky130_fd_sc_hd__a21oi_4 _26539_ (.A1(_10527_),
    .A2(_10528_),
    .B1(_10525_),
    .Y(_10621_));
 sky130_fd_sc_hd__o2bb2ai_2 _26540_ (.A1_N(_10620_),
    .A2_N(_10621_),
    .B1(_10620_),
    .B2(_10621_),
    .Y(_10622_));
 sky130_fd_sc_hd__buf_1 _26541_ (.A(_09919_),
    .X(_10623_));
 sky130_fd_sc_hd__o22a_1 _26542_ (.A1(_10353_),
    .A2(_06882_),
    .B1(_10623_),
    .B2(_07020_),
    .X(_10624_));
 sky130_fd_sc_hd__and4_2 _26543_ (.A(_10355_),
    .B(_13547_),
    .C(_13081_),
    .D(_07024_),
    .X(_10625_));
 sky130_fd_sc_hd__nor2_2 _26544_ (.A(_10624_),
    .B(_10625_),
    .Y(_10626_));
 sky130_fd_sc_hd__nor2_4 _26545_ (.A(_10358_),
    .B(_10375_),
    .Y(_10627_));
 sky130_fd_sc_hd__a2bb2o_2 _26546_ (.A1_N(_10626_),
    .A2_N(_10627_),
    .B1(_10626_),
    .B2(_10627_),
    .X(_10628_));
 sky130_fd_sc_hd__o2bb2ai_2 _26547_ (.A1_N(_10622_),
    .A2_N(_10628_),
    .B1(_10622_),
    .B2(_10628_),
    .Y(_10629_));
 sky130_fd_sc_hd__o22a_1 _26548_ (.A1(_10529_),
    .A2(_10530_),
    .B1(_10531_),
    .B2(_10536_),
    .X(_10630_));
 sky130_fd_sc_hd__o2bb2ai_1 _26549_ (.A1_N(_10629_),
    .A2_N(_10630_),
    .B1(_10629_),
    .B2(_10630_),
    .Y(_10631_));
 sky130_fd_sc_hd__a21oi_2 _26550_ (.A1(_10544_),
    .A2(_10545_),
    .B1(_10543_),
    .Y(_10632_));
 sky130_fd_sc_hd__a21oi_4 _26551_ (.A1(_10534_),
    .A2(_10535_),
    .B1(_10533_),
    .Y(_10633_));
 sky130_fd_sc_hd__o22a_1 _26552_ (.A1(_10465_),
    .A2(_09783_),
    .B1(_07269_),
    .B2(_09895_),
    .X(_10634_));
 sky130_fd_sc_hd__and4_2 _26553_ (.A(_13089_),
    .B(_13535_),
    .C(_13093_),
    .D(_07450_),
    .X(_10635_));
 sky130_fd_sc_hd__nor2_2 _26554_ (.A(_10634_),
    .B(_10635_),
    .Y(_10636_));
 sky130_fd_sc_hd__nor2_2 _26555_ (.A(_07075_),
    .B(_07881_),
    .Y(_10637_));
 sky130_fd_sc_hd__a2bb2o_1 _26556_ (.A1_N(_10636_),
    .A2_N(_10637_),
    .B1(_10636_),
    .B2(_10637_),
    .X(_10638_));
 sky130_fd_sc_hd__a2bb2o_1 _26557_ (.A1_N(_10633_),
    .A2_N(_10638_),
    .B1(_10633_),
    .B2(_10638_),
    .X(_10639_));
 sky130_fd_sc_hd__a2bb2o_1 _26558_ (.A1_N(_10632_),
    .A2_N(_10639_),
    .B1(_10632_),
    .B2(_10639_),
    .X(_10640_));
 sky130_fd_sc_hd__o2bb2ai_1 _26559_ (.A1_N(_10631_),
    .A2_N(_10640_),
    .B1(_10631_),
    .B2(_10640_),
    .Y(_10641_));
 sky130_fd_sc_hd__o22a_1 _26560_ (.A1(_10537_),
    .A2(_10538_),
    .B1(_10539_),
    .B2(_10548_),
    .X(_10642_));
 sky130_fd_sc_hd__o2bb2a_1 _26561_ (.A1_N(_10641_),
    .A2_N(_10642_),
    .B1(_10641_),
    .B2(_10642_),
    .X(_10643_));
 sky130_vsdinv _26562_ (.A(_10643_),
    .Y(_10644_));
 sky130_fd_sc_hd__o22a_1 _26563_ (.A1(_10570_),
    .A2(_10571_),
    .B1(_10562_),
    .B2(_10572_),
    .X(_10645_));
 sky130_fd_sc_hd__o22a_1 _26564_ (.A1(_10541_),
    .A2(_10546_),
    .B1(_10540_),
    .B2(_10547_),
    .X(_10646_));
 sky130_fd_sc_hd__nor2_1 _26565_ (.A(_10479_),
    .B(_08499_),
    .Y(_10647_));
 sky130_fd_sc_hd__or2_2 _26566_ (.A(_08660_),
    .B(_08736_),
    .X(_10648_));
 sky130_vsdinv _26567_ (.A(_10648_),
    .Y(_10649_));
 sky130_fd_sc_hd__a2bb2o_1 _26568_ (.A1_N(_10647_),
    .A2_N(_10649_),
    .B1(_10647_),
    .B2(_10649_),
    .X(_10650_));
 sky130_fd_sc_hd__a2bb2o_1 _26569_ (.A1_N(_10561_),
    .A2_N(_10650_),
    .B1(_10561_),
    .B2(_10650_),
    .X(_10651_));
 sky130_fd_sc_hd__o22a_1 _26570_ (.A1(_10563_),
    .A2(_07871_),
    .B1(_10564_),
    .B2(_10480_),
    .X(_10652_));
 sky130_fd_sc_hd__buf_1 _26571_ (.A(_09554_),
    .X(_10653_));
 sky130_fd_sc_hd__buf_1 _26572_ (.A(_09555_),
    .X(_10654_));
 sky130_fd_sc_hd__and4_2 _26573_ (.A(_10653_),
    .B(_07878_),
    .C(_10654_),
    .D(_08024_),
    .X(_10655_));
 sky130_fd_sc_hd__nor2_2 _26574_ (.A(_10652_),
    .B(_10655_),
    .Y(_10656_));
 sky130_fd_sc_hd__nor2_2 _26575_ (.A(_06690_),
    .B(_10323_),
    .Y(_10657_));
 sky130_fd_sc_hd__a2bb2o_1 _26576_ (.A1_N(_10656_),
    .A2_N(_10657_),
    .B1(_10656_),
    .B2(_10657_),
    .X(_10658_));
 sky130_fd_sc_hd__a21oi_2 _26577_ (.A1(_10567_),
    .A2(_10569_),
    .B1(_10566_),
    .Y(_10659_));
 sky130_fd_sc_hd__a2bb2o_1 _26578_ (.A1_N(_10658_),
    .A2_N(_10659_),
    .B1(_10658_),
    .B2(_10659_),
    .X(_10660_));
 sky130_fd_sc_hd__a2bb2o_1 _26579_ (.A1_N(_10651_),
    .A2_N(_10660_),
    .B1(_10651_),
    .B2(_10660_),
    .X(_10661_));
 sky130_fd_sc_hd__a2bb2o_1 _26580_ (.A1_N(_10646_),
    .A2_N(_10661_),
    .B1(_10646_),
    .B2(_10661_),
    .X(_10662_));
 sky130_fd_sc_hd__a2bb2o_1 _26581_ (.A1_N(_10645_),
    .A2_N(_10662_),
    .B1(_10645_),
    .B2(_10662_),
    .X(_10663_));
 sky130_vsdinv _26582_ (.A(_10663_),
    .Y(_10664_));
 sky130_fd_sc_hd__a22o_1 _26583_ (.A1(_10644_),
    .A2(_10663_),
    .B1(_10643_),
    .B2(_10664_),
    .X(_10665_));
 sky130_fd_sc_hd__o22a_1 _26584_ (.A1(_10549_),
    .A2(_10550_),
    .B1(_10552_),
    .B2(_10575_),
    .X(_10666_));
 sky130_fd_sc_hd__a2bb2o_1 _26585_ (.A1_N(_10665_),
    .A2_N(_10666_),
    .B1(_10665_),
    .B2(_10666_),
    .X(_10667_));
 sky130_fd_sc_hd__o22a_1 _26586_ (.A1(_10587_),
    .A2(_10589_),
    .B1(_10424_),
    .B2(_10591_),
    .X(_10668_));
 sky130_fd_sc_hd__o22a_1 _26587_ (.A1(_10554_),
    .A2(_10573_),
    .B1(_10553_),
    .B2(_10574_),
    .X(_10669_));
 sky130_fd_sc_hd__buf_1 _26588_ (.A(_10585_),
    .X(_10670_));
 sky130_fd_sc_hd__o21ba_1 _26589_ (.A1(_10557_),
    .A2(_10560_),
    .B1_N(_10556_),
    .X(_10671_));
 sky130_fd_sc_hd__a2bb2o_1 _26590_ (.A1_N(_10588_),
    .A2_N(_10671_),
    .B1(_10582_),
    .B2(_10671_),
    .X(_10672_));
 sky130_fd_sc_hd__a2bb2o_1 _26591_ (.A1_N(_10670_),
    .A2_N(_10672_),
    .B1(_10670_),
    .B2(_10672_),
    .X(_10673_));
 sky130_fd_sc_hd__o22a_1 _26592_ (.A1(_10588_),
    .A2(_10583_),
    .B1(_10584_),
    .B2(_10670_),
    .X(_10674_));
 sky130_fd_sc_hd__o2bb2ai_1 _26593_ (.A1_N(_10673_),
    .A2_N(_10674_),
    .B1(_10673_),
    .B2(_10674_),
    .Y(_10675_));
 sky130_fd_sc_hd__a2bb2o_1 _26594_ (.A1_N(_10295_),
    .A2_N(_10675_),
    .B1(_10295_),
    .B2(_10675_),
    .X(_10676_));
 sky130_fd_sc_hd__a2bb2o_1 _26595_ (.A1_N(_10669_),
    .A2_N(_10676_),
    .B1(_10669_),
    .B2(_10676_),
    .X(_10677_));
 sky130_fd_sc_hd__a2bb2o_1 _26596_ (.A1_N(_10668_),
    .A2_N(_10677_),
    .B1(_10668_),
    .B2(_10677_),
    .X(_10678_));
 sky130_fd_sc_hd__a2bb2o_1 _26597_ (.A1_N(_10667_),
    .A2_N(_10678_),
    .B1(_10667_),
    .B2(_10678_),
    .X(_10679_));
 sky130_fd_sc_hd__o22a_1 _26598_ (.A1(_10577_),
    .A2(_10578_),
    .B1(_10579_),
    .B2(_10594_),
    .X(_10680_));
 sky130_fd_sc_hd__a2bb2o_1 _26599_ (.A1_N(_10679_),
    .A2_N(_10680_),
    .B1(_10679_),
    .B2(_10680_),
    .X(_10681_));
 sky130_fd_sc_hd__buf_1 _26600_ (.A(_10519_),
    .X(_10682_));
 sky130_fd_sc_hd__buf_1 _26601_ (.A(_10682_),
    .X(_10683_));
 sky130_fd_sc_hd__buf_1 _26602_ (.A(_10514_),
    .X(_10684_));
 sky130_fd_sc_hd__o22a_1 _26603_ (.A1(_10581_),
    .A2(_10592_),
    .B1(_10580_),
    .B2(_10593_),
    .X(_10685_));
 sky130_fd_sc_hd__a2bb2o_1 _26604_ (.A1_N(_10684_),
    .A2_N(_10685_),
    .B1(_10684_),
    .B2(_10685_),
    .X(_10686_));
 sky130_fd_sc_hd__a2bb2o_1 _26605_ (.A1_N(_10683_),
    .A2_N(_10686_),
    .B1(_10683_),
    .B2(_10686_),
    .X(_10687_));
 sky130_fd_sc_hd__a2bb2o_1 _26606_ (.A1_N(_10681_),
    .A2_N(_10687_),
    .B1(_10681_),
    .B2(_10687_),
    .X(_10688_));
 sky130_fd_sc_hd__o22a_1 _26607_ (.A1(_10595_),
    .A2(_10596_),
    .B1(_10524_),
    .B2(_10597_),
    .X(_10689_));
 sky130_fd_sc_hd__a2bb2o_1 _26608_ (.A1_N(_10688_),
    .A2_N(_10689_),
    .B1(_10688_),
    .B2(_10689_),
    .X(_10690_));
 sky130_fd_sc_hd__a2bb2o_1 _26609_ (.A1_N(_10614_),
    .A2_N(_10690_),
    .B1(_10614_),
    .B2(_10690_),
    .X(_10691_));
 sky130_fd_sc_hd__o22a_1 _26610_ (.A1(_10598_),
    .A2(_10599_),
    .B1(_10518_),
    .B2(_10600_),
    .X(_10692_));
 sky130_fd_sc_hd__a2bb2o_1 _26611_ (.A1_N(_10691_),
    .A2_N(_10692_),
    .B1(_10691_),
    .B2(_10692_),
    .X(_10693_));
 sky130_fd_sc_hd__a2bb2o_1 _26612_ (.A1_N(_10517_),
    .A2_N(_10693_),
    .B1(_10517_),
    .B2(_10693_),
    .X(_10694_));
 sky130_fd_sc_hd__o22a_1 _26613_ (.A1(_10601_),
    .A2(_10602_),
    .B1(_10411_),
    .B2(_10603_),
    .X(_10695_));
 sky130_fd_sc_hd__and2_1 _26614_ (.A(_10694_),
    .B(_10695_),
    .X(_10696_));
 sky130_fd_sc_hd__or2_1 _26615_ (.A(_10694_),
    .B(_10695_),
    .X(_10697_));
 sky130_fd_sc_hd__or2b_1 _26616_ (.A(_10696_),
    .B_N(_10697_),
    .X(_10698_));
 sky130_fd_sc_hd__o21ai_1 _26617_ (.A1(_10607_),
    .A2(_10609_),
    .B1(_10606_),
    .Y(_10699_));
 sky130_fd_sc_hd__a2bb2o_1 _26618_ (.A1_N(_10698_),
    .A2_N(_10699_),
    .B1(_10698_),
    .B2(_10699_),
    .X(_02670_));
 sky130_fd_sc_hd__and4_2 _26619_ (.A(_10342_),
    .B(_10248_),
    .C(_13066_),
    .D(_07192_),
    .X(_10700_));
 sky130_fd_sc_hd__o22a_1 _26620_ (.A1(_11719_),
    .A2(_07188_),
    .B1(_10616_),
    .B2(_06651_),
    .X(_10701_));
 sky130_fd_sc_hd__nor2_2 _26621_ (.A(_10700_),
    .B(_10701_),
    .Y(_10702_));
 sky130_fd_sc_hd__nor2_4 _26622_ (.A(_10348_),
    .B(_07178_),
    .Y(_10703_));
 sky130_fd_sc_hd__a2bb2o_2 _26623_ (.A1_N(_10702_),
    .A2_N(_10703_),
    .B1(_10702_),
    .B2(_10703_),
    .X(_10704_));
 sky130_fd_sc_hd__a21oi_4 _26624_ (.A1(_10618_),
    .A2(_10619_),
    .B1(_10615_),
    .Y(_10705_));
 sky130_fd_sc_hd__o2bb2ai_4 _26625_ (.A1_N(_10704_),
    .A2_N(_10705_),
    .B1(_10704_),
    .B2(_10705_),
    .Y(_10706_));
 sky130_fd_sc_hd__o22a_1 _26626_ (.A1(_10353_),
    .A2(_07020_),
    .B1(_10623_),
    .B2(_07459_),
    .X(_10707_));
 sky130_fd_sc_hd__and4_2 _26627_ (.A(_13075_),
    .B(_13543_),
    .C(_13081_),
    .D(_13540_),
    .X(_10708_));
 sky130_fd_sc_hd__nor2_2 _26628_ (.A(_10707_),
    .B(_10708_),
    .Y(_10709_));
 sky130_fd_sc_hd__buf_2 _26629_ (.A(_07198_),
    .X(_10710_));
 sky130_fd_sc_hd__nor2_4 _26630_ (.A(_10358_),
    .B(_10710_),
    .Y(_10711_));
 sky130_fd_sc_hd__a2bb2o_2 _26631_ (.A1_N(_10709_),
    .A2_N(_10711_),
    .B1(_10709_),
    .B2(_10711_),
    .X(_10712_));
 sky130_fd_sc_hd__o2bb2ai_4 _26632_ (.A1_N(_10706_),
    .A2_N(_10712_),
    .B1(_10706_),
    .B2(_10712_),
    .Y(_10713_));
 sky130_fd_sc_hd__o22a_2 _26633_ (.A1(_10620_),
    .A2(_10621_),
    .B1(_10622_),
    .B2(_10628_),
    .X(_10714_));
 sky130_fd_sc_hd__o2bb2ai_2 _26634_ (.A1_N(_10713_),
    .A2_N(_10714_),
    .B1(_10713_),
    .B2(_10714_),
    .Y(_10715_));
 sky130_fd_sc_hd__a21oi_2 _26635_ (.A1(_10636_),
    .A2(_10637_),
    .B1(_10635_),
    .Y(_10716_));
 sky130_fd_sc_hd__a21oi_4 _26636_ (.A1(_10626_),
    .A2(_10627_),
    .B1(_10625_),
    .Y(_10717_));
 sky130_fd_sc_hd__o22a_1 _26637_ (.A1(_10465_),
    .A2(_07737_),
    .B1(_07269_),
    .B2(_10012_),
    .X(_10718_));
 sky130_fd_sc_hd__and4_1 _26638_ (.A(_13089_),
    .B(_07450_),
    .C(_10371_),
    .D(_07588_),
    .X(_10719_));
 sky130_fd_sc_hd__nor2_2 _26639_ (.A(_10718_),
    .B(_10719_),
    .Y(_10720_));
 sky130_fd_sc_hd__nor2_2 _26640_ (.A(_07075_),
    .B(_08027_),
    .Y(_10721_));
 sky130_fd_sc_hd__a2bb2o_1 _26641_ (.A1_N(_10720_),
    .A2_N(_10721_),
    .B1(_10720_),
    .B2(_10721_),
    .X(_10722_));
 sky130_fd_sc_hd__a2bb2o_1 _26642_ (.A1_N(_10717_),
    .A2_N(_10722_),
    .B1(_10717_),
    .B2(_10722_),
    .X(_10723_));
 sky130_fd_sc_hd__a2bb2o_2 _26643_ (.A1_N(_10716_),
    .A2_N(_10723_),
    .B1(_10716_),
    .B2(_10723_),
    .X(_10724_));
 sky130_fd_sc_hd__o2bb2ai_2 _26644_ (.A1_N(_10715_),
    .A2_N(_10724_),
    .B1(_10715_),
    .B2(_10724_),
    .Y(_10725_));
 sky130_fd_sc_hd__o22a_1 _26645_ (.A1(_10629_),
    .A2(_10630_),
    .B1(_10631_),
    .B2(_10640_),
    .X(_10726_));
 sky130_fd_sc_hd__o2bb2ai_1 _26646_ (.A1_N(_10725_),
    .A2_N(_10726_),
    .B1(_10725_),
    .B2(_10726_),
    .Y(_10727_));
 sky130_fd_sc_hd__o22a_1 _26647_ (.A1(_10658_),
    .A2(_10659_),
    .B1(_10651_),
    .B2(_10660_),
    .X(_10728_));
 sky130_fd_sc_hd__o22a_1 _26648_ (.A1(_10633_),
    .A2(_10638_),
    .B1(_10632_),
    .B2(_10639_),
    .X(_10729_));
 sky130_fd_sc_hd__or2_1 _26649_ (.A(_11703_),
    .B(_09545_),
    .X(_10730_));
 sky130_fd_sc_hd__a32o_1 _26650_ (.A1(_08816_),
    .A2(_13108_),
    .A3(_10649_),
    .B1(_10648_),
    .B2(_10730_),
    .X(_10731_));
 sky130_fd_sc_hd__a2bb2o_2 _26651_ (.A1_N(_10560_),
    .A2_N(_10731_),
    .B1(_10560_),
    .B2(_10731_),
    .X(_10732_));
 sky130_fd_sc_hd__buf_1 _26652_ (.A(_10732_),
    .X(_10733_));
 sky130_fd_sc_hd__o22a_1 _26653_ (.A1(_10215_),
    .A2(_09258_),
    .B1(_10216_),
    .B2(_07891_),
    .X(_10734_));
 sky130_fd_sc_hd__and4_1 _26654_ (.A(_10653_),
    .B(_13516_),
    .C(_10654_),
    .D(_08172_),
    .X(_10735_));
 sky130_fd_sc_hd__nor2_1 _26655_ (.A(_10734_),
    .B(_10735_),
    .Y(_10736_));
 sky130_fd_sc_hd__nor2_1 _26656_ (.A(_06690_),
    .B(_08500_),
    .Y(_10737_));
 sky130_fd_sc_hd__a2bb2o_1 _26657_ (.A1_N(_10736_),
    .A2_N(_10737_),
    .B1(_10736_),
    .B2(_10737_),
    .X(_10738_));
 sky130_fd_sc_hd__a21oi_4 _26658_ (.A1(_10656_),
    .A2(_10657_),
    .B1(_10655_),
    .Y(_10739_));
 sky130_fd_sc_hd__a2bb2o_1 _26659_ (.A1_N(_10738_),
    .A2_N(_10739_),
    .B1(_10738_),
    .B2(_10739_),
    .X(_10740_));
 sky130_fd_sc_hd__a2bb2o_1 _26660_ (.A1_N(_10733_),
    .A2_N(_10740_),
    .B1(_10733_),
    .B2(_10740_),
    .X(_10741_));
 sky130_fd_sc_hd__a2bb2o_1 _26661_ (.A1_N(_10729_),
    .A2_N(_10741_),
    .B1(_10729_),
    .B2(_10741_),
    .X(_10742_));
 sky130_fd_sc_hd__a2bb2o_1 _26662_ (.A1_N(_10728_),
    .A2_N(_10742_),
    .B1(_10728_),
    .B2(_10742_),
    .X(_10743_));
 sky130_fd_sc_hd__o2bb2ai_1 _26663_ (.A1_N(_10727_),
    .A2_N(_10743_),
    .B1(_10727_),
    .B2(_10743_),
    .Y(_10744_));
 sky130_fd_sc_hd__o22a_1 _26664_ (.A1(_10641_),
    .A2(_10642_),
    .B1(_10644_),
    .B2(_10663_),
    .X(_10745_));
 sky130_fd_sc_hd__o2bb2a_1 _26665_ (.A1_N(_10744_),
    .A2_N(_10745_),
    .B1(_10744_),
    .B2(_10745_),
    .X(_10746_));
 sky130_vsdinv _26666_ (.A(_10746_),
    .Y(_10747_));
 sky130_fd_sc_hd__o22a_1 _26667_ (.A1(_10673_),
    .A2(_10674_),
    .B1(_10291_),
    .B2(_10675_),
    .X(_10748_));
 sky130_fd_sc_hd__o22a_1 _26668_ (.A1(_10646_),
    .A2(_10661_),
    .B1(_10645_),
    .B2(_10662_),
    .X(_10749_));
 sky130_fd_sc_hd__o22a_1 _26669_ (.A1(_10588_),
    .A2(_10671_),
    .B1(_10670_),
    .B2(_10672_),
    .X(_10750_));
 sky130_fd_sc_hd__buf_2 _26670_ (.A(_08499_),
    .X(_10751_));
 sky130_fd_sc_hd__o32a_1 _26671_ (.A1(_10479_),
    .A2(_10751_),
    .A3(_10648_),
    .B1(_10561_),
    .B2(_10650_),
    .X(_10752_));
 sky130_vsdinv _26672_ (.A(_10752_),
    .Y(_10753_));
 sky130_fd_sc_hd__nor2_1 _26673_ (.A(_10199_),
    .B(_10432_),
    .Y(_10754_));
 sky130_fd_sc_hd__a21oi_1 _26674_ (.A1(_13126_),
    .A2(_10433_),
    .B1(_10754_),
    .Y(_10755_));
 sky130_fd_sc_hd__a2bb2o_1 _26675_ (.A1_N(_10753_),
    .A2_N(_10755_),
    .B1(_10753_),
    .B2(_10755_),
    .X(_10756_));
 sky130_fd_sc_hd__o2bb2ai_1 _26676_ (.A1_N(_10750_),
    .A2_N(_10756_),
    .B1(_10750_),
    .B2(_10756_),
    .Y(_10757_));
 sky130_fd_sc_hd__a2bb2o_1 _26677_ (.A1_N(_10314_),
    .A2_N(_10757_),
    .B1(_10314_),
    .B2(_10757_),
    .X(_10758_));
 sky130_fd_sc_hd__a2bb2o_1 _26678_ (.A1_N(_10749_),
    .A2_N(_10758_),
    .B1(_10749_),
    .B2(_10758_),
    .X(_10759_));
 sky130_fd_sc_hd__a2bb2o_1 _26679_ (.A1_N(_10748_),
    .A2_N(_10759_),
    .B1(_10748_),
    .B2(_10759_),
    .X(_10760_));
 sky130_vsdinv _26680_ (.A(_10760_),
    .Y(_10761_));
 sky130_fd_sc_hd__a22o_1 _26681_ (.A1(_10747_),
    .A2(_10760_),
    .B1(_10746_),
    .B2(_10761_),
    .X(_10762_));
 sky130_fd_sc_hd__o22a_1 _26682_ (.A1(_10665_),
    .A2(_10666_),
    .B1(_10667_),
    .B2(_10678_),
    .X(_10763_));
 sky130_fd_sc_hd__a2bb2o_1 _26683_ (.A1_N(_10762_),
    .A2_N(_10763_),
    .B1(_10762_),
    .B2(_10763_),
    .X(_10764_));
 sky130_fd_sc_hd__buf_1 _26684_ (.A(_10682_),
    .X(_10765_));
 sky130_fd_sc_hd__o22a_1 _26685_ (.A1(_10669_),
    .A2(_10676_),
    .B1(_10668_),
    .B2(_10677_),
    .X(_10766_));
 sky130_fd_sc_hd__a2bb2o_1 _26686_ (.A1_N(_10421_),
    .A2_N(_10766_),
    .B1(_10421_),
    .B2(_10766_),
    .X(_10767_));
 sky130_fd_sc_hd__a2bb2o_1 _26687_ (.A1_N(_10765_),
    .A2_N(_10767_),
    .B1(_10765_),
    .B2(_10767_),
    .X(_10768_));
 sky130_fd_sc_hd__a2bb2o_1 _26688_ (.A1_N(_10764_),
    .A2_N(_10768_),
    .B1(_10764_),
    .B2(_10768_),
    .X(_10769_));
 sky130_fd_sc_hd__o22a_1 _26689_ (.A1(_10679_),
    .A2(_10680_),
    .B1(_10681_),
    .B2(_10687_),
    .X(_10770_));
 sky130_fd_sc_hd__a2bb2o_1 _26690_ (.A1_N(_10769_),
    .A2_N(_10770_),
    .B1(_10769_),
    .B2(_10770_),
    .X(_10771_));
 sky130_fd_sc_hd__clkbuf_2 _26691_ (.A(_10275_),
    .X(_10772_));
 sky130_fd_sc_hd__o22a_1 _26692_ (.A1(_10610_),
    .A2(_10685_),
    .B1(_10611_),
    .B2(_10686_),
    .X(_10773_));
 sky130_fd_sc_hd__or2_1 _26693_ (.A(_10278_),
    .B(_10773_),
    .X(_10774_));
 sky130_fd_sc_hd__a21bo_1 _26694_ (.A1(_10772_),
    .A2(_10773_),
    .B1_N(_10774_),
    .X(_10775_));
 sky130_fd_sc_hd__a2bb2o_1 _26695_ (.A1_N(_10771_),
    .A2_N(_10775_),
    .B1(_10771_),
    .B2(_10775_),
    .X(_10776_));
 sky130_fd_sc_hd__o22a_1 _26696_ (.A1(_10688_),
    .A2(_10689_),
    .B1(_10614_),
    .B2(_10690_),
    .X(_10777_));
 sky130_fd_sc_hd__a2bb2o_1 _26697_ (.A1_N(_10776_),
    .A2_N(_10777_),
    .B1(_10776_),
    .B2(_10777_),
    .X(_10778_));
 sky130_fd_sc_hd__a2bb2o_1 _26698_ (.A1_N(_10613_),
    .A2_N(_10778_),
    .B1(_10613_),
    .B2(_10778_),
    .X(_10779_));
 sky130_fd_sc_hd__o22a_1 _26699_ (.A1(_10691_),
    .A2(_10692_),
    .B1(_10517_),
    .B2(_10693_),
    .X(_10780_));
 sky130_fd_sc_hd__or2_1 _26700_ (.A(_10779_),
    .B(_10780_),
    .X(_10781_));
 sky130_fd_sc_hd__a21bo_1 _26701_ (.A1(_10779_),
    .A2(_10780_),
    .B1_N(_10781_),
    .X(_10782_));
 sky130_fd_sc_hd__buf_1 _26702_ (.A(_10782_),
    .X(_10783_));
 sky130_fd_sc_hd__or2_1 _26703_ (.A(_10607_),
    .B(_10698_),
    .X(_10784_));
 sky130_fd_sc_hd__or3_1 _26704_ (.A(_10399_),
    .B(_10513_),
    .C(_10784_),
    .X(_10785_));
 sky130_fd_sc_hd__o221a_1 _26705_ (.A1(_10606_),
    .A2(_10696_),
    .B1(_10608_),
    .B2(_10784_),
    .C1(_10697_),
    .X(_10786_));
 sky130_fd_sc_hd__o21ai_1 _26706_ (.A1(_10406_),
    .A2(_10785_),
    .B1(_10786_),
    .Y(_10787_));
 sky130_vsdinv _26707_ (.A(_10787_),
    .Y(_10788_));
 sky130_vsdinv _26708_ (.A(_10783_),
    .Y(_10789_));
 sky130_fd_sc_hd__o22a_1 _26709_ (.A1(_10783_),
    .A2(_10788_),
    .B1(_10789_),
    .B2(_10787_),
    .X(_02671_));
 sky130_fd_sc_hd__o21ai_1 _26710_ (.A1(_10783_),
    .A2(_10788_),
    .B1(_10781_),
    .Y(_10790_));
 sky130_fd_sc_hd__buf_1 _26711_ (.A(_10140_),
    .X(_10791_));
 sky130_fd_sc_hd__and4_2 _26712_ (.A(_10791_),
    .B(_06878_),
    .C(_13066_),
    .D(_06884_),
    .X(_10792_));
 sky130_fd_sc_hd__o22a_1 _26713_ (.A1(_11719_),
    .A2(_13551_),
    .B1(_10616_),
    .B2(_09025_),
    .X(_10793_));
 sky130_fd_sc_hd__nor2_2 _26714_ (.A(_10792_),
    .B(_10793_),
    .Y(_10794_));
 sky130_fd_sc_hd__clkbuf_4 _26715_ (.A(_07972_),
    .X(_10795_));
 sky130_fd_sc_hd__nor2_4 _26716_ (.A(_10795_),
    .B(_07321_),
    .Y(_10796_));
 sky130_fd_sc_hd__a2bb2o_2 _26717_ (.A1_N(_10794_),
    .A2_N(_10796_),
    .B1(_10794_),
    .B2(_10796_),
    .X(_10797_));
 sky130_fd_sc_hd__a21oi_4 _26718_ (.A1(_10702_),
    .A2(_10703_),
    .B1(_10700_),
    .Y(_10798_));
 sky130_fd_sc_hd__o2bb2ai_2 _26719_ (.A1_N(_10797_),
    .A2_N(_10798_),
    .B1(_10797_),
    .B2(_10798_),
    .Y(_10799_));
 sky130_fd_sc_hd__buf_1 _26720_ (.A(_09918_),
    .X(_10800_));
 sky130_fd_sc_hd__o22a_1 _26721_ (.A1(_10800_),
    .A2(_07459_),
    .B1(_10623_),
    .B2(_10327_),
    .X(_10801_));
 sky130_fd_sc_hd__and4_1 _26722_ (.A(_13075_),
    .B(_13540_),
    .C(_13081_),
    .D(_13536_),
    .X(_10802_));
 sky130_fd_sc_hd__nor2_2 _26723_ (.A(_10801_),
    .B(_10802_),
    .Y(_10803_));
 sky130_fd_sc_hd__clkbuf_2 _26724_ (.A(_07532_),
    .X(_10804_));
 sky130_fd_sc_hd__clkbuf_2 _26725_ (.A(_10329_),
    .X(_10805_));
 sky130_fd_sc_hd__nor2_2 _26726_ (.A(_10804_),
    .B(_10805_),
    .Y(_10806_));
 sky130_fd_sc_hd__a2bb2o_2 _26727_ (.A1_N(_10803_),
    .A2_N(_10806_),
    .B1(_10803_),
    .B2(_10806_),
    .X(_10807_));
 sky130_fd_sc_hd__o2bb2ai_2 _26728_ (.A1_N(_10799_),
    .A2_N(_10807_),
    .B1(_10799_),
    .B2(_10807_),
    .Y(_10808_));
 sky130_fd_sc_hd__o22a_2 _26729_ (.A1(_10704_),
    .A2(_10705_),
    .B1(_10706_),
    .B2(_10712_),
    .X(_10809_));
 sky130_fd_sc_hd__o2bb2ai_2 _26730_ (.A1_N(_10808_),
    .A2_N(_10809_),
    .B1(_10808_),
    .B2(_10809_),
    .Y(_10810_));
 sky130_fd_sc_hd__a21oi_2 _26731_ (.A1(_10720_),
    .A2(_10721_),
    .B1(_10719_),
    .Y(_10811_));
 sky130_fd_sc_hd__a21oi_4 _26732_ (.A1(_10709_),
    .A2(_10711_),
    .B1(_10708_),
    .Y(_10812_));
 sky130_fd_sc_hd__o22a_1 _26733_ (.A1(_10465_),
    .A2(_10012_),
    .B1(_10368_),
    .B2(_09007_),
    .X(_10813_));
 sky130_fd_sc_hd__and4_1 _26734_ (.A(_10370_),
    .B(_07588_),
    .C(_10371_),
    .D(_07878_),
    .X(_10814_));
 sky130_fd_sc_hd__nor2_2 _26735_ (.A(_10813_),
    .B(_10814_),
    .Y(_10815_));
 sky130_fd_sc_hd__nor2_2 _26736_ (.A(_10374_),
    .B(_08175_),
    .Y(_10816_));
 sky130_fd_sc_hd__a2bb2o_1 _26737_ (.A1_N(_10815_),
    .A2_N(_10816_),
    .B1(_10815_),
    .B2(_10816_),
    .X(_10817_));
 sky130_fd_sc_hd__a2bb2o_1 _26738_ (.A1_N(_10812_),
    .A2_N(_10817_),
    .B1(_10812_),
    .B2(_10817_),
    .X(_10818_));
 sky130_fd_sc_hd__a2bb2o_2 _26739_ (.A1_N(_10811_),
    .A2_N(_10818_),
    .B1(_10811_),
    .B2(_10818_),
    .X(_10819_));
 sky130_fd_sc_hd__o2bb2ai_2 _26740_ (.A1_N(_10810_),
    .A2_N(_10819_),
    .B1(_10810_),
    .B2(_10819_),
    .Y(_10820_));
 sky130_fd_sc_hd__o22a_1 _26741_ (.A1(_10713_),
    .A2(_10714_),
    .B1(_10715_),
    .B2(_10724_),
    .X(_10821_));
 sky130_fd_sc_hd__o2bb2ai_1 _26742_ (.A1_N(_10820_),
    .A2_N(_10821_),
    .B1(_10820_),
    .B2(_10821_),
    .Y(_10822_));
 sky130_fd_sc_hd__buf_1 _26743_ (.A(_10732_),
    .X(_10823_));
 sky130_fd_sc_hd__o22a_1 _26744_ (.A1(_10738_),
    .A2(_10739_),
    .B1(_10823_),
    .B2(_10740_),
    .X(_10824_));
 sky130_fd_sc_hd__o22a_1 _26745_ (.A1(_10717_),
    .A2(_10722_),
    .B1(_10716_),
    .B2(_10723_),
    .X(_10825_));
 sky130_fd_sc_hd__o22a_1 _26746_ (.A1(_10563_),
    .A2(_08839_),
    .B1(_10564_),
    .B2(_08498_),
    .X(_10826_));
 sky130_fd_sc_hd__and4_1 _26747_ (.A(_10653_),
    .B(_08172_),
    .C(_10654_),
    .D(_08820_),
    .X(_10827_));
 sky130_fd_sc_hd__nor2_2 _26748_ (.A(_10826_),
    .B(_10827_),
    .Y(_10828_));
 sky130_fd_sc_hd__or2_2 _26749_ (.A(_11703_),
    .B(_06803_),
    .X(_10829_));
 sky130_vsdinv _26750_ (.A(_10829_),
    .Y(_10830_));
 sky130_fd_sc_hd__buf_1 _26751_ (.A(_10830_),
    .X(_10831_));
 sky130_fd_sc_hd__a2bb2o_1 _26752_ (.A1_N(_10828_),
    .A2_N(_10831_),
    .B1(_10828_),
    .B2(_10831_),
    .X(_10832_));
 sky130_fd_sc_hd__a31o_1 _26753_ (.A1(\pcpi_mul.rs2[21] ),
    .A2(_13507_),
    .A3(_10736_),
    .B1(_10735_),
    .X(_10833_));
 sky130_vsdinv _26754_ (.A(_10833_),
    .Y(_10834_));
 sky130_vsdinv _26755_ (.A(_10832_),
    .Y(_10835_));
 sky130_fd_sc_hd__a22o_1 _26756_ (.A1(_10832_),
    .A2(_10834_),
    .B1(_10835_),
    .B2(_10833_),
    .X(_10836_));
 sky130_fd_sc_hd__a2bb2o_1 _26757_ (.A1_N(_10733_),
    .A2_N(_10836_),
    .B1(_10732_),
    .B2(_10836_),
    .X(_10837_));
 sky130_fd_sc_hd__a2bb2o_1 _26758_ (.A1_N(_10825_),
    .A2_N(_10837_),
    .B1(_10825_),
    .B2(_10837_),
    .X(_10838_));
 sky130_fd_sc_hd__a2bb2o_1 _26759_ (.A1_N(_10824_),
    .A2_N(_10838_),
    .B1(_10824_),
    .B2(_10838_),
    .X(_10839_));
 sky130_fd_sc_hd__o2bb2ai_1 _26760_ (.A1_N(_10822_),
    .A2_N(_10839_),
    .B1(_10822_),
    .B2(_10839_),
    .Y(_10840_));
 sky130_fd_sc_hd__o22a_1 _26761_ (.A1(_10725_),
    .A2(_10726_),
    .B1(_10727_),
    .B2(_10743_),
    .X(_10841_));
 sky130_fd_sc_hd__o2bb2a_1 _26762_ (.A1_N(_10840_),
    .A2_N(_10841_),
    .B1(_10840_),
    .B2(_10841_),
    .X(_10842_));
 sky130_vsdinv _26763_ (.A(_10842_),
    .Y(_10843_));
 sky130_fd_sc_hd__o22a_1 _26764_ (.A1(_10750_),
    .A2(_10756_),
    .B1(_10291_),
    .B2(_10757_),
    .X(_10844_));
 sky130_fd_sc_hd__o22a_1 _26765_ (.A1(_10729_),
    .A2(_10741_),
    .B1(_10728_),
    .B2(_10742_),
    .X(_10845_));
 sky130_fd_sc_hd__o22a_2 _26766_ (.A1(_10648_),
    .A2(_10730_),
    .B1(_10559_),
    .B2(_10731_),
    .X(_10846_));
 sky130_fd_sc_hd__o22ai_1 _26767_ (.A1(_06001_),
    .A2(_10430_),
    .B1(_10753_),
    .B2(_10754_),
    .Y(_10847_));
 sky130_fd_sc_hd__o2bb2a_1 _26768_ (.A1_N(_10846_),
    .A2_N(_10847_),
    .B1(_10846_),
    .B2(_10847_),
    .X(_10848_));
 sky130_fd_sc_hd__a2bb2o_1 _26769_ (.A1_N(_10290_),
    .A2_N(_10848_),
    .B1(_10290_),
    .B2(_10848_),
    .X(_10849_));
 sky130_fd_sc_hd__a2bb2o_1 _26770_ (.A1_N(_10845_),
    .A2_N(_10849_),
    .B1(_10845_),
    .B2(_10849_),
    .X(_10850_));
 sky130_fd_sc_hd__a2bb2o_1 _26771_ (.A1_N(_10844_),
    .A2_N(_10850_),
    .B1(_10844_),
    .B2(_10850_),
    .X(_10851_));
 sky130_vsdinv _26772_ (.A(_10851_),
    .Y(_10852_));
 sky130_fd_sc_hd__a22o_1 _26773_ (.A1(_10843_),
    .A2(_10851_),
    .B1(_10842_),
    .B2(_10852_),
    .X(_10853_));
 sky130_fd_sc_hd__o22a_1 _26774_ (.A1(_10744_),
    .A2(_10745_),
    .B1(_10747_),
    .B2(_10760_),
    .X(_10854_));
 sky130_fd_sc_hd__a2bb2o_1 _26775_ (.A1_N(_10853_),
    .A2_N(_10854_),
    .B1(_10853_),
    .B2(_10854_),
    .X(_10855_));
 sky130_fd_sc_hd__o22a_1 _26776_ (.A1(_10749_),
    .A2(_10758_),
    .B1(_10748_),
    .B2(_10759_),
    .X(_10856_));
 sky130_fd_sc_hd__a2bb2o_1 _26777_ (.A1_N(_10514_),
    .A2_N(_10856_),
    .B1(_10514_),
    .B2(_10856_),
    .X(_10857_));
 sky130_fd_sc_hd__a2bb2o_1 _26778_ (.A1_N(_10765_),
    .A2_N(_10857_),
    .B1(_10520_),
    .B2(_10857_),
    .X(_10858_));
 sky130_fd_sc_hd__a2bb2o_1 _26779_ (.A1_N(_10855_),
    .A2_N(_10858_),
    .B1(_10855_),
    .B2(_10858_),
    .X(_10859_));
 sky130_fd_sc_hd__o22a_1 _26780_ (.A1(_10762_),
    .A2(_10763_),
    .B1(_10764_),
    .B2(_10768_),
    .X(_10860_));
 sky130_fd_sc_hd__a2bb2o_1 _26781_ (.A1_N(_10859_),
    .A2_N(_10860_),
    .B1(_10859_),
    .B2(_10860_),
    .X(_10861_));
 sky130_fd_sc_hd__o22a_1 _26782_ (.A1(_10515_),
    .A2(_10766_),
    .B1(_10682_),
    .B2(_10767_),
    .X(_10862_));
 sky130_fd_sc_hd__or2_1 _26783_ (.A(_10410_),
    .B(_10862_),
    .X(_10863_));
 sky130_fd_sc_hd__a21bo_1 _26784_ (.A1(_10276_),
    .A2(_10862_),
    .B1_N(_10863_),
    .X(_10864_));
 sky130_fd_sc_hd__a2bb2o_1 _26785_ (.A1_N(_10861_),
    .A2_N(_10864_),
    .B1(_10861_),
    .B2(_10864_),
    .X(_10865_));
 sky130_fd_sc_hd__o22a_1 _26786_ (.A1(_10769_),
    .A2(_10770_),
    .B1(_10771_),
    .B2(_10775_),
    .X(_10866_));
 sky130_fd_sc_hd__a2bb2o_1 _26787_ (.A1_N(_10865_),
    .A2_N(_10866_),
    .B1(_10865_),
    .B2(_10866_),
    .X(_10867_));
 sky130_fd_sc_hd__a2bb2o_1 _26788_ (.A1_N(_10774_),
    .A2_N(_10867_),
    .B1(_10774_),
    .B2(_10867_),
    .X(_10868_));
 sky130_fd_sc_hd__o22a_1 _26789_ (.A1(_10776_),
    .A2(_10777_),
    .B1(_10613_),
    .B2(_10778_),
    .X(_10869_));
 sky130_fd_sc_hd__or2_1 _26790_ (.A(_10868_),
    .B(_10869_),
    .X(_10870_));
 sky130_fd_sc_hd__a21bo_1 _26791_ (.A1(_10868_),
    .A2(_10869_),
    .B1_N(_10870_),
    .X(_10871_));
 sky130_fd_sc_hd__a2bb2o_1 _26792_ (.A1_N(_10790_),
    .A2_N(_10871_),
    .B1(_10790_),
    .B2(_10871_),
    .X(_02672_));
 sky130_fd_sc_hd__and4_2 _26793_ (.A(_10791_),
    .B(_06763_),
    .C(_13067_),
    .D(_13542_),
    .X(_10872_));
 sky130_fd_sc_hd__buf_1 _26794_ (.A(_10616_),
    .X(_10873_));
 sky130_fd_sc_hd__o22a_1 _26795_ (.A1(_11719_),
    .A2(_13547_),
    .B1(_10873_),
    .B2(_07020_),
    .X(_10874_));
 sky130_fd_sc_hd__nor2_2 _26796_ (.A(_10872_),
    .B(_10874_),
    .Y(_10875_));
 sky130_fd_sc_hd__nor2_4 _26797_ (.A(_10795_),
    .B(_10375_),
    .Y(_10876_));
 sky130_fd_sc_hd__a2bb2o_2 _26798_ (.A1_N(_10875_),
    .A2_N(_10876_),
    .B1(_10875_),
    .B2(_10876_),
    .X(_10877_));
 sky130_fd_sc_hd__a21oi_4 _26799_ (.A1(_10794_),
    .A2(_10796_),
    .B1(_10792_),
    .Y(_10878_));
 sky130_fd_sc_hd__o2bb2ai_4 _26800_ (.A1_N(_10877_),
    .A2_N(_10878_),
    .B1(_10877_),
    .B2(_10878_),
    .Y(_10879_));
 sky130_fd_sc_hd__buf_1 _26801_ (.A(_10623_),
    .X(_10880_));
 sky130_fd_sc_hd__o22a_1 _26802_ (.A1(_10800_),
    .A2(_10327_),
    .B1(_10880_),
    .B2(_10329_),
    .X(_10881_));
 sky130_fd_sc_hd__and4_2 _26803_ (.A(_13075_),
    .B(_13537_),
    .C(_13082_),
    .D(_13530_),
    .X(_10882_));
 sky130_fd_sc_hd__nor2_2 _26804_ (.A(_10881_),
    .B(_10882_),
    .Y(_10883_));
 sky130_fd_sc_hd__nor2_2 _26805_ (.A(_10804_),
    .B(_10334_),
    .Y(_10884_));
 sky130_fd_sc_hd__a2bb2o_2 _26806_ (.A1_N(_10883_),
    .A2_N(_10884_),
    .B1(_10883_),
    .B2(_10884_),
    .X(_10885_));
 sky130_fd_sc_hd__o2bb2ai_4 _26807_ (.A1_N(_10879_),
    .A2_N(_10885_),
    .B1(_10879_),
    .B2(_10885_),
    .Y(_10886_));
 sky130_fd_sc_hd__o22a_2 _26808_ (.A1(_10797_),
    .A2(_10798_),
    .B1(_10799_),
    .B2(_10807_),
    .X(_10887_));
 sky130_fd_sc_hd__o2bb2ai_2 _26809_ (.A1_N(_10886_),
    .A2_N(_10887_),
    .B1(_10886_),
    .B2(_10887_),
    .Y(_10888_));
 sky130_fd_sc_hd__a21oi_2 _26810_ (.A1(_10815_),
    .A2(_10816_),
    .B1(_10814_),
    .Y(_10889_));
 sky130_fd_sc_hd__a21oi_2 _26811_ (.A1(_10803_),
    .A2(_10806_),
    .B1(_10802_),
    .Y(_10890_));
 sky130_fd_sc_hd__o22a_1 _26812_ (.A1(_10367_),
    .A2(_09007_),
    .B1(_10368_),
    .B2(_10480_),
    .X(_10891_));
 sky130_fd_sc_hd__and4_1 _26813_ (.A(_10370_),
    .B(_13521_),
    .C(_13094_),
    .D(_08024_),
    .X(_10892_));
 sky130_fd_sc_hd__nor2_2 _26814_ (.A(_10891_),
    .B(_10892_),
    .Y(_10893_));
 sky130_fd_sc_hd__nor2_2 _26815_ (.A(_10374_),
    .B(_10323_),
    .Y(_10894_));
 sky130_fd_sc_hd__a2bb2o_1 _26816_ (.A1_N(_10893_),
    .A2_N(_10894_),
    .B1(_10893_),
    .B2(_10894_),
    .X(_10895_));
 sky130_fd_sc_hd__a2bb2o_1 _26817_ (.A1_N(_10890_),
    .A2_N(_10895_),
    .B1(_10890_),
    .B2(_10895_),
    .X(_10896_));
 sky130_fd_sc_hd__a2bb2o_2 _26818_ (.A1_N(_10889_),
    .A2_N(_10896_),
    .B1(_10889_),
    .B2(_10896_),
    .X(_10897_));
 sky130_fd_sc_hd__o2bb2ai_2 _26819_ (.A1_N(_10888_),
    .A2_N(_10897_),
    .B1(_10888_),
    .B2(_10897_),
    .Y(_10898_));
 sky130_fd_sc_hd__o22a_1 _26820_ (.A1(_10808_),
    .A2(_10809_),
    .B1(_10810_),
    .B2(_10819_),
    .X(_10899_));
 sky130_fd_sc_hd__o2bb2ai_1 _26821_ (.A1_N(_10898_),
    .A2_N(_10899_),
    .B1(_10898_),
    .B2(_10899_),
    .Y(_10900_));
 sky130_fd_sc_hd__o22a_1 _26822_ (.A1(_10832_),
    .A2(_10834_),
    .B1(_10823_),
    .B2(_10836_),
    .X(_10901_));
 sky130_fd_sc_hd__o22a_1 _26823_ (.A1(_10812_),
    .A2(_10817_),
    .B1(_10811_),
    .B2(_10818_),
    .X(_10902_));
 sky130_fd_sc_hd__buf_1 _26824_ (.A(_10732_),
    .X(_10903_));
 sky130_fd_sc_hd__a31o_1 _26825_ (.A1(_10088_),
    .A2(\pcpi_mul.rs2[21] ),
    .A3(_10828_),
    .B1(_10827_),
    .X(_10904_));
 sky130_vsdinv _26826_ (.A(_10904_),
    .Y(_10905_));
 sky130_fd_sc_hd__o22a_1 _26827_ (.A1(_10563_),
    .A2(_09239_),
    .B1(_08661_),
    .B2(_10564_),
    .X(_10906_));
 sky130_fd_sc_hd__and4_1 _26828_ (.A(_10653_),
    .B(_13506_),
    .C(_08815_),
    .D(_10654_),
    .X(_10907_));
 sky130_fd_sc_hd__nor2_1 _26829_ (.A(_10906_),
    .B(_10907_),
    .Y(_10908_));
 sky130_fd_sc_hd__o2bb2a_1 _26830_ (.A1_N(_10831_),
    .A2_N(_10908_),
    .B1(_10830_),
    .B2(_10908_),
    .X(_10909_));
 sky130_vsdinv _26831_ (.A(_10909_),
    .Y(_10910_));
 sky130_fd_sc_hd__a22o_1 _26832_ (.A1(_10905_),
    .A2(_10910_),
    .B1(_10904_),
    .B2(_10909_),
    .X(_10911_));
 sky130_fd_sc_hd__a2bb2o_1 _26833_ (.A1_N(_10903_),
    .A2_N(_10911_),
    .B1(_10733_),
    .B2(_10911_),
    .X(_10912_));
 sky130_fd_sc_hd__a2bb2o_1 _26834_ (.A1_N(_10902_),
    .A2_N(_10912_),
    .B1(_10902_),
    .B2(_10912_),
    .X(_10913_));
 sky130_fd_sc_hd__a2bb2o_1 _26835_ (.A1_N(_10901_),
    .A2_N(_10913_),
    .B1(_10901_),
    .B2(_10913_),
    .X(_10914_));
 sky130_fd_sc_hd__o2bb2ai_1 _26836_ (.A1_N(_10900_),
    .A2_N(_10914_),
    .B1(_10900_),
    .B2(_10914_),
    .Y(_10915_));
 sky130_fd_sc_hd__o22a_1 _26837_ (.A1(_10820_),
    .A2(_10821_),
    .B1(_10822_),
    .B2(_10839_),
    .X(_10916_));
 sky130_fd_sc_hd__o2bb2a_1 _26838_ (.A1_N(_10915_),
    .A2_N(_10916_),
    .B1(_10915_),
    .B2(_10916_),
    .X(_10917_));
 sky130_vsdinv _26839_ (.A(_10917_),
    .Y(_10918_));
 sky130_fd_sc_hd__or3_4 _26840_ (.A(_06001_),
    .B(_10430_),
    .C(_10846_),
    .X(_10919_));
 sky130_fd_sc_hd__o21a_1 _26841_ (.A1(_10291_),
    .A2(_10848_),
    .B1(_10919_),
    .X(_10920_));
 sky130_fd_sc_hd__o22a_1 _26842_ (.A1(_10825_),
    .A2(_10837_),
    .B1(_10824_),
    .B2(_10838_),
    .X(_10921_));
 sky130_vsdinv _26843_ (.A(_10919_),
    .Y(_10922_));
 sky130_fd_sc_hd__and3_1 _26844_ (.A(_10582_),
    .B(_10846_),
    .C(_10585_),
    .X(_10923_));
 sky130_fd_sc_hd__or2_1 _26845_ (.A(_10922_),
    .B(_10923_),
    .X(_10924_));
 sky130_fd_sc_hd__a2bb2o_1 _26846_ (.A1_N(_10294_),
    .A2_N(_10924_),
    .B1(_10294_),
    .B2(_10924_),
    .X(_10925_));
 sky130_fd_sc_hd__buf_1 _26847_ (.A(_10925_),
    .X(_10926_));
 sky130_fd_sc_hd__a2bb2o_1 _26848_ (.A1_N(_10921_),
    .A2_N(_10926_),
    .B1(_10921_),
    .B2(_10925_),
    .X(_10927_));
 sky130_fd_sc_hd__a2bb2o_1 _26849_ (.A1_N(_10920_),
    .A2_N(_10927_),
    .B1(_10920_),
    .B2(_10927_),
    .X(_10928_));
 sky130_vsdinv _26850_ (.A(_10928_),
    .Y(_10929_));
 sky130_fd_sc_hd__a22o_1 _26851_ (.A1(_10918_),
    .A2(_10928_),
    .B1(_10917_),
    .B2(_10929_),
    .X(_10930_));
 sky130_fd_sc_hd__o22a_1 _26852_ (.A1(_10840_),
    .A2(_10841_),
    .B1(_10843_),
    .B2(_10851_),
    .X(_10931_));
 sky130_fd_sc_hd__a2bb2o_1 _26853_ (.A1_N(_10930_),
    .A2_N(_10931_),
    .B1(_10930_),
    .B2(_10931_),
    .X(_10932_));
 sky130_fd_sc_hd__o22a_1 _26854_ (.A1(_10845_),
    .A2(_10849_),
    .B1(_10844_),
    .B2(_10850_),
    .X(_10933_));
 sky130_fd_sc_hd__a2bb2o_1 _26855_ (.A1_N(_10684_),
    .A2_N(_10933_),
    .B1(_10521_),
    .B2(_10933_),
    .X(_10934_));
 sky130_fd_sc_hd__a2bb2o_1 _26856_ (.A1_N(_10520_),
    .A2_N(_10934_),
    .B1(_10611_),
    .B2(_10934_),
    .X(_10935_));
 sky130_fd_sc_hd__a2bb2o_1 _26857_ (.A1_N(_10932_),
    .A2_N(_10935_),
    .B1(_10932_),
    .B2(_10935_),
    .X(_10936_));
 sky130_fd_sc_hd__o22a_1 _26858_ (.A1(_10853_),
    .A2(_10854_),
    .B1(_10855_),
    .B2(_10858_),
    .X(_10937_));
 sky130_fd_sc_hd__a2bb2o_1 _26859_ (.A1_N(_10936_),
    .A2_N(_10937_),
    .B1(_10936_),
    .B2(_10937_),
    .X(_10938_));
 sky130_fd_sc_hd__o22a_1 _26860_ (.A1(_10515_),
    .A2(_10856_),
    .B1(_10682_),
    .B2(_10857_),
    .X(_10939_));
 sky130_fd_sc_hd__or2_1 _26861_ (.A(_10410_),
    .B(_10939_),
    .X(_10940_));
 sky130_fd_sc_hd__a21bo_1 _26862_ (.A1(_10276_),
    .A2(_10939_),
    .B1_N(_10940_),
    .X(_10941_));
 sky130_fd_sc_hd__a2bb2o_1 _26863_ (.A1_N(_10938_),
    .A2_N(_10941_),
    .B1(_10938_),
    .B2(_10941_),
    .X(_10942_));
 sky130_fd_sc_hd__o22a_1 _26864_ (.A1(_10859_),
    .A2(_10860_),
    .B1(_10861_),
    .B2(_10864_),
    .X(_10943_));
 sky130_fd_sc_hd__a2bb2o_1 _26865_ (.A1_N(_10942_),
    .A2_N(_10943_),
    .B1(_10942_),
    .B2(_10943_),
    .X(_10944_));
 sky130_fd_sc_hd__a2bb2o_1 _26866_ (.A1_N(_10863_),
    .A2_N(_10944_),
    .B1(_10863_),
    .B2(_10944_),
    .X(_10945_));
 sky130_fd_sc_hd__o22a_1 _26867_ (.A1(_10865_),
    .A2(_10866_),
    .B1(_10774_),
    .B2(_10867_),
    .X(_10946_));
 sky130_fd_sc_hd__or2_1 _26868_ (.A(_10945_),
    .B(_10946_),
    .X(_10947_));
 sky130_fd_sc_hd__a21bo_1 _26869_ (.A1(_10945_),
    .A2(_10946_),
    .B1_N(_10947_),
    .X(_10948_));
 sky130_fd_sc_hd__a22o_1 _26870_ (.A1(_10868_),
    .A2(_10869_),
    .B1(_10781_),
    .B2(_10870_),
    .X(_10949_));
 sky130_fd_sc_hd__o31a_1 _26871_ (.A1(_10783_),
    .A2(_10871_),
    .A3(_10788_),
    .B1(_10949_),
    .X(_10950_));
 sky130_fd_sc_hd__a2bb2oi_1 _26872_ (.A1_N(_10948_),
    .A2_N(_10950_),
    .B1(_10948_),
    .B2(_10950_),
    .Y(_02673_));
 sky130_fd_sc_hd__and4_2 _26873_ (.A(_10791_),
    .B(_07171_),
    .C(_13067_),
    .D(_07175_),
    .X(_10951_));
 sky130_fd_sc_hd__o22a_1 _26874_ (.A1(_11720_),
    .A2(_13543_),
    .B1(_10873_),
    .B2(_07459_),
    .X(_10952_));
 sky130_fd_sc_hd__nor2_2 _26875_ (.A(_10951_),
    .B(_10952_),
    .Y(_10953_));
 sky130_fd_sc_hd__nor2_4 _26876_ (.A(_10795_),
    .B(_10710_),
    .Y(_10954_));
 sky130_fd_sc_hd__a2bb2o_2 _26877_ (.A1_N(_10953_),
    .A2_N(_10954_),
    .B1(_10953_),
    .B2(_10954_),
    .X(_10955_));
 sky130_fd_sc_hd__a21oi_4 _26878_ (.A1(_10875_),
    .A2(_10876_),
    .B1(_10872_),
    .Y(_10956_));
 sky130_fd_sc_hd__o2bb2ai_2 _26879_ (.A1_N(_10955_),
    .A2_N(_10956_),
    .B1(_10955_),
    .B2(_10956_),
    .Y(_10957_));
 sky130_fd_sc_hd__o22a_1 _26880_ (.A1(_10800_),
    .A2(_10329_),
    .B1(_10880_),
    .B2(_10334_),
    .X(_10958_));
 sky130_fd_sc_hd__and4_1 _26881_ (.A(_13076_),
    .B(_13531_),
    .C(_13082_),
    .D(_13525_),
    .X(_10959_));
 sky130_fd_sc_hd__nor2_2 _26882_ (.A(_10958_),
    .B(_10959_),
    .Y(_10960_));
 sky130_fd_sc_hd__nor2_2 _26883_ (.A(_10804_),
    .B(_10489_),
    .Y(_10961_));
 sky130_fd_sc_hd__a2bb2o_2 _26884_ (.A1_N(_10960_),
    .A2_N(_10961_),
    .B1(_10960_),
    .B2(_10961_),
    .X(_10962_));
 sky130_fd_sc_hd__o2bb2ai_2 _26885_ (.A1_N(_10957_),
    .A2_N(_10962_),
    .B1(_10957_),
    .B2(_10962_),
    .Y(_10963_));
 sky130_fd_sc_hd__o22a_2 _26886_ (.A1(_10877_),
    .A2(_10878_),
    .B1(_10879_),
    .B2(_10885_),
    .X(_10964_));
 sky130_fd_sc_hd__o2bb2ai_2 _26887_ (.A1_N(_10963_),
    .A2_N(_10964_),
    .B1(_10963_),
    .B2(_10964_),
    .Y(_10965_));
 sky130_fd_sc_hd__a21oi_2 _26888_ (.A1(_10893_),
    .A2(_10894_),
    .B1(_10892_),
    .Y(_10966_));
 sky130_fd_sc_hd__a21oi_2 _26889_ (.A1(_10883_),
    .A2(_10884_),
    .B1(_10882_),
    .Y(_10967_));
 sky130_fd_sc_hd__o22a_1 _26890_ (.A1(_10367_),
    .A2(_08175_),
    .B1(_07270_),
    .B2(_07892_),
    .X(_10968_));
 sky130_fd_sc_hd__and4_2 _26891_ (.A(_13090_),
    .B(_13517_),
    .C(_13094_),
    .D(_13511_),
    .X(_10969_));
 sky130_fd_sc_hd__nor2_2 _26892_ (.A(_10968_),
    .B(_10969_),
    .Y(_10970_));
 sky130_fd_sc_hd__nor2_2 _26893_ (.A(_07076_),
    .B(_08500_),
    .Y(_10971_));
 sky130_fd_sc_hd__a2bb2o_1 _26894_ (.A1_N(_10970_),
    .A2_N(_10971_),
    .B1(_10970_),
    .B2(_10971_),
    .X(_10972_));
 sky130_fd_sc_hd__a2bb2o_1 _26895_ (.A1_N(_10967_),
    .A2_N(_10972_),
    .B1(_10967_),
    .B2(_10972_),
    .X(_10973_));
 sky130_fd_sc_hd__a2bb2o_2 _26896_ (.A1_N(_10966_),
    .A2_N(_10973_),
    .B1(_10966_),
    .B2(_10973_),
    .X(_10974_));
 sky130_fd_sc_hd__o2bb2ai_2 _26897_ (.A1_N(_10965_),
    .A2_N(_10974_),
    .B1(_10965_),
    .B2(_10974_),
    .Y(_10975_));
 sky130_fd_sc_hd__o22a_1 _26898_ (.A1(_10886_),
    .A2(_10887_),
    .B1(_10888_),
    .B2(_10897_),
    .X(_10976_));
 sky130_fd_sc_hd__o2bb2ai_1 _26899_ (.A1_N(_10975_),
    .A2_N(_10976_),
    .B1(_10975_),
    .B2(_10976_),
    .Y(_10977_));
 sky130_fd_sc_hd__o22a_1 _26900_ (.A1(_10905_),
    .A2(_10910_),
    .B1(_10823_),
    .B2(_10911_),
    .X(_10978_));
 sky130_fd_sc_hd__o22a_1 _26901_ (.A1(_10890_),
    .A2(_10895_),
    .B1(_10889_),
    .B2(_10896_),
    .X(_10979_));
 sky130_fd_sc_hd__buf_1 _26902_ (.A(_11704_),
    .X(_10980_));
 sky130_fd_sc_hd__o22a_1 _26903_ (.A1(_10980_),
    .A2(_10328_),
    .B1(_10980_),
    .B2(_10326_),
    .X(_10981_));
 sky130_fd_sc_hd__or4_4 _26904_ (.A(_11705_),
    .B(_10328_),
    .C(_11705_),
    .D(_10326_),
    .X(_10982_));
 sky130_fd_sc_hd__or2b_2 _26905_ (.A(_10981_),
    .B_N(_10982_),
    .X(_10983_));
 sky130_fd_sc_hd__o22a_1 _26906_ (.A1(_10831_),
    .A2(_10907_),
    .B1(_10333_),
    .B2(_10906_),
    .X(_10984_));
 sky130_fd_sc_hd__a2bb2oi_2 _26907_ (.A1_N(_10983_),
    .A2_N(_10984_),
    .B1(_10983_),
    .B2(_10984_),
    .Y(_10985_));
 sky130_fd_sc_hd__a2bb2o_1 _26908_ (.A1_N(_10903_),
    .A2_N(_10985_),
    .B1(_10903_),
    .B2(_10985_),
    .X(_10986_));
 sky130_fd_sc_hd__a2bb2o_1 _26909_ (.A1_N(_10979_),
    .A2_N(_10986_),
    .B1(_10979_),
    .B2(_10986_),
    .X(_10987_));
 sky130_fd_sc_hd__a2bb2o_1 _26910_ (.A1_N(_10978_),
    .A2_N(_10987_),
    .B1(_10978_),
    .B2(_10987_),
    .X(_10988_));
 sky130_fd_sc_hd__o2bb2ai_1 _26911_ (.A1_N(_10977_),
    .A2_N(_10988_),
    .B1(_10977_),
    .B2(_10988_),
    .Y(_10989_));
 sky130_fd_sc_hd__o22a_1 _26912_ (.A1(_10898_),
    .A2(_10899_),
    .B1(_10900_),
    .B2(_10914_),
    .X(_10990_));
 sky130_fd_sc_hd__o2bb2a_1 _26913_ (.A1_N(_10989_),
    .A2_N(_10990_),
    .B1(_10989_),
    .B2(_10990_),
    .X(_10991_));
 sky130_vsdinv _26914_ (.A(_10991_),
    .Y(_10992_));
 sky130_fd_sc_hd__o21a_1 _26915_ (.A1(_10314_),
    .A2(_10924_),
    .B1(_10919_),
    .X(_10993_));
 sky130_fd_sc_hd__buf_1 _26916_ (.A(_10993_),
    .X(_10994_));
 sky130_fd_sc_hd__o22a_1 _26917_ (.A1(_10902_),
    .A2(_10912_),
    .B1(_10901_),
    .B2(_10913_),
    .X(_10995_));
 sky130_fd_sc_hd__a2bb2o_1 _26918_ (.A1_N(_10926_),
    .A2_N(_10995_),
    .B1(_10926_),
    .B2(_10995_),
    .X(_10996_));
 sky130_fd_sc_hd__a2bb2o_1 _26919_ (.A1_N(_10994_),
    .A2_N(_10996_),
    .B1(_10993_),
    .B2(_10996_),
    .X(_10997_));
 sky130_vsdinv _26920_ (.A(_10997_),
    .Y(_10998_));
 sky130_fd_sc_hd__a22o_1 _26921_ (.A1(_10992_),
    .A2(_10997_),
    .B1(_10991_),
    .B2(_10998_),
    .X(_10999_));
 sky130_fd_sc_hd__o22a_1 _26922_ (.A1(_10915_),
    .A2(_10916_),
    .B1(_10918_),
    .B2(_10928_),
    .X(_11000_));
 sky130_fd_sc_hd__a2bb2o_1 _26923_ (.A1_N(_10999_),
    .A2_N(_11000_),
    .B1(_10999_),
    .B2(_11000_),
    .X(_11001_));
 sky130_fd_sc_hd__buf_1 _26924_ (.A(_10926_),
    .X(_11002_));
 sky130_fd_sc_hd__o22a_1 _26925_ (.A1(_10921_),
    .A2(_11002_),
    .B1(_10920_),
    .B2(_10927_),
    .X(_11003_));
 sky130_fd_sc_hd__a2bb2o_1 _26926_ (.A1_N(_10515_),
    .A2_N(_11003_),
    .B1(_10684_),
    .B2(_11003_),
    .X(_11004_));
 sky130_fd_sc_hd__a2bb2o_1 _26927_ (.A1_N(_10683_),
    .A2_N(_11004_),
    .B1(_10765_),
    .B2(_11004_),
    .X(_11005_));
 sky130_fd_sc_hd__a2bb2o_1 _26928_ (.A1_N(_11001_),
    .A2_N(_11005_),
    .B1(_11001_),
    .B2(_11005_),
    .X(_11006_));
 sky130_fd_sc_hd__o22a_1 _26929_ (.A1(_10930_),
    .A2(_10931_),
    .B1(_10932_),
    .B2(_10935_),
    .X(_11007_));
 sky130_fd_sc_hd__a2bb2o_1 _26930_ (.A1_N(_11006_),
    .A2_N(_11007_),
    .B1(_11006_),
    .B2(_11007_),
    .X(_11008_));
 sky130_fd_sc_hd__o22a_1 _26931_ (.A1(_10610_),
    .A2(_10933_),
    .B1(_10611_),
    .B2(_10934_),
    .X(_11009_));
 sky130_fd_sc_hd__or2_1 _26932_ (.A(_10278_),
    .B(_11009_),
    .X(_11010_));
 sky130_fd_sc_hd__a21bo_1 _26933_ (.A1(_10772_),
    .A2(_11009_),
    .B1_N(_11010_),
    .X(_11011_));
 sky130_fd_sc_hd__a2bb2o_1 _26934_ (.A1_N(_11008_),
    .A2_N(_11011_),
    .B1(_11008_),
    .B2(_11011_),
    .X(_11012_));
 sky130_fd_sc_hd__o22a_1 _26935_ (.A1(_10936_),
    .A2(_10937_),
    .B1(_10938_),
    .B2(_10941_),
    .X(_11013_));
 sky130_fd_sc_hd__a2bb2o_1 _26936_ (.A1_N(_11012_),
    .A2_N(_11013_),
    .B1(_11012_),
    .B2(_11013_),
    .X(_11014_));
 sky130_fd_sc_hd__a2bb2o_1 _26937_ (.A1_N(_10940_),
    .A2_N(_11014_),
    .B1(_10940_),
    .B2(_11014_),
    .X(_11015_));
 sky130_fd_sc_hd__o22a_1 _26938_ (.A1(_10942_),
    .A2(_10943_),
    .B1(_10863_),
    .B2(_10944_),
    .X(_11016_));
 sky130_fd_sc_hd__and2_1 _26939_ (.A(_11015_),
    .B(_11016_),
    .X(_11017_));
 sky130_fd_sc_hd__or2_1 _26940_ (.A(_11015_),
    .B(_11016_),
    .X(_11018_));
 sky130_fd_sc_hd__or2b_1 _26941_ (.A(_11017_),
    .B_N(_11018_),
    .X(_11019_));
 sky130_fd_sc_hd__o21ai_1 _26942_ (.A1(_10948_),
    .A2(_10950_),
    .B1(_10947_),
    .Y(_11020_));
 sky130_fd_sc_hd__a2bb2o_1 _26943_ (.A1_N(_11019_),
    .A2_N(_11020_),
    .B1(_11019_),
    .B2(_11020_),
    .X(_02674_));
 sky130_fd_sc_hd__buf_1 _26944_ (.A(_10791_),
    .X(_11021_));
 sky130_fd_sc_hd__buf_1 _26945_ (.A(_13067_),
    .X(_11022_));
 sky130_fd_sc_hd__and4_1 _26946_ (.A(_11021_),
    .B(_10375_),
    .C(_11022_),
    .D(_13537_),
    .X(_11023_));
 sky130_fd_sc_hd__buf_1 _26947_ (.A(_10873_),
    .X(_11024_));
 sky130_fd_sc_hd__o22a_1 _26948_ (.A1(_11720_),
    .A2(_13540_),
    .B1(_11024_),
    .B2(_10710_),
    .X(_11025_));
 sky130_fd_sc_hd__nor2_2 _26949_ (.A(_11023_),
    .B(_11025_),
    .Y(_11026_));
 sky130_fd_sc_hd__clkbuf_4 _26950_ (.A(_10795_),
    .X(_11027_));
 sky130_fd_sc_hd__nor2_4 _26951_ (.A(_11027_),
    .B(_10805_),
    .Y(_11028_));
 sky130_fd_sc_hd__a2bb2o_2 _26952_ (.A1_N(_11026_),
    .A2_N(_11028_),
    .B1(_11026_),
    .B2(_11028_),
    .X(_11029_));
 sky130_fd_sc_hd__a21oi_4 _26953_ (.A1(_10953_),
    .A2(_10954_),
    .B1(_10951_),
    .Y(_11030_));
 sky130_fd_sc_hd__o2bb2ai_4 _26954_ (.A1_N(_11029_),
    .A2_N(_11030_),
    .B1(_11029_),
    .B2(_11030_),
    .Y(_11031_));
 sky130_fd_sc_hd__buf_1 _26955_ (.A(_10800_),
    .X(_11032_));
 sky130_fd_sc_hd__clkbuf_2 _26956_ (.A(_10334_),
    .X(_11033_));
 sky130_fd_sc_hd__buf_1 _26957_ (.A(_10880_),
    .X(_11034_));
 sky130_fd_sc_hd__clkbuf_2 _26958_ (.A(_10489_),
    .X(_11035_));
 sky130_fd_sc_hd__o22a_1 _26959_ (.A1(_11032_),
    .A2(_11033_),
    .B1(_11034_),
    .B2(_11035_),
    .X(_11036_));
 sky130_fd_sc_hd__and4_2 _26960_ (.A(_13076_),
    .B(_13526_),
    .C(_13083_),
    .D(_13522_),
    .X(_11037_));
 sky130_fd_sc_hd__nor2_2 _26961_ (.A(_11036_),
    .B(_11037_),
    .Y(_11038_));
 sky130_fd_sc_hd__buf_2 _26962_ (.A(_10804_),
    .X(_11039_));
 sky130_fd_sc_hd__buf_2 _26963_ (.A(_10568_),
    .X(_11040_));
 sky130_fd_sc_hd__nor2_4 _26964_ (.A(_11039_),
    .B(_11040_),
    .Y(_11041_));
 sky130_fd_sc_hd__a2bb2o_2 _26965_ (.A1_N(_11038_),
    .A2_N(_11041_),
    .B1(_11038_),
    .B2(_11041_),
    .X(_11042_));
 sky130_fd_sc_hd__o2bb2ai_4 _26966_ (.A1_N(_11031_),
    .A2_N(_11042_),
    .B1(_11031_),
    .B2(_11042_),
    .Y(_11043_));
 sky130_fd_sc_hd__o22a_2 _26967_ (.A1(_10955_),
    .A2(_10956_),
    .B1(_10957_),
    .B2(_10962_),
    .X(_11044_));
 sky130_fd_sc_hd__o2bb2ai_2 _26968_ (.A1_N(_11043_),
    .A2_N(_11044_),
    .B1(_11043_),
    .B2(_11044_),
    .Y(_11045_));
 sky130_fd_sc_hd__a21oi_4 _26969_ (.A1(_10970_),
    .A2(_10971_),
    .B1(_10969_),
    .Y(_11046_));
 sky130_fd_sc_hd__a21oi_2 _26970_ (.A1(_10960_),
    .A2(_10961_),
    .B1(_10959_),
    .Y(_11047_));
 sky130_fd_sc_hd__clkbuf_2 _26971_ (.A(_10305_),
    .X(_11048_));
 sky130_fd_sc_hd__buf_1 _26972_ (.A(_10367_),
    .X(_11049_));
 sky130_fd_sc_hd__clkbuf_2 _26973_ (.A(_10323_),
    .X(_11050_));
 sky130_fd_sc_hd__o22a_1 _26974_ (.A1(_11049_),
    .A2(_11050_),
    .B1(_07270_),
    .B2(_10751_),
    .X(_11051_));
 sky130_fd_sc_hd__and4_1 _26975_ (.A(_13090_),
    .B(_13512_),
    .C(_13094_),
    .D(_13507_),
    .X(_11052_));
 sky130_fd_sc_hd__or2_1 _26976_ (.A(_11051_),
    .B(_11052_),
    .X(_11053_));
 sky130_vsdinv _26977_ (.A(_11053_),
    .Y(_11054_));
 sky130_fd_sc_hd__or2_1 _26978_ (.A(_11706_),
    .B(_07076_),
    .X(_11055_));
 sky130_fd_sc_hd__buf_1 _26979_ (.A(_11055_),
    .X(_11056_));
 sky130_fd_sc_hd__a32o_1 _26980_ (.A1(_11048_),
    .A2(\pcpi_mul.rs2[24] ),
    .A3(_11054_),
    .B1(_11053_),
    .B2(_11056_),
    .X(_11057_));
 sky130_fd_sc_hd__a2bb2o_1 _26981_ (.A1_N(_11047_),
    .A2_N(_11057_),
    .B1(_11047_),
    .B2(_11057_),
    .X(_11058_));
 sky130_fd_sc_hd__a2bb2o_2 _26982_ (.A1_N(_11046_),
    .A2_N(_11058_),
    .B1(_11046_),
    .B2(_11058_),
    .X(_11059_));
 sky130_fd_sc_hd__o2bb2ai_2 _26983_ (.A1_N(_11045_),
    .A2_N(_11059_),
    .B1(_11045_),
    .B2(_11059_),
    .Y(_11060_));
 sky130_fd_sc_hd__o22a_1 _26984_ (.A1(_10963_),
    .A2(_10964_),
    .B1(_10965_),
    .B2(_10974_),
    .X(_11061_));
 sky130_fd_sc_hd__o2bb2ai_1 _26985_ (.A1_N(_11060_),
    .A2_N(_11061_),
    .B1(_11060_),
    .B2(_11061_),
    .Y(_11062_));
 sky130_fd_sc_hd__buf_1 _26986_ (.A(_10903_),
    .X(_11063_));
 sky130_fd_sc_hd__or2_2 _26987_ (.A(_10333_),
    .B(_10982_),
    .X(_11064_));
 sky130_fd_sc_hd__o21a_1 _26988_ (.A1(_11063_),
    .A2(_10985_),
    .B1(_11064_),
    .X(_11065_));
 sky130_fd_sc_hd__o22a_1 _26989_ (.A1(_10967_),
    .A2(_10972_),
    .B1(_10966_),
    .B2(_10973_),
    .X(_11066_));
 sky130_vsdinv _26990_ (.A(_11064_),
    .Y(_11067_));
 sky130_fd_sc_hd__and2_1 _26991_ (.A(_10829_),
    .B(_10981_),
    .X(_11068_));
 sky130_fd_sc_hd__or2_1 _26992_ (.A(_11067_),
    .B(_11068_),
    .X(_11069_));
 sky130_fd_sc_hd__a2bb2o_1 _26993_ (.A1_N(_11063_),
    .A2_N(_11069_),
    .B1(_10823_),
    .B2(_11069_),
    .X(_11070_));
 sky130_fd_sc_hd__buf_1 _26994_ (.A(_11070_),
    .X(_11071_));
 sky130_fd_sc_hd__buf_1 _26995_ (.A(_11070_),
    .X(_11072_));
 sky130_fd_sc_hd__a2bb2o_1 _26996_ (.A1_N(_11066_),
    .A2_N(_11071_),
    .B1(_11066_),
    .B2(_11072_),
    .X(_11073_));
 sky130_fd_sc_hd__a2bb2o_1 _26997_ (.A1_N(_11065_),
    .A2_N(_11073_),
    .B1(_11065_),
    .B2(_11073_),
    .X(_11074_));
 sky130_fd_sc_hd__o2bb2ai_1 _26998_ (.A1_N(_11062_),
    .A2_N(_11074_),
    .B1(_11062_),
    .B2(_11074_),
    .Y(_11075_));
 sky130_fd_sc_hd__o22a_1 _26999_ (.A1(_10975_),
    .A2(_10976_),
    .B1(_10977_),
    .B2(_10988_),
    .X(_11076_));
 sky130_fd_sc_hd__o2bb2a_1 _27000_ (.A1_N(_11075_),
    .A2_N(_11076_),
    .B1(_11075_),
    .B2(_11076_),
    .X(_11077_));
 sky130_vsdinv _27001_ (.A(_11077_),
    .Y(_11078_));
 sky130_fd_sc_hd__buf_1 _27002_ (.A(_10994_),
    .X(_11079_));
 sky130_fd_sc_hd__buf_1 _27003_ (.A(_11002_),
    .X(_11080_));
 sky130_fd_sc_hd__o22a_1 _27004_ (.A1(_10979_),
    .A2(_10986_),
    .B1(_10978_),
    .B2(_10987_),
    .X(_11081_));
 sky130_fd_sc_hd__a2bb2o_1 _27005_ (.A1_N(_11080_),
    .A2_N(_11081_),
    .B1(_11080_),
    .B2(_11081_),
    .X(_11082_));
 sky130_fd_sc_hd__a2bb2o_1 _27006_ (.A1_N(_11079_),
    .A2_N(_11082_),
    .B1(_11079_),
    .B2(_11082_),
    .X(_11083_));
 sky130_vsdinv _27007_ (.A(_11083_),
    .Y(_11084_));
 sky130_fd_sc_hd__a22o_1 _27008_ (.A1(_11078_),
    .A2(_11083_),
    .B1(_11077_),
    .B2(_11084_),
    .X(_11085_));
 sky130_fd_sc_hd__o22a_1 _27009_ (.A1(_10989_),
    .A2(_10990_),
    .B1(_10992_),
    .B2(_10997_),
    .X(_11086_));
 sky130_fd_sc_hd__a2bb2o_1 _27010_ (.A1_N(_11085_),
    .A2_N(_11086_),
    .B1(_11085_),
    .B2(_11086_),
    .X(_11087_));
 sky130_fd_sc_hd__buf_1 _27011_ (.A(_10683_),
    .X(_11088_));
 sky130_fd_sc_hd__buf_1 _27012_ (.A(_11088_),
    .X(_11089_));
 sky130_fd_sc_hd__buf_1 _27013_ (.A(_10610_),
    .X(_11090_));
 sky130_fd_sc_hd__buf_1 _27014_ (.A(_11090_),
    .X(_11091_));
 sky130_fd_sc_hd__buf_1 _27015_ (.A(_11002_),
    .X(_11092_));
 sky130_fd_sc_hd__buf_1 _27016_ (.A(_10994_),
    .X(_11093_));
 sky130_fd_sc_hd__o22a_1 _27017_ (.A1(_11092_),
    .A2(_10995_),
    .B1(_11093_),
    .B2(_10996_),
    .X(_11094_));
 sky130_fd_sc_hd__a2bb2o_1 _27018_ (.A1_N(_11091_),
    .A2_N(_11094_),
    .B1(_11091_),
    .B2(_11094_),
    .X(_11095_));
 sky130_fd_sc_hd__a2bb2o_1 _27019_ (.A1_N(_11089_),
    .A2_N(_11095_),
    .B1(_11089_),
    .B2(_11095_),
    .X(_11096_));
 sky130_fd_sc_hd__a2bb2o_1 _27020_ (.A1_N(_11087_),
    .A2_N(_11096_),
    .B1(_11087_),
    .B2(_11096_),
    .X(_11097_));
 sky130_fd_sc_hd__o22a_1 _27021_ (.A1(_10999_),
    .A2(_11000_),
    .B1(_11001_),
    .B2(_11005_),
    .X(_11098_));
 sky130_fd_sc_hd__a2bb2o_1 _27022_ (.A1_N(_11097_),
    .A2_N(_11098_),
    .B1(_11097_),
    .B2(_11098_),
    .X(_11099_));
 sky130_fd_sc_hd__buf_1 _27023_ (.A(_10772_),
    .X(_11100_));
 sky130_fd_sc_hd__clkbuf_2 _27024_ (.A(_11100_),
    .X(_11101_));
 sky130_fd_sc_hd__buf_1 _27025_ (.A(_11090_),
    .X(_11102_));
 sky130_fd_sc_hd__buf_1 _27026_ (.A(_11088_),
    .X(_11103_));
 sky130_fd_sc_hd__o22a_1 _27027_ (.A1(_11102_),
    .A2(_11003_),
    .B1(_11103_),
    .B2(_11004_),
    .X(_11104_));
 sky130_fd_sc_hd__buf_1 _27028_ (.A(_10772_),
    .X(_11105_));
 sky130_fd_sc_hd__or2_1 _27029_ (.A(_11105_),
    .B(_11104_),
    .X(_11106_));
 sky130_fd_sc_hd__a21bo_1 _27030_ (.A1(_11101_),
    .A2(_11104_),
    .B1_N(_11106_),
    .X(_11107_));
 sky130_fd_sc_hd__a2bb2o_1 _27031_ (.A1_N(_11099_),
    .A2_N(_11107_),
    .B1(_11099_),
    .B2(_11107_),
    .X(_11108_));
 sky130_fd_sc_hd__o22a_1 _27032_ (.A1(_11006_),
    .A2(_11007_),
    .B1(_11008_),
    .B2(_11011_),
    .X(_11109_));
 sky130_fd_sc_hd__a2bb2o_1 _27033_ (.A1_N(_11108_),
    .A2_N(_11109_),
    .B1(_11108_),
    .B2(_11109_),
    .X(_11110_));
 sky130_fd_sc_hd__a2bb2o_1 _27034_ (.A1_N(_11010_),
    .A2_N(_11110_),
    .B1(_11010_),
    .B2(_11110_),
    .X(_11111_));
 sky130_fd_sc_hd__o22a_1 _27035_ (.A1(_11012_),
    .A2(_11013_),
    .B1(_10940_),
    .B2(_11014_),
    .X(_11112_));
 sky130_fd_sc_hd__or2_1 _27036_ (.A(_11111_),
    .B(_11112_),
    .X(_11113_));
 sky130_fd_sc_hd__a21bo_1 _27037_ (.A1(_11111_),
    .A2(_11112_),
    .B1_N(_11113_),
    .X(_11114_));
 sky130_fd_sc_hd__buf_1 _27038_ (.A(_11114_),
    .X(_11115_));
 sky130_fd_sc_hd__or2_1 _27039_ (.A(_10948_),
    .B(_11019_),
    .X(_11116_));
 sky130_fd_sc_hd__or3_1 _27040_ (.A(_10782_),
    .B(_10871_),
    .C(_11116_),
    .X(_11117_));
 sky130_fd_sc_hd__or2_1 _27041_ (.A(_10785_),
    .B(_11117_),
    .X(_11118_));
 sky130_fd_sc_hd__o221a_1 _27042_ (.A1(_10947_),
    .A2(_11017_),
    .B1(_10949_),
    .B2(_11116_),
    .C1(_11018_),
    .X(_11119_));
 sky130_fd_sc_hd__o221a_2 _27043_ (.A1(_10786_),
    .A2(_11117_),
    .B1(_10406_),
    .B2(_11118_),
    .C1(_11119_),
    .X(_11120_));
 sky130_fd_sc_hd__buf_1 _27044_ (.A(_11120_),
    .X(_11121_));
 sky130_fd_sc_hd__a2bb2oi_1 _27045_ (.A1_N(_11115_),
    .A2_N(_11121_),
    .B1(_11115_),
    .B2(_11121_),
    .Y(_02675_));
 sky130_fd_sc_hd__and4_2 _27046_ (.A(_11021_),
    .B(_10710_),
    .C(_11022_),
    .D(_13531_),
    .X(_11122_));
 sky130_fd_sc_hd__o22a_1 _27047_ (.A1(_11721_),
    .A2(_13537_),
    .B1(_11024_),
    .B2(_10805_),
    .X(_11123_));
 sky130_fd_sc_hd__nor2_2 _27048_ (.A(_11122_),
    .B(_11123_),
    .Y(_11124_));
 sky130_fd_sc_hd__nor2_4 _27049_ (.A(_11027_),
    .B(_11033_),
    .Y(_11125_));
 sky130_fd_sc_hd__a2bb2o_2 _27050_ (.A1_N(_11124_),
    .A2_N(_11125_),
    .B1(_11124_),
    .B2(_11125_),
    .X(_11126_));
 sky130_fd_sc_hd__a21oi_4 _27051_ (.A1(_11026_),
    .A2(_11028_),
    .B1(_11023_),
    .Y(_11127_));
 sky130_fd_sc_hd__o2bb2ai_4 _27052_ (.A1_N(_11126_),
    .A2_N(_11127_),
    .B1(_11126_),
    .B2(_11127_),
    .Y(_11128_));
 sky130_fd_sc_hd__o22a_1 _27053_ (.A1(_11032_),
    .A2(_11035_),
    .B1(_11034_),
    .B2(_10568_),
    .X(_11129_));
 sky130_fd_sc_hd__and4_2 _27054_ (.A(_13077_),
    .B(_13522_),
    .C(_13083_),
    .D(_13517_),
    .X(_11130_));
 sky130_fd_sc_hd__nor2_2 _27055_ (.A(_11129_),
    .B(_11130_),
    .Y(_11131_));
 sky130_fd_sc_hd__buf_2 _27056_ (.A(_11050_),
    .X(_11132_));
 sky130_fd_sc_hd__nor2_4 _27057_ (.A(_11039_),
    .B(_11132_),
    .Y(_11133_));
 sky130_fd_sc_hd__a2bb2o_2 _27058_ (.A1_N(_11131_),
    .A2_N(_11133_),
    .B1(_11131_),
    .B2(_11133_),
    .X(_11134_));
 sky130_fd_sc_hd__o2bb2ai_4 _27059_ (.A1_N(_11128_),
    .A2_N(_11134_),
    .B1(_11128_),
    .B2(_11134_),
    .Y(_11135_));
 sky130_fd_sc_hd__o22a_2 _27060_ (.A1(_11029_),
    .A2(_11030_),
    .B1(_11031_),
    .B2(_11042_),
    .X(_11136_));
 sky130_fd_sc_hd__o2bb2ai_2 _27061_ (.A1_N(_11135_),
    .A2_N(_11136_),
    .B1(_11135_),
    .B2(_11136_),
    .Y(_11137_));
 sky130_fd_sc_hd__buf_1 _27062_ (.A(_11055_),
    .X(_11138_));
 sky130_fd_sc_hd__o21ba_1 _27063_ (.A1(_11053_),
    .A2(_11138_),
    .B1_N(_11052_),
    .X(_11139_));
 sky130_fd_sc_hd__a21oi_4 _27064_ (.A1(_11038_),
    .A2(_11041_),
    .B1(_11037_),
    .Y(_11140_));
 sky130_fd_sc_hd__clkbuf_2 _27065_ (.A(_10751_),
    .X(_11141_));
 sky130_fd_sc_hd__nor2_1 _27066_ (.A(_11049_),
    .B(_11141_),
    .Y(_11142_));
 sky130_fd_sc_hd__or2_2 _27067_ (.A(_10980_),
    .B(_07270_),
    .X(_11143_));
 sky130_vsdinv _27068_ (.A(_11143_),
    .Y(_11144_));
 sky130_fd_sc_hd__a2bb2o_1 _27069_ (.A1_N(_11142_),
    .A2_N(_11144_),
    .B1(_11142_),
    .B2(_11144_),
    .X(_11145_));
 sky130_fd_sc_hd__a2bb2o_1 _27070_ (.A1_N(_11138_),
    .A2_N(_11145_),
    .B1(_11056_),
    .B2(_11145_),
    .X(_11146_));
 sky130_fd_sc_hd__a2bb2o_1 _27071_ (.A1_N(_11140_),
    .A2_N(_11146_),
    .B1(_11140_),
    .B2(_11146_),
    .X(_11147_));
 sky130_fd_sc_hd__a2bb2o_2 _27072_ (.A1_N(_11139_),
    .A2_N(_11147_),
    .B1(_11139_),
    .B2(_11147_),
    .X(_11148_));
 sky130_fd_sc_hd__o2bb2ai_2 _27073_ (.A1_N(_11137_),
    .A2_N(_11148_),
    .B1(_11137_),
    .B2(_11148_),
    .Y(_11149_));
 sky130_fd_sc_hd__o22a_1 _27074_ (.A1(_11043_),
    .A2(_11044_),
    .B1(_11045_),
    .B2(_11059_),
    .X(_11150_));
 sky130_fd_sc_hd__o2bb2ai_1 _27075_ (.A1_N(_11149_),
    .A2_N(_11150_),
    .B1(_11149_),
    .B2(_11150_),
    .Y(_11151_));
 sky130_fd_sc_hd__o21a_1 _27076_ (.A1(_11063_),
    .A2(_11069_),
    .B1(_11064_),
    .X(_11152_));
 sky130_fd_sc_hd__buf_1 _27077_ (.A(_11152_),
    .X(_11153_));
 sky130_fd_sc_hd__o22a_1 _27078_ (.A1(_11047_),
    .A2(_11057_),
    .B1(_11046_),
    .B2(_11058_),
    .X(_11154_));
 sky130_fd_sc_hd__a2bb2o_1 _27079_ (.A1_N(_11072_),
    .A2_N(_11154_),
    .B1(_11072_),
    .B2(_11154_),
    .X(_11155_));
 sky130_fd_sc_hd__a2bb2o_1 _27080_ (.A1_N(_11153_),
    .A2_N(_11155_),
    .B1(_11153_),
    .B2(_11155_),
    .X(_11156_));
 sky130_fd_sc_hd__o2bb2ai_1 _27081_ (.A1_N(_11151_),
    .A2_N(_11156_),
    .B1(_11151_),
    .B2(_11156_),
    .Y(_11157_));
 sky130_fd_sc_hd__o22a_1 _27082_ (.A1(_11060_),
    .A2(_11061_),
    .B1(_11062_),
    .B2(_11074_),
    .X(_11158_));
 sky130_fd_sc_hd__o2bb2a_1 _27083_ (.A1_N(_11157_),
    .A2_N(_11158_),
    .B1(_11157_),
    .B2(_11158_),
    .X(_11159_));
 sky130_vsdinv _27084_ (.A(_11159_),
    .Y(_11160_));
 sky130_fd_sc_hd__buf_1 _27085_ (.A(_11002_),
    .X(_11161_));
 sky130_fd_sc_hd__buf_1 _27086_ (.A(_11071_),
    .X(_11162_));
 sky130_fd_sc_hd__o22a_1 _27087_ (.A1(_11066_),
    .A2(_11162_),
    .B1(_11065_),
    .B2(_11073_),
    .X(_11163_));
 sky130_fd_sc_hd__a2bb2o_1 _27088_ (.A1_N(_11161_),
    .A2_N(_11163_),
    .B1(_11161_),
    .B2(_11163_),
    .X(_11164_));
 sky130_fd_sc_hd__buf_1 _27089_ (.A(_10994_),
    .X(_11165_));
 sky130_fd_sc_hd__a2bb2o_1 _27090_ (.A1_N(_11079_),
    .A2_N(_11164_),
    .B1(_11165_),
    .B2(_11164_),
    .X(_11166_));
 sky130_vsdinv _27091_ (.A(_11166_),
    .Y(_11167_));
 sky130_fd_sc_hd__a22o_1 _27092_ (.A1(_11160_),
    .A2(_11166_),
    .B1(_11159_),
    .B2(_11167_),
    .X(_11168_));
 sky130_fd_sc_hd__o22a_1 _27093_ (.A1(_11075_),
    .A2(_11076_),
    .B1(_11078_),
    .B2(_11083_),
    .X(_11169_));
 sky130_fd_sc_hd__a2bb2o_1 _27094_ (.A1_N(_11168_),
    .A2_N(_11169_),
    .B1(_11168_),
    .B2(_11169_),
    .X(_11170_));
 sky130_fd_sc_hd__buf_1 _27095_ (.A(_11088_),
    .X(_11171_));
 sky130_fd_sc_hd__o22a_1 _27096_ (.A1(_11092_),
    .A2(_11081_),
    .B1(_11093_),
    .B2(_11082_),
    .X(_11172_));
 sky130_fd_sc_hd__a2bb2o_1 _27097_ (.A1_N(_11091_),
    .A2_N(_11172_),
    .B1(_11090_),
    .B2(_11172_),
    .X(_11173_));
 sky130_fd_sc_hd__a2bb2o_1 _27098_ (.A1_N(_11171_),
    .A2_N(_11173_),
    .B1(_11171_),
    .B2(_11173_),
    .X(_11174_));
 sky130_fd_sc_hd__a2bb2o_1 _27099_ (.A1_N(_11170_),
    .A2_N(_11174_),
    .B1(_11170_),
    .B2(_11174_),
    .X(_11175_));
 sky130_fd_sc_hd__o22a_1 _27100_ (.A1(_11085_),
    .A2(_11086_),
    .B1(_11087_),
    .B2(_11096_),
    .X(_11176_));
 sky130_fd_sc_hd__a2bb2o_1 _27101_ (.A1_N(_11175_),
    .A2_N(_11176_),
    .B1(_11175_),
    .B2(_11176_),
    .X(_11177_));
 sky130_fd_sc_hd__o22a_1 _27102_ (.A1(_11102_),
    .A2(_11094_),
    .B1(_11103_),
    .B2(_11095_),
    .X(_11178_));
 sky130_fd_sc_hd__or2_1 _27103_ (.A(_11105_),
    .B(_11178_),
    .X(_11179_));
 sky130_fd_sc_hd__a21bo_1 _27104_ (.A1(_11100_),
    .A2(_11178_),
    .B1_N(_11179_),
    .X(_11180_));
 sky130_fd_sc_hd__a2bb2o_1 _27105_ (.A1_N(_11177_),
    .A2_N(_11180_),
    .B1(_11177_),
    .B2(_11180_),
    .X(_11181_));
 sky130_fd_sc_hd__o22a_1 _27106_ (.A1(_11097_),
    .A2(_11098_),
    .B1(_11099_),
    .B2(_11107_),
    .X(_11182_));
 sky130_fd_sc_hd__a2bb2o_1 _27107_ (.A1_N(_11181_),
    .A2_N(_11182_),
    .B1(_11181_),
    .B2(_11182_),
    .X(_11183_));
 sky130_fd_sc_hd__a2bb2o_1 _27108_ (.A1_N(_11106_),
    .A2_N(_11183_),
    .B1(_11106_),
    .B2(_11183_),
    .X(_11184_));
 sky130_fd_sc_hd__o22a_1 _27109_ (.A1(_11108_),
    .A2(_11109_),
    .B1(_11010_),
    .B2(_11110_),
    .X(_11185_));
 sky130_fd_sc_hd__or2_1 _27110_ (.A(_11184_),
    .B(_11185_),
    .X(_11186_));
 sky130_fd_sc_hd__a21bo_1 _27111_ (.A1(_11184_),
    .A2(_11185_),
    .B1_N(_11186_),
    .X(_11187_));
 sky130_fd_sc_hd__o21ai_1 _27112_ (.A1(_11115_),
    .A2(_11121_),
    .B1(_11113_),
    .Y(_11188_));
 sky130_fd_sc_hd__a2bb2o_1 _27113_ (.A1_N(_11187_),
    .A2_N(_11188_),
    .B1(_11187_),
    .B2(_11188_),
    .X(_02676_));
 sky130_fd_sc_hd__buf_1 _27114_ (.A(_11021_),
    .X(_11189_));
 sky130_fd_sc_hd__and4_2 _27115_ (.A(_11189_),
    .B(_10805_),
    .C(_11022_),
    .D(_13526_),
    .X(_11190_));
 sky130_fd_sc_hd__o22a_1 _27116_ (.A1(_11721_),
    .A2(_13531_),
    .B1(_11024_),
    .B2(_11033_),
    .X(_11191_));
 sky130_fd_sc_hd__nor2_4 _27117_ (.A(_11190_),
    .B(_11191_),
    .Y(_11192_));
 sky130_fd_sc_hd__nor2_4 _27118_ (.A(_11027_),
    .B(_11035_),
    .Y(_11193_));
 sky130_fd_sc_hd__a2bb2o_2 _27119_ (.A1_N(_11192_),
    .A2_N(_11193_),
    .B1(_11192_),
    .B2(_11193_),
    .X(_11194_));
 sky130_fd_sc_hd__a21oi_4 _27120_ (.A1(_11124_),
    .A2(_11125_),
    .B1(_11122_),
    .Y(_11195_));
 sky130_fd_sc_hd__o2bb2ai_2 _27121_ (.A1_N(_11194_),
    .A2_N(_11195_),
    .B1(_11194_),
    .B2(_11195_),
    .Y(_11196_));
 sky130_fd_sc_hd__buf_1 _27122_ (.A(_11032_),
    .X(_11197_));
 sky130_fd_sc_hd__o22a_1 _27123_ (.A1(_11197_),
    .A2(_11040_),
    .B1(_11034_),
    .B2(_11132_),
    .X(_11198_));
 sky130_fd_sc_hd__and4_2 _27124_ (.A(_13077_),
    .B(_13518_),
    .C(_13083_),
    .D(_13513_),
    .X(_11199_));
 sky130_fd_sc_hd__nor2_2 _27125_ (.A(_11198_),
    .B(_11199_),
    .Y(_11200_));
 sky130_fd_sc_hd__nor2_2 _27126_ (.A(_11039_),
    .B(_11141_),
    .Y(_11201_));
 sky130_fd_sc_hd__a2bb2o_2 _27127_ (.A1_N(_11200_),
    .A2_N(_11201_),
    .B1(_11200_),
    .B2(_11201_),
    .X(_11202_));
 sky130_fd_sc_hd__o2bb2ai_2 _27128_ (.A1_N(_11196_),
    .A2_N(_11202_),
    .B1(_11196_),
    .B2(_11202_),
    .Y(_11203_));
 sky130_fd_sc_hd__o22a_2 _27129_ (.A1(_11126_),
    .A2(_11127_),
    .B1(_11128_),
    .B2(_11134_),
    .X(_11204_));
 sky130_fd_sc_hd__o2bb2ai_2 _27130_ (.A1_N(_11203_),
    .A2_N(_11204_),
    .B1(_11203_),
    .B2(_11204_),
    .Y(_11205_));
 sky130_fd_sc_hd__clkbuf_2 _27131_ (.A(_11141_),
    .X(_11206_));
 sky130_fd_sc_hd__o32a_1 _27132_ (.A1(_11049_),
    .A2(_11206_),
    .A3(_11143_),
    .B1(_11138_),
    .B2(_11145_),
    .X(_11207_));
 sky130_fd_sc_hd__a21oi_4 _27133_ (.A1(_11131_),
    .A2(_11133_),
    .B1(_11130_),
    .Y(_11208_));
 sky130_fd_sc_hd__or2_1 _27134_ (.A(_10980_),
    .B(_11049_),
    .X(_11209_));
 sky130_fd_sc_hd__a32o_1 _27135_ (.A1(_11048_),
    .A2(_13090_),
    .A3(_11144_),
    .B1(_11143_),
    .B2(_11209_),
    .X(_11210_));
 sky130_fd_sc_hd__a2bb2o_1 _27136_ (.A1_N(_11056_),
    .A2_N(_11210_),
    .B1(_11056_),
    .B2(_11210_),
    .X(_11211_));
 sky130_fd_sc_hd__buf_1 _27137_ (.A(_11211_),
    .X(_11212_));
 sky130_fd_sc_hd__a2bb2o_1 _27138_ (.A1_N(_11208_),
    .A2_N(_11212_),
    .B1(_11208_),
    .B2(_11211_),
    .X(_11213_));
 sky130_fd_sc_hd__a2bb2o_2 _27139_ (.A1_N(_11207_),
    .A2_N(_11213_),
    .B1(_11207_),
    .B2(_11213_),
    .X(_11214_));
 sky130_fd_sc_hd__o2bb2ai_2 _27140_ (.A1_N(_11205_),
    .A2_N(_11214_),
    .B1(_11205_),
    .B2(_11214_),
    .Y(_11215_));
 sky130_fd_sc_hd__o22a_1 _27141_ (.A1(_11135_),
    .A2(_11136_),
    .B1(_11137_),
    .B2(_11148_),
    .X(_11216_));
 sky130_fd_sc_hd__o2bb2ai_1 _27142_ (.A1_N(_11215_),
    .A2_N(_11216_),
    .B1(_11215_),
    .B2(_11216_),
    .Y(_11217_));
 sky130_fd_sc_hd__buf_1 _27143_ (.A(_11152_),
    .X(_11218_));
 sky130_fd_sc_hd__o22a_1 _27144_ (.A1(_11140_),
    .A2(_11146_),
    .B1(_11139_),
    .B2(_11147_),
    .X(_11219_));
 sky130_fd_sc_hd__a2bb2o_1 _27145_ (.A1_N(_11071_),
    .A2_N(_11219_),
    .B1(_11071_),
    .B2(_11219_),
    .X(_11220_));
 sky130_fd_sc_hd__a2bb2o_1 _27146_ (.A1_N(_11218_),
    .A2_N(_11220_),
    .B1(_11153_),
    .B2(_11220_),
    .X(_11221_));
 sky130_fd_sc_hd__o2bb2ai_1 _27147_ (.A1_N(_11217_),
    .A2_N(_11221_),
    .B1(_11217_),
    .B2(_11221_),
    .Y(_11222_));
 sky130_fd_sc_hd__o22a_1 _27148_ (.A1(_11149_),
    .A2(_11150_),
    .B1(_11151_),
    .B2(_11156_),
    .X(_11223_));
 sky130_fd_sc_hd__o2bb2a_1 _27149_ (.A1_N(_11222_),
    .A2_N(_11223_),
    .B1(_11222_),
    .B2(_11223_),
    .X(_11224_));
 sky130_vsdinv _27150_ (.A(_11224_),
    .Y(_11225_));
 sky130_fd_sc_hd__buf_1 _27151_ (.A(_11072_),
    .X(_11226_));
 sky130_fd_sc_hd__o22a_1 _27152_ (.A1(_11226_),
    .A2(_11154_),
    .B1(_11218_),
    .B2(_11155_),
    .X(_11227_));
 sky130_fd_sc_hd__a2bb2o_1 _27153_ (.A1_N(_11161_),
    .A2_N(_11227_),
    .B1(_11161_),
    .B2(_11227_),
    .X(_11228_));
 sky130_fd_sc_hd__a2bb2o_1 _27154_ (.A1_N(_11165_),
    .A2_N(_11228_),
    .B1(_11165_),
    .B2(_11228_),
    .X(_11229_));
 sky130_vsdinv _27155_ (.A(_11229_),
    .Y(_11230_));
 sky130_fd_sc_hd__a22o_1 _27156_ (.A1(_11225_),
    .A2(_11229_),
    .B1(_11224_),
    .B2(_11230_),
    .X(_11231_));
 sky130_fd_sc_hd__o22a_1 _27157_ (.A1(_11157_),
    .A2(_11158_),
    .B1(_11160_),
    .B2(_11166_),
    .X(_11232_));
 sky130_fd_sc_hd__a2bb2o_1 _27158_ (.A1_N(_11231_),
    .A2_N(_11232_),
    .B1(_11231_),
    .B2(_11232_),
    .X(_11233_));
 sky130_fd_sc_hd__buf_1 _27159_ (.A(_11090_),
    .X(_11234_));
 sky130_fd_sc_hd__buf_1 _27160_ (.A(_11092_),
    .X(_11235_));
 sky130_fd_sc_hd__o22a_1 _27161_ (.A1(_11235_),
    .A2(_11163_),
    .B1(_11093_),
    .B2(_11164_),
    .X(_11236_));
 sky130_fd_sc_hd__a2bb2o_1 _27162_ (.A1_N(_11234_),
    .A2_N(_11236_),
    .B1(_11091_),
    .B2(_11236_),
    .X(_11237_));
 sky130_fd_sc_hd__a2bb2o_1 _27163_ (.A1_N(_11171_),
    .A2_N(_11237_),
    .B1(_11171_),
    .B2(_11237_),
    .X(_11238_));
 sky130_fd_sc_hd__a2bb2o_1 _27164_ (.A1_N(_11233_),
    .A2_N(_11238_),
    .B1(_11233_),
    .B2(_11238_),
    .X(_11239_));
 sky130_fd_sc_hd__o22a_1 _27165_ (.A1(_11168_),
    .A2(_11169_),
    .B1(_11170_),
    .B2(_11174_),
    .X(_11240_));
 sky130_fd_sc_hd__a2bb2o_1 _27166_ (.A1_N(_11239_),
    .A2_N(_11240_),
    .B1(_11239_),
    .B2(_11240_),
    .X(_11241_));
 sky130_fd_sc_hd__o22a_1 _27167_ (.A1(_11102_),
    .A2(_11172_),
    .B1(_11088_),
    .B2(_11173_),
    .X(_11242_));
 sky130_fd_sc_hd__or2_1 _27168_ (.A(_11105_),
    .B(_11242_),
    .X(_11243_));
 sky130_fd_sc_hd__a21bo_1 _27169_ (.A1(_11100_),
    .A2(_11242_),
    .B1_N(_11243_),
    .X(_11244_));
 sky130_fd_sc_hd__a2bb2o_1 _27170_ (.A1_N(_11241_),
    .A2_N(_11244_),
    .B1(_11241_),
    .B2(_11244_),
    .X(_11245_));
 sky130_fd_sc_hd__o22a_1 _27171_ (.A1(_11175_),
    .A2(_11176_),
    .B1(_11177_),
    .B2(_11180_),
    .X(_11246_));
 sky130_fd_sc_hd__a2bb2o_1 _27172_ (.A1_N(_11245_),
    .A2_N(_11246_),
    .B1(_11245_),
    .B2(_11246_),
    .X(_11247_));
 sky130_fd_sc_hd__a2bb2o_1 _27173_ (.A1_N(_11179_),
    .A2_N(_11247_),
    .B1(_11179_),
    .B2(_11247_),
    .X(_11248_));
 sky130_fd_sc_hd__o22a_1 _27174_ (.A1(_11181_),
    .A2(_11182_),
    .B1(_11106_),
    .B2(_11183_),
    .X(_11249_));
 sky130_fd_sc_hd__or2_1 _27175_ (.A(_11248_),
    .B(_11249_),
    .X(_11250_));
 sky130_fd_sc_hd__a21bo_1 _27176_ (.A1(_11248_),
    .A2(_11249_),
    .B1_N(_11250_),
    .X(_11251_));
 sky130_fd_sc_hd__a22o_1 _27177_ (.A1(_11184_),
    .A2(_11185_),
    .B1(_11113_),
    .B2(_11186_),
    .X(_11252_));
 sky130_fd_sc_hd__o31a_1 _27178_ (.A1(_11115_),
    .A2(_11187_),
    .A3(_11121_),
    .B1(_11252_),
    .X(_11253_));
 sky130_fd_sc_hd__a2bb2oi_1 _27179_ (.A1_N(_11251_),
    .A2_N(_11253_),
    .B1(_11251_),
    .B2(_11253_),
    .Y(_02677_));
 sky130_fd_sc_hd__and4_2 _27180_ (.A(_11189_),
    .B(_11033_),
    .C(_13068_),
    .D(_13521_),
    .X(_11254_));
 sky130_fd_sc_hd__buf_1 _27181_ (.A(_10873_),
    .X(_11255_));
 sky130_fd_sc_hd__o22a_1 _27182_ (.A1(_11721_),
    .A2(_13526_),
    .B1(_11255_),
    .B2(_10489_),
    .X(_11256_));
 sky130_fd_sc_hd__nor2_2 _27183_ (.A(_11254_),
    .B(_11256_),
    .Y(_11257_));
 sky130_fd_sc_hd__buf_2 _27184_ (.A(_11027_),
    .X(_11258_));
 sky130_fd_sc_hd__nor2_4 _27185_ (.A(_11258_),
    .B(_11040_),
    .Y(_11259_));
 sky130_fd_sc_hd__a2bb2o_2 _27186_ (.A1_N(_11257_),
    .A2_N(_11259_),
    .B1(_11257_),
    .B2(_11259_),
    .X(_11260_));
 sky130_fd_sc_hd__a21oi_4 _27187_ (.A1(_11192_),
    .A2(_11193_),
    .B1(_11190_),
    .Y(_11261_));
 sky130_fd_sc_hd__o2bb2ai_4 _27188_ (.A1_N(_11260_),
    .A2_N(_11261_),
    .B1(_11260_),
    .B2(_11261_),
    .Y(_11262_));
 sky130_fd_sc_hd__buf_1 _27189_ (.A(_11048_),
    .X(_11263_));
 sky130_fd_sc_hd__o22a_1 _27190_ (.A1(_11032_),
    .A2(_11050_),
    .B1(_11034_),
    .B2(_11141_),
    .X(_11264_));
 sky130_fd_sc_hd__and4_1 _27191_ (.A(_13076_),
    .B(_13513_),
    .C(_13082_),
    .D(_13508_),
    .X(_11265_));
 sky130_fd_sc_hd__or2_1 _27192_ (.A(_11264_),
    .B(_11265_),
    .X(_11266_));
 sky130_vsdinv _27193_ (.A(_11266_),
    .Y(_11267_));
 sky130_fd_sc_hd__or2_1 _27194_ (.A(_11707_),
    .B(_11039_),
    .X(_11268_));
 sky130_fd_sc_hd__a32o_2 _27195_ (.A1(_11263_),
    .A2(\pcpi_mul.rs2[27] ),
    .A3(_11267_),
    .B1(_11266_),
    .B2(_11268_),
    .X(_11269_));
 sky130_fd_sc_hd__o2bb2ai_4 _27196_ (.A1_N(_11262_),
    .A2_N(_11269_),
    .B1(_11262_),
    .B2(_11269_),
    .Y(_11270_));
 sky130_fd_sc_hd__o22a_2 _27197_ (.A1(_11194_),
    .A2(_11195_),
    .B1(_11196_),
    .B2(_11202_),
    .X(_11271_));
 sky130_fd_sc_hd__o2bb2ai_2 _27198_ (.A1_N(_11270_),
    .A2_N(_11271_),
    .B1(_11270_),
    .B2(_11271_),
    .Y(_11272_));
 sky130_fd_sc_hd__o22a_1 _27199_ (.A1(_11143_),
    .A2(_11209_),
    .B1(_11138_),
    .B2(_11210_),
    .X(_11273_));
 sky130_fd_sc_hd__a21oi_2 _27200_ (.A1(_11200_),
    .A2(_11201_),
    .B1(_11199_),
    .Y(_11274_));
 sky130_fd_sc_hd__a2bb2o_1 _27201_ (.A1_N(_11212_),
    .A2_N(_11274_),
    .B1(_11212_),
    .B2(_11274_),
    .X(_11275_));
 sky130_fd_sc_hd__a2bb2o_2 _27202_ (.A1_N(_11273_),
    .A2_N(_11275_),
    .B1(_11273_),
    .B2(_11275_),
    .X(_11276_));
 sky130_fd_sc_hd__o2bb2ai_2 _27203_ (.A1_N(_11272_),
    .A2_N(_11276_),
    .B1(_11272_),
    .B2(_11276_),
    .Y(_11277_));
 sky130_fd_sc_hd__o22a_1 _27204_ (.A1(_11203_),
    .A2(_11204_),
    .B1(_11205_),
    .B2(_11214_),
    .X(_11278_));
 sky130_fd_sc_hd__o2bb2ai_1 _27205_ (.A1_N(_11277_),
    .A2_N(_11278_),
    .B1(_11277_),
    .B2(_11278_),
    .Y(_11279_));
 sky130_fd_sc_hd__buf_1 _27206_ (.A(_11153_),
    .X(_11280_));
 sky130_fd_sc_hd__buf_1 _27207_ (.A(_11211_),
    .X(_11281_));
 sky130_fd_sc_hd__o22a_1 _27208_ (.A1(_11208_),
    .A2(_11281_),
    .B1(_11207_),
    .B2(_11213_),
    .X(_11282_));
 sky130_fd_sc_hd__a2bb2o_1 _27209_ (.A1_N(_11226_),
    .A2_N(_11282_),
    .B1(_11226_),
    .B2(_11282_),
    .X(_11283_));
 sky130_fd_sc_hd__a2bb2o_1 _27210_ (.A1_N(_11280_),
    .A2_N(_11283_),
    .B1(_11218_),
    .B2(_11283_),
    .X(_11284_));
 sky130_fd_sc_hd__o2bb2ai_1 _27211_ (.A1_N(_11279_),
    .A2_N(_11284_),
    .B1(_11279_),
    .B2(_11284_),
    .Y(_11285_));
 sky130_fd_sc_hd__o22a_1 _27212_ (.A1(_11215_),
    .A2(_11216_),
    .B1(_11217_),
    .B2(_11221_),
    .X(_11286_));
 sky130_fd_sc_hd__o2bb2a_1 _27213_ (.A1_N(_11285_),
    .A2_N(_11286_),
    .B1(_11285_),
    .B2(_11286_),
    .X(_11287_));
 sky130_vsdinv _27214_ (.A(_11287_),
    .Y(_11288_));
 sky130_fd_sc_hd__o22a_1 _27215_ (.A1(_11162_),
    .A2(_11219_),
    .B1(_11218_),
    .B2(_11220_),
    .X(_11289_));
 sky130_fd_sc_hd__a2bb2o_1 _27216_ (.A1_N(_11080_),
    .A2_N(_11289_),
    .B1(_11080_),
    .B2(_11289_),
    .X(_11290_));
 sky130_fd_sc_hd__a2bb2o_1 _27217_ (.A1_N(_11093_),
    .A2_N(_11290_),
    .B1(_11079_),
    .B2(_11290_),
    .X(_11291_));
 sky130_vsdinv _27218_ (.A(_11291_),
    .Y(_11292_));
 sky130_fd_sc_hd__a22o_1 _27219_ (.A1(_11288_),
    .A2(_11291_),
    .B1(_11287_),
    .B2(_11292_),
    .X(_11293_));
 sky130_fd_sc_hd__o22a_1 _27220_ (.A1(_11222_),
    .A2(_11223_),
    .B1(_11225_),
    .B2(_11229_),
    .X(_11294_));
 sky130_fd_sc_hd__a2bb2o_1 _27221_ (.A1_N(_11293_),
    .A2_N(_11294_),
    .B1(_11293_),
    .B2(_11294_),
    .X(_11295_));
 sky130_fd_sc_hd__buf_1 _27222_ (.A(_11165_),
    .X(_11296_));
 sky130_fd_sc_hd__o22a_1 _27223_ (.A1(_11235_),
    .A2(_11227_),
    .B1(_11296_),
    .B2(_11228_),
    .X(_11297_));
 sky130_fd_sc_hd__a2bb2o_1 _27224_ (.A1_N(_11234_),
    .A2_N(_11297_),
    .B1(_11234_),
    .B2(_11297_),
    .X(_11298_));
 sky130_fd_sc_hd__a2bb2o_1 _27225_ (.A1_N(_11089_),
    .A2_N(_11298_),
    .B1(_11089_),
    .B2(_11298_),
    .X(_11299_));
 sky130_fd_sc_hd__a2bb2o_1 _27226_ (.A1_N(_11295_),
    .A2_N(_11299_),
    .B1(_11295_),
    .B2(_11299_),
    .X(_11300_));
 sky130_fd_sc_hd__o22a_1 _27227_ (.A1(_11231_),
    .A2(_11232_),
    .B1(_11233_),
    .B2(_11238_),
    .X(_11301_));
 sky130_fd_sc_hd__a2bb2o_1 _27228_ (.A1_N(_11300_),
    .A2_N(_11301_),
    .B1(_11300_),
    .B2(_11301_),
    .X(_11302_));
 sky130_fd_sc_hd__o22a_1 _27229_ (.A1(_11102_),
    .A2(_11236_),
    .B1(_11103_),
    .B2(_11237_),
    .X(_11303_));
 sky130_fd_sc_hd__or2_1 _27230_ (.A(_11105_),
    .B(_11303_),
    .X(_11304_));
 sky130_fd_sc_hd__a21bo_1 _27231_ (.A1(_11100_),
    .A2(_11303_),
    .B1_N(_11304_),
    .X(_11305_));
 sky130_fd_sc_hd__a2bb2o_1 _27232_ (.A1_N(_11302_),
    .A2_N(_11305_),
    .B1(_11302_),
    .B2(_11305_),
    .X(_11306_));
 sky130_fd_sc_hd__o22a_1 _27233_ (.A1(_11239_),
    .A2(_11240_),
    .B1(_11241_),
    .B2(_11244_),
    .X(_11307_));
 sky130_fd_sc_hd__a2bb2o_1 _27234_ (.A1_N(_11306_),
    .A2_N(_11307_),
    .B1(_11306_),
    .B2(_11307_),
    .X(_11308_));
 sky130_fd_sc_hd__a2bb2o_1 _27235_ (.A1_N(_11243_),
    .A2_N(_11308_),
    .B1(_11243_),
    .B2(_11308_),
    .X(_11309_));
 sky130_fd_sc_hd__o22a_1 _27236_ (.A1(_11245_),
    .A2(_11246_),
    .B1(_11179_),
    .B2(_11247_),
    .X(_11310_));
 sky130_fd_sc_hd__and2_1 _27237_ (.A(_11309_),
    .B(_11310_),
    .X(_11311_));
 sky130_fd_sc_hd__or2_1 _27238_ (.A(_11309_),
    .B(_11310_),
    .X(_11312_));
 sky130_fd_sc_hd__or2b_1 _27239_ (.A(_11311_),
    .B_N(_11312_),
    .X(_11313_));
 sky130_fd_sc_hd__o21ai_1 _27240_ (.A1(_11251_),
    .A2(_11253_),
    .B1(_11250_),
    .Y(_11314_));
 sky130_fd_sc_hd__a2bb2o_1 _27241_ (.A1_N(_11313_),
    .A2_N(_11314_),
    .B1(_11313_),
    .B2(_11314_),
    .X(_02678_));
 sky130_fd_sc_hd__and4_2 _27242_ (.A(_11189_),
    .B(_11035_),
    .C(_13068_),
    .D(_13518_),
    .X(_11315_));
 sky130_fd_sc_hd__o22a_1 _27243_ (.A1(_11722_),
    .A2(_13522_),
    .B1(_11255_),
    .B2(_11040_),
    .X(_11316_));
 sky130_fd_sc_hd__nor2_2 _27244_ (.A(_11315_),
    .B(_11316_),
    .Y(_11317_));
 sky130_fd_sc_hd__nor2_4 _27245_ (.A(_11258_),
    .B(_11132_),
    .Y(_11318_));
 sky130_fd_sc_hd__a2bb2o_2 _27246_ (.A1_N(_11317_),
    .A2_N(_11318_),
    .B1(_11317_),
    .B2(_11318_),
    .X(_11319_));
 sky130_fd_sc_hd__a21oi_4 _27247_ (.A1(_11257_),
    .A2(_11259_),
    .B1(_11254_),
    .Y(_11320_));
 sky130_fd_sc_hd__o2bb2ai_2 _27248_ (.A1_N(_11319_),
    .A2_N(_11320_),
    .B1(_11319_),
    .B2(_11320_),
    .Y(_11321_));
 sky130_fd_sc_hd__buf_1 _27249_ (.A(_11268_),
    .X(_11322_));
 sky130_fd_sc_hd__buf_1 _27250_ (.A(_11322_),
    .X(_11323_));
 sky130_fd_sc_hd__nor2_1 _27251_ (.A(_11197_),
    .B(_11206_),
    .Y(_11324_));
 sky130_fd_sc_hd__or2_2 _27252_ (.A(_11706_),
    .B(_10880_),
    .X(_11325_));
 sky130_vsdinv _27253_ (.A(_11325_),
    .Y(_11326_));
 sky130_fd_sc_hd__a2bb2o_1 _27254_ (.A1_N(_11324_),
    .A2_N(_11326_),
    .B1(_11324_),
    .B2(_11326_),
    .X(_11327_));
 sky130_fd_sc_hd__a2bb2o_2 _27255_ (.A1_N(_11323_),
    .A2_N(_11327_),
    .B1(_11323_),
    .B2(_11327_),
    .X(_11328_));
 sky130_fd_sc_hd__o2bb2ai_2 _27256_ (.A1_N(_11321_),
    .A2_N(_11328_),
    .B1(_11321_),
    .B2(_11328_),
    .Y(_11329_));
 sky130_fd_sc_hd__o22a_2 _27257_ (.A1(_11260_),
    .A2(_11261_),
    .B1(_11262_),
    .B2(_11269_),
    .X(_11330_));
 sky130_fd_sc_hd__o2bb2ai_1 _27258_ (.A1_N(_11329_),
    .A2_N(_11330_),
    .B1(_11329_),
    .B2(_11330_),
    .Y(_11331_));
 sky130_fd_sc_hd__buf_1 _27259_ (.A(_11273_),
    .X(_11332_));
 sky130_fd_sc_hd__buf_1 _27260_ (.A(_11332_),
    .X(_11333_));
 sky130_fd_sc_hd__buf_1 _27261_ (.A(_11212_),
    .X(_11334_));
 sky130_fd_sc_hd__o21ba_1 _27262_ (.A1(_11266_),
    .A2(_11323_),
    .B1_N(_11265_),
    .X(_11335_));
 sky130_fd_sc_hd__a2bb2o_1 _27263_ (.A1_N(_11334_),
    .A2_N(_11335_),
    .B1(_11334_),
    .B2(_11335_),
    .X(_11336_));
 sky130_fd_sc_hd__a2bb2o_1 _27264_ (.A1_N(_11333_),
    .A2_N(_11336_),
    .B1(_11333_),
    .B2(_11336_),
    .X(_11337_));
 sky130_fd_sc_hd__o2bb2ai_1 _27265_ (.A1_N(_11331_),
    .A2_N(_11337_),
    .B1(_11331_),
    .B2(_11337_),
    .Y(_11338_));
 sky130_fd_sc_hd__o22a_1 _27266_ (.A1(_11270_),
    .A2(_11271_),
    .B1(_11272_),
    .B2(_11276_),
    .X(_11339_));
 sky130_fd_sc_hd__o2bb2ai_1 _27267_ (.A1_N(_11338_),
    .A2_N(_11339_),
    .B1(_11338_),
    .B2(_11339_),
    .Y(_11340_));
 sky130_fd_sc_hd__buf_1 _27268_ (.A(_11280_),
    .X(_11341_));
 sky130_fd_sc_hd__buf_1 _27269_ (.A(_11226_),
    .X(_11342_));
 sky130_fd_sc_hd__buf_1 _27270_ (.A(_11281_),
    .X(_11343_));
 sky130_fd_sc_hd__o22a_1 _27271_ (.A1(_11343_),
    .A2(_11274_),
    .B1(_11332_),
    .B2(_11275_),
    .X(_11344_));
 sky130_fd_sc_hd__a2bb2o_1 _27272_ (.A1_N(_11342_),
    .A2_N(_11344_),
    .B1(_11162_),
    .B2(_11344_),
    .X(_11345_));
 sky130_fd_sc_hd__a2bb2o_1 _27273_ (.A1_N(_11341_),
    .A2_N(_11345_),
    .B1(_11280_),
    .B2(_11345_),
    .X(_11346_));
 sky130_fd_sc_hd__o2bb2ai_1 _27274_ (.A1_N(_11340_),
    .A2_N(_11346_),
    .B1(_11340_),
    .B2(_11346_),
    .Y(_11347_));
 sky130_fd_sc_hd__o22a_1 _27275_ (.A1(_11277_),
    .A2(_11278_),
    .B1(_11279_),
    .B2(_11284_),
    .X(_11348_));
 sky130_fd_sc_hd__o2bb2a_1 _27276_ (.A1_N(_11347_),
    .A2_N(_11348_),
    .B1(_11347_),
    .B2(_11348_),
    .X(_11349_));
 sky130_vsdinv _27277_ (.A(_11349_),
    .Y(_11350_));
 sky130_fd_sc_hd__buf_1 _27278_ (.A(_11296_),
    .X(_11351_));
 sky130_fd_sc_hd__buf_1 _27279_ (.A(_11092_),
    .X(_11352_));
 sky130_fd_sc_hd__buf_1 _27280_ (.A(_11162_),
    .X(_11353_));
 sky130_fd_sc_hd__buf_1 _27281_ (.A(_11280_),
    .X(_11354_));
 sky130_fd_sc_hd__o22a_1 _27282_ (.A1(_11353_),
    .A2(_11282_),
    .B1(_11354_),
    .B2(_11283_),
    .X(_11355_));
 sky130_fd_sc_hd__a2bb2o_1 _27283_ (.A1_N(_11352_),
    .A2_N(_11355_),
    .B1(_11352_),
    .B2(_11355_),
    .X(_11356_));
 sky130_fd_sc_hd__a2bb2o_1 _27284_ (.A1_N(_11351_),
    .A2_N(_11356_),
    .B1(_11351_),
    .B2(_11356_),
    .X(_11357_));
 sky130_vsdinv _27285_ (.A(_11357_),
    .Y(_11358_));
 sky130_fd_sc_hd__a22o_1 _27286_ (.A1(_11350_),
    .A2(_11357_),
    .B1(_11349_),
    .B2(_11358_),
    .X(_11359_));
 sky130_fd_sc_hd__o22a_1 _27287_ (.A1(_11285_),
    .A2(_11286_),
    .B1(_11288_),
    .B2(_11291_),
    .X(_11360_));
 sky130_fd_sc_hd__a2bb2o_1 _27288_ (.A1_N(_11359_),
    .A2_N(_11360_),
    .B1(_11359_),
    .B2(_11360_),
    .X(_11361_));
 sky130_fd_sc_hd__buf_1 _27289_ (.A(_11103_),
    .X(_11362_));
 sky130_fd_sc_hd__buf_1 _27290_ (.A(_11362_),
    .X(_11363_));
 sky130_fd_sc_hd__buf_1 _27291_ (.A(_11234_),
    .X(_11364_));
 sky130_fd_sc_hd__buf_1 _27292_ (.A(_11235_),
    .X(_11365_));
 sky130_fd_sc_hd__o22a_1 _27293_ (.A1(_11365_),
    .A2(_11289_),
    .B1(_11351_),
    .B2(_11290_),
    .X(_11366_));
 sky130_fd_sc_hd__a2bb2o_1 _27294_ (.A1_N(_11364_),
    .A2_N(_11366_),
    .B1(_11364_),
    .B2(_11366_),
    .X(_11367_));
 sky130_fd_sc_hd__buf_1 _27295_ (.A(_11362_),
    .X(_11368_));
 sky130_fd_sc_hd__a2bb2o_1 _27296_ (.A1_N(_11363_),
    .A2_N(_11367_),
    .B1(_11368_),
    .B2(_11367_),
    .X(_11369_));
 sky130_fd_sc_hd__a2bb2o_1 _27297_ (.A1_N(_11361_),
    .A2_N(_11369_),
    .B1(_11361_),
    .B2(_11369_),
    .X(_11370_));
 sky130_fd_sc_hd__o22a_1 _27298_ (.A1(_11293_),
    .A2(_11294_),
    .B1(_11295_),
    .B2(_11299_),
    .X(_11371_));
 sky130_fd_sc_hd__a2bb2o_1 _27299_ (.A1_N(_11370_),
    .A2_N(_11371_),
    .B1(_11370_),
    .B2(_11371_),
    .X(_11372_));
 sky130_fd_sc_hd__buf_1 _27300_ (.A(_11101_),
    .X(_11373_));
 sky130_fd_sc_hd__buf_1 _27301_ (.A(_11364_),
    .X(_11374_));
 sky130_fd_sc_hd__o22a_1 _27302_ (.A1(_11374_),
    .A2(_11297_),
    .B1(_11363_),
    .B2(_11298_),
    .X(_11375_));
 sky130_fd_sc_hd__or2_1 _27303_ (.A(_11373_),
    .B(_11375_),
    .X(_11376_));
 sky130_fd_sc_hd__a21bo_1 _27304_ (.A1(_11373_),
    .A2(_11375_),
    .B1_N(_11376_),
    .X(_11377_));
 sky130_fd_sc_hd__a2bb2o_1 _27305_ (.A1_N(_11372_),
    .A2_N(_11377_),
    .B1(_11372_),
    .B2(_11377_),
    .X(_11378_));
 sky130_fd_sc_hd__o22a_1 _27306_ (.A1(_11300_),
    .A2(_11301_),
    .B1(_11302_),
    .B2(_11305_),
    .X(_11379_));
 sky130_fd_sc_hd__a2bb2o_1 _27307_ (.A1_N(_11378_),
    .A2_N(_11379_),
    .B1(_11378_),
    .B2(_11379_),
    .X(_11380_));
 sky130_fd_sc_hd__a2bb2o_1 _27308_ (.A1_N(_11304_),
    .A2_N(_11380_),
    .B1(_11304_),
    .B2(_11380_),
    .X(_11381_));
 sky130_fd_sc_hd__o22a_1 _27309_ (.A1(_11306_),
    .A2(_11307_),
    .B1(_11243_),
    .B2(_11308_),
    .X(_11382_));
 sky130_fd_sc_hd__or2_1 _27310_ (.A(_11381_),
    .B(_11382_),
    .X(_11383_));
 sky130_vsdinv _27311_ (.A(_11383_),
    .Y(_11384_));
 sky130_fd_sc_hd__a21oi_4 _27312_ (.A1(_11381_),
    .A2(_11382_),
    .B1(_11384_),
    .Y(_11385_));
 sky130_vsdinv _27313_ (.A(_11385_),
    .Y(_11386_));
 sky130_fd_sc_hd__or2_1 _27314_ (.A(_11251_),
    .B(_11313_),
    .X(_11387_));
 sky130_fd_sc_hd__o221a_1 _27315_ (.A1(_11250_),
    .A2(_11311_),
    .B1(_11252_),
    .B2(_11387_),
    .C1(_11312_),
    .X(_11388_));
 sky130_fd_sc_hd__o41a_2 _27316_ (.A1(_11114_),
    .A2(_11187_),
    .A3(_11387_),
    .A4(_11120_),
    .B1(_11388_),
    .X(_11389_));
 sky130_vsdinv _27317_ (.A(_11389_),
    .Y(_11390_));
 sky130_fd_sc_hd__o22a_1 _27318_ (.A1(_11386_),
    .A2(_11389_),
    .B1(_11385_),
    .B2(_11390_),
    .X(_02679_));
 sky130_fd_sc_hd__and4_1 _27319_ (.A(_11189_),
    .B(_10568_),
    .C(_13068_),
    .D(_13513_),
    .X(_11391_));
 sky130_fd_sc_hd__o22a_1 _27320_ (.A1(_11722_),
    .A2(_13518_),
    .B1(_11255_),
    .B2(_11132_),
    .X(_11392_));
 sky130_fd_sc_hd__nor2_2 _27321_ (.A(_11391_),
    .B(_11392_),
    .Y(_11393_));
 sky130_fd_sc_hd__nor2_1 _27322_ (.A(_11258_),
    .B(_11206_),
    .Y(_11394_));
 sky130_fd_sc_hd__a2bb2o_2 _27323_ (.A1_N(_11393_),
    .A2_N(_11394_),
    .B1(_11393_),
    .B2(_11394_),
    .X(_11395_));
 sky130_fd_sc_hd__a21oi_4 _27324_ (.A1(_11317_),
    .A2(_11318_),
    .B1(_11315_),
    .Y(_11396_));
 sky130_fd_sc_hd__o2bb2ai_2 _27325_ (.A1_N(_11395_),
    .A2_N(_11396_),
    .B1(_11395_),
    .B2(_11396_),
    .Y(_11397_));
 sky130_fd_sc_hd__or2_1 _27326_ (.A(_11706_),
    .B(_11197_),
    .X(_11398_));
 sky130_fd_sc_hd__a32o_1 _27327_ (.A1(_11048_),
    .A2(_13077_),
    .A3(_11326_),
    .B1(_11325_),
    .B2(_11398_),
    .X(_11399_));
 sky130_fd_sc_hd__a2bb2o_1 _27328_ (.A1_N(_11322_),
    .A2_N(_11399_),
    .B1(_11322_),
    .B2(_11399_),
    .X(_11400_));
 sky130_fd_sc_hd__buf_1 _27329_ (.A(_11400_),
    .X(_11401_));
 sky130_fd_sc_hd__buf_1 _27330_ (.A(_11400_),
    .X(_11402_));
 sky130_fd_sc_hd__o2bb2ai_2 _27331_ (.A1_N(_11397_),
    .A2_N(_11401_),
    .B1(_11397_),
    .B2(_11402_),
    .Y(_11403_));
 sky130_fd_sc_hd__o22a_1 _27332_ (.A1(_11319_),
    .A2(_11320_),
    .B1(_11321_),
    .B2(_11328_),
    .X(_11404_));
 sky130_fd_sc_hd__o2bb2ai_2 _27333_ (.A1_N(_11403_),
    .A2_N(_11404_),
    .B1(_11403_),
    .B2(_11404_),
    .Y(_11405_));
 sky130_fd_sc_hd__buf_1 _27334_ (.A(_11332_),
    .X(_11406_));
 sky130_fd_sc_hd__o32a_1 _27335_ (.A1(_11197_),
    .A2(_11206_),
    .A3(_11325_),
    .B1(_11323_),
    .B2(_11327_),
    .X(_11407_));
 sky130_fd_sc_hd__a2bb2o_1 _27336_ (.A1_N(_11334_),
    .A2_N(_11407_),
    .B1(_11334_),
    .B2(_11407_),
    .X(_11408_));
 sky130_fd_sc_hd__a2bb2o_2 _27337_ (.A1_N(_11406_),
    .A2_N(_11408_),
    .B1(_11406_),
    .B2(_11408_),
    .X(_11409_));
 sky130_fd_sc_hd__o2bb2ai_2 _27338_ (.A1_N(_11405_),
    .A2_N(_11409_),
    .B1(_11405_),
    .B2(_11409_),
    .Y(_11410_));
 sky130_fd_sc_hd__o22a_1 _27339_ (.A1(_11329_),
    .A2(_11330_),
    .B1(_11331_),
    .B2(_11337_),
    .X(_11411_));
 sky130_fd_sc_hd__o2bb2ai_1 _27340_ (.A1_N(_11410_),
    .A2_N(_11411_),
    .B1(_11410_),
    .B2(_11411_),
    .Y(_11412_));
 sky130_fd_sc_hd__o22a_1 _27341_ (.A1(_11343_),
    .A2(_11335_),
    .B1(_11333_),
    .B2(_11336_),
    .X(_11413_));
 sky130_fd_sc_hd__a2bb2o_1 _27342_ (.A1_N(_11342_),
    .A2_N(_11413_),
    .B1(_11342_),
    .B2(_11413_),
    .X(_11414_));
 sky130_fd_sc_hd__a2bb2o_1 _27343_ (.A1_N(_11341_),
    .A2_N(_11414_),
    .B1(_11341_),
    .B2(_11414_),
    .X(_11415_));
 sky130_fd_sc_hd__o2bb2ai_1 _27344_ (.A1_N(_11412_),
    .A2_N(_11415_),
    .B1(_11412_),
    .B2(_11415_),
    .Y(_11416_));
 sky130_fd_sc_hd__o22a_1 _27345_ (.A1(_11338_),
    .A2(_11339_),
    .B1(_11340_),
    .B2(_11346_),
    .X(_11417_));
 sky130_fd_sc_hd__o2bb2a_1 _27346_ (.A1_N(_11416_),
    .A2_N(_11417_),
    .B1(_11416_),
    .B2(_11417_),
    .X(_11418_));
 sky130_vsdinv _27347_ (.A(_11418_),
    .Y(_11419_));
 sky130_fd_sc_hd__o22a_1 _27348_ (.A1(_11353_),
    .A2(_11344_),
    .B1(_11341_),
    .B2(_11345_),
    .X(_11420_));
 sky130_fd_sc_hd__a2bb2o_1 _27349_ (.A1_N(_11352_),
    .A2_N(_11420_),
    .B1(_11235_),
    .B2(_11420_),
    .X(_11421_));
 sky130_fd_sc_hd__a2bb2o_1 _27350_ (.A1_N(_11351_),
    .A2_N(_11421_),
    .B1(_11296_),
    .B2(_11421_),
    .X(_11422_));
 sky130_vsdinv _27351_ (.A(_11422_),
    .Y(_11423_));
 sky130_fd_sc_hd__a22o_1 _27352_ (.A1(_11419_),
    .A2(_11422_),
    .B1(_11418_),
    .B2(_11423_),
    .X(_11424_));
 sky130_fd_sc_hd__o22a_1 _27353_ (.A1(_11347_),
    .A2(_11348_),
    .B1(_11350_),
    .B2(_11357_),
    .X(_11425_));
 sky130_fd_sc_hd__a2bb2o_1 _27354_ (.A1_N(_11424_),
    .A2_N(_11425_),
    .B1(_11424_),
    .B2(_11425_),
    .X(_11426_));
 sky130_fd_sc_hd__clkbuf_1 _27355_ (.A(_11364_),
    .X(_11427_));
 sky130_fd_sc_hd__clkbuf_2 _27356_ (.A(_11296_),
    .X(_11428_));
 sky130_fd_sc_hd__o22a_1 _27357_ (.A1(_11365_),
    .A2(_11355_),
    .B1(_11428_),
    .B2(_11356_),
    .X(_11429_));
 sky130_fd_sc_hd__a2bb2o_1 _27358_ (.A1_N(_11427_),
    .A2_N(_11429_),
    .B1(_11427_),
    .B2(_11429_),
    .X(_11430_));
 sky130_fd_sc_hd__a2bb2o_1 _27359_ (.A1_N(_11368_),
    .A2_N(_11430_),
    .B1(_11368_),
    .B2(_11430_),
    .X(_11431_));
 sky130_fd_sc_hd__a2bb2o_1 _27360_ (.A1_N(_11426_),
    .A2_N(_11431_),
    .B1(_11426_),
    .B2(_11431_),
    .X(_11432_));
 sky130_fd_sc_hd__o22a_1 _27361_ (.A1(_11359_),
    .A2(_11360_),
    .B1(_11361_),
    .B2(_11369_),
    .X(_11433_));
 sky130_fd_sc_hd__a2bb2o_1 _27362_ (.A1_N(_11432_),
    .A2_N(_11433_),
    .B1(_11432_),
    .B2(_11433_),
    .X(_11434_));
 sky130_fd_sc_hd__o22a_1 _27363_ (.A1(_11374_),
    .A2(_11366_),
    .B1(_11362_),
    .B2(_11367_),
    .X(_11435_));
 sky130_fd_sc_hd__or2_1 _27364_ (.A(_11101_),
    .B(_11435_),
    .X(_11436_));
 sky130_fd_sc_hd__a21bo_1 _27365_ (.A1(_11373_),
    .A2(_11435_),
    .B1_N(_11436_),
    .X(_11437_));
 sky130_fd_sc_hd__a2bb2o_1 _27366_ (.A1_N(_11434_),
    .A2_N(_11437_),
    .B1(_11434_),
    .B2(_11437_),
    .X(_11438_));
 sky130_fd_sc_hd__o22a_1 _27367_ (.A1(_11370_),
    .A2(_11371_),
    .B1(_11372_),
    .B2(_11377_),
    .X(_11439_));
 sky130_fd_sc_hd__a2bb2o_1 _27368_ (.A1_N(_11438_),
    .A2_N(_11439_),
    .B1(_11438_),
    .B2(_11439_),
    .X(_11440_));
 sky130_fd_sc_hd__a2bb2o_2 _27369_ (.A1_N(_11376_),
    .A2_N(_11440_),
    .B1(_11376_),
    .B2(_11440_),
    .X(_11441_));
 sky130_fd_sc_hd__o22a_2 _27370_ (.A1(_11378_),
    .A2(_11379_),
    .B1(_11304_),
    .B2(_11380_),
    .X(_11442_));
 sky130_fd_sc_hd__nor2_2 _27371_ (.A(_11441_),
    .B(_11442_),
    .Y(_11443_));
 sky130_fd_sc_hd__a21oi_4 _27372_ (.A1(_11441_),
    .A2(_11442_),
    .B1(_11443_),
    .Y(_11444_));
 sky130_vsdinv _27373_ (.A(_11444_),
    .Y(_11445_));
 sky130_fd_sc_hd__o21ai_1 _27374_ (.A1(_11386_),
    .A2(_11389_),
    .B1(_11383_),
    .Y(_11446_));
 sky130_fd_sc_hd__a2bb2o_1 _27375_ (.A1_N(_11445_),
    .A2_N(_11446_),
    .B1(_11445_),
    .B2(_11446_),
    .X(_02680_));
 sky130_fd_sc_hd__and4_1 _27376_ (.A(_11021_),
    .B(_11050_),
    .C(_11022_),
    .D(_13507_),
    .X(_11447_));
 sky130_fd_sc_hd__o22a_1 _27377_ (.A1(_11720_),
    .A2(_13512_),
    .B1(_11024_),
    .B2(_10751_),
    .X(_11448_));
 sky130_fd_sc_hd__or2_1 _27378_ (.A(_11447_),
    .B(_11448_),
    .X(_11449_));
 sky130_vsdinv _27379_ (.A(_11449_),
    .Y(_11450_));
 sky130_fd_sc_hd__or2_1 _27380_ (.A(_11707_),
    .B(_11258_),
    .X(_11451_));
 sky130_fd_sc_hd__a32o_1 _27381_ (.A1(_11263_),
    .A2(_13071_),
    .A3(_11450_),
    .B1(_11449_),
    .B2(_11451_),
    .X(_11452_));
 sky130_fd_sc_hd__a31o_1 _27382_ (.A1(\pcpi_mul.rs2[30] ),
    .A2(_13508_),
    .A3(_11393_),
    .B1(_11391_),
    .X(_11453_));
 sky130_vsdinv _27383_ (.A(_11453_),
    .Y(_11454_));
 sky130_vsdinv _27384_ (.A(_11452_),
    .Y(_11455_));
 sky130_fd_sc_hd__a22o_1 _27385_ (.A1(_11452_),
    .A2(_11454_),
    .B1(_11455_),
    .B2(_11453_),
    .X(_11456_));
 sky130_fd_sc_hd__a2bb2o_1 _27386_ (.A1_N(_11402_),
    .A2_N(_11456_),
    .B1(_11402_),
    .B2(_11456_),
    .X(_11457_));
 sky130_fd_sc_hd__o22a_1 _27387_ (.A1(_11395_),
    .A2(_11396_),
    .B1(_11397_),
    .B2(_11402_),
    .X(_11458_));
 sky130_fd_sc_hd__o2bb2a_1 _27388_ (.A1_N(_11457_),
    .A2_N(_11458_),
    .B1(_11457_),
    .B2(_11458_),
    .X(_11459_));
 sky130_vsdinv _27389_ (.A(_11459_),
    .Y(_11460_));
 sky130_fd_sc_hd__o22a_1 _27390_ (.A1(_11325_),
    .A2(_11398_),
    .B1(_11322_),
    .B2(_11399_),
    .X(_11461_));
 sky130_fd_sc_hd__a2bb2o_1 _27391_ (.A1_N(_11281_),
    .A2_N(_11461_),
    .B1(_11281_),
    .B2(_11461_),
    .X(_11462_));
 sky130_fd_sc_hd__a2bb2o_1 _27392_ (.A1_N(_11333_),
    .A2_N(_11462_),
    .B1(_11332_),
    .B2(_11462_),
    .X(_11463_));
 sky130_vsdinv _27393_ (.A(_11463_),
    .Y(_11464_));
 sky130_fd_sc_hd__a22o_1 _27394_ (.A1(_11460_),
    .A2(_11463_),
    .B1(_11459_),
    .B2(_11464_),
    .X(_11465_));
 sky130_fd_sc_hd__o22a_1 _27395_ (.A1(_11403_),
    .A2(_11404_),
    .B1(_11405_),
    .B2(_11409_),
    .X(_11466_));
 sky130_fd_sc_hd__o2bb2ai_1 _27396_ (.A1_N(_11465_),
    .A2_N(_11466_),
    .B1(_11465_),
    .B2(_11466_),
    .Y(_11467_));
 sky130_fd_sc_hd__o22a_1 _27397_ (.A1(_11343_),
    .A2(_11407_),
    .B1(_11406_),
    .B2(_11408_),
    .X(_11468_));
 sky130_fd_sc_hd__a2bb2o_1 _27398_ (.A1_N(_11353_),
    .A2_N(_11468_),
    .B1(_11342_),
    .B2(_11468_),
    .X(_11469_));
 sky130_fd_sc_hd__a2bb2o_1 _27399_ (.A1_N(_11354_),
    .A2_N(_11469_),
    .B1(_11354_),
    .B2(_11469_),
    .X(_11470_));
 sky130_fd_sc_hd__o2bb2ai_1 _27400_ (.A1_N(_11467_),
    .A2_N(_11470_),
    .B1(_11467_),
    .B2(_11470_),
    .Y(_11471_));
 sky130_fd_sc_hd__o22a_1 _27401_ (.A1(_11410_),
    .A2(_11411_),
    .B1(_11412_),
    .B2(_11415_),
    .X(_11472_));
 sky130_fd_sc_hd__o2bb2a_1 _27402_ (.A1_N(_11471_),
    .A2_N(_11472_),
    .B1(_11471_),
    .B2(_11472_),
    .X(_11473_));
 sky130_fd_sc_hd__o22a_2 _27403_ (.A1(_11353_),
    .A2(_11413_),
    .B1(_11354_),
    .B2(_11414_),
    .X(_11474_));
 sky130_fd_sc_hd__a2bb2o_1 _27404_ (.A1_N(_11365_),
    .A2_N(_11474_),
    .B1(_11352_),
    .B2(_11474_),
    .X(_11475_));
 sky130_fd_sc_hd__a2bb2oi_2 _27405_ (.A1_N(_11428_),
    .A2_N(_11475_),
    .B1(_11428_),
    .B2(_11475_),
    .Y(_11476_));
 sky130_fd_sc_hd__a2bb2o_1 _27406_ (.A1_N(_11473_),
    .A2_N(_11476_),
    .B1(_11473_),
    .B2(_11476_),
    .X(_11477_));
 sky130_fd_sc_hd__o22a_1 _27407_ (.A1(_11416_),
    .A2(_11417_),
    .B1(_11419_),
    .B2(_11422_),
    .X(_11478_));
 sky130_fd_sc_hd__a2bb2o_1 _27408_ (.A1_N(_11477_),
    .A2_N(_11478_),
    .B1(_11477_),
    .B2(_11478_),
    .X(_11479_));
 sky130_fd_sc_hd__o22a_1 _27409_ (.A1(_11365_),
    .A2(_11420_),
    .B1(_11428_),
    .B2(_11421_),
    .X(_11480_));
 sky130_fd_sc_hd__a2bb2o_1 _27410_ (.A1_N(_11427_),
    .A2_N(_11480_),
    .B1(_11427_),
    .B2(_11480_),
    .X(_11481_));
 sky130_fd_sc_hd__a2bb2o_1 _27411_ (.A1_N(_11368_),
    .A2_N(_11481_),
    .B1(_11362_),
    .B2(_11481_),
    .X(_11482_));
 sky130_fd_sc_hd__a2bb2o_1 _27412_ (.A1_N(_11479_),
    .A2_N(_11482_),
    .B1(_11479_),
    .B2(_11482_),
    .X(_11483_));
 sky130_fd_sc_hd__o22a_1 _27413_ (.A1(_11424_),
    .A2(_11425_),
    .B1(_11426_),
    .B2(_11431_),
    .X(_11484_));
 sky130_fd_sc_hd__a2bb2o_1 _27414_ (.A1_N(_11483_),
    .A2_N(_11484_),
    .B1(_11483_),
    .B2(_11484_),
    .X(_11485_));
 sky130_fd_sc_hd__o22ai_2 _27415_ (.A1(_11374_),
    .A2(_11429_),
    .B1(_11363_),
    .B2(_11430_),
    .Y(_11486_));
 sky130_fd_sc_hd__or2_1 _27416_ (.A(_11101_),
    .B(_11486_),
    .X(_11487_));
 sky130_fd_sc_hd__a21boi_2 _27417_ (.A1(_11373_),
    .A2(_11486_),
    .B1_N(_11487_),
    .Y(_11488_));
 sky130_fd_sc_hd__a2bb2o_1 _27418_ (.A1_N(_11485_),
    .A2_N(_11488_),
    .B1(_11485_),
    .B2(_11488_),
    .X(_11489_));
 sky130_fd_sc_hd__o22a_1 _27419_ (.A1(_11432_),
    .A2(_11433_),
    .B1(_11434_),
    .B2(_11437_),
    .X(_11490_));
 sky130_fd_sc_hd__a2bb2o_1 _27420_ (.A1_N(_11489_),
    .A2_N(_11490_),
    .B1(_11489_),
    .B2(_11490_),
    .X(_11491_));
 sky130_fd_sc_hd__a2bb2o_1 _27421_ (.A1_N(_11436_),
    .A2_N(_11491_),
    .B1(_11436_),
    .B2(_11491_),
    .X(_11492_));
 sky130_fd_sc_hd__o22a_1 _27422_ (.A1(_11438_),
    .A2(_11439_),
    .B1(_11376_),
    .B2(_11440_),
    .X(_11493_));
 sky130_fd_sc_hd__a2bb2o_1 _27423_ (.A1_N(_11492_),
    .A2_N(_11493_),
    .B1(_11492_),
    .B2(_11493_),
    .X(_11494_));
 sky130_fd_sc_hd__o2bb2a_1 _27424_ (.A1_N(_11441_),
    .A2_N(_11442_),
    .B1(_11384_),
    .B2(_11443_),
    .X(_11495_));
 sky130_fd_sc_hd__a31oi_4 _27425_ (.A1(_11385_),
    .A2(_11444_),
    .A3(_11390_),
    .B1(_11495_),
    .Y(_11496_));
 sky130_fd_sc_hd__a2bb2oi_1 _27426_ (.A1_N(_11494_),
    .A2_N(_11496_),
    .B1(_11494_),
    .B2(_11496_),
    .Y(_02681_));
 sky130_fd_sc_hd__o22a_1 _27427_ (.A1(_11492_),
    .A2(_11493_),
    .B1(_11494_),
    .B2(_11496_),
    .X(_11497_));
 sky130_fd_sc_hd__o22a_1 _27428_ (.A1(_11477_),
    .A2(_11478_),
    .B1(_11479_),
    .B2(_11482_),
    .X(_11498_));
 sky130_fd_sc_hd__o22ai_1 _27429_ (.A1(_11465_),
    .A2(_11466_),
    .B1(_11467_),
    .B2(_11470_),
    .Y(_11499_));
 sky130_fd_sc_hd__o2bb2a_1 _27430_ (.A1_N(_11498_),
    .A2_N(_11499_),
    .B1(_11498_),
    .B2(_11499_),
    .X(_11500_));
 sky130_fd_sc_hd__or2b_1 _27431_ (.A(_11068_),
    .B_N(_11468_),
    .X(_11501_));
 sky130_fd_sc_hd__a2bb2o_1 _27432_ (.A1_N(_11067_),
    .A2_N(_11468_),
    .B1(_11063_),
    .B2(_11501_),
    .X(_11502_));
 sky130_fd_sc_hd__a2bb2o_1 _27433_ (.A1_N(_11401_),
    .A2_N(_11502_),
    .B1(_11401_),
    .B2(_11502_),
    .X(_11503_));
 sky130_vsdinv _27434_ (.A(_11503_),
    .Y(_11504_));
 sky130_fd_sc_hd__a32o_1 _27435_ (.A1(_11263_),
    .A2(_13071_),
    .A3(_11503_),
    .B1(_11451_),
    .B2(_11504_),
    .X(_11505_));
 sky130_vsdinv _27436_ (.A(_11505_),
    .Y(_11506_));
 sky130_fd_sc_hd__a22o_1 _27437_ (.A1(_11464_),
    .A2(_11505_),
    .B1(_11463_),
    .B2(_11506_),
    .X(_11507_));
 sky130_fd_sc_hd__o2bb2a_1 _27438_ (.A1_N(_11500_),
    .A2_N(_11507_),
    .B1(_11500_),
    .B2(_11507_),
    .X(_11508_));
 sky130_fd_sc_hd__o22a_1 _27439_ (.A1(_11343_),
    .A2(_11461_),
    .B1(_11406_),
    .B2(_11462_),
    .X(_11509_));
 sky130_fd_sc_hd__or2_1 _27440_ (.A(_11707_),
    .B(_11255_),
    .X(_11510_));
 sky130_fd_sc_hd__o22a_2 _27441_ (.A1(_10281_),
    .A2(_10414_),
    .B1(_10418_),
    .B2(_10417_),
    .X(_11511_));
 sky130_fd_sc_hd__o22a_1 _27442_ (.A1(_11489_),
    .A2(_11490_),
    .B1(_11436_),
    .B2(_11491_),
    .X(_11512_));
 sky130_fd_sc_hd__o2bb2a_1 _27443_ (.A1_N(_11511_),
    .A2_N(_11512_),
    .B1(_11511_),
    .B2(_11512_),
    .X(_11513_));
 sky130_fd_sc_hd__a2bb2o_1 _27444_ (.A1_N(_11510_),
    .A2_N(_11513_),
    .B1(_11510_),
    .B2(_11513_),
    .X(_11514_));
 sky130_fd_sc_hd__o2bb2a_1 _27445_ (.A1_N(_11509_),
    .A2_N(_11514_),
    .B1(_11509_),
    .B2(_11514_),
    .X(_11515_));
 sky130_fd_sc_hd__o2bb2ai_1 _27446_ (.A1_N(_11508_),
    .A2_N(_11515_),
    .B1(_11508_),
    .B2(_11515_),
    .Y(_11516_));
 sky130_fd_sc_hd__a2bb2o_1 _27447_ (.A1_N(_11471_),
    .A2_N(_11472_),
    .B1(_11473_),
    .B2(_11476_),
    .X(_11517_));
 sky130_fd_sc_hd__o22a_1 _27448_ (.A1(_11457_),
    .A2(_11458_),
    .B1(_11460_),
    .B2(_11463_),
    .X(_11518_));
 sky130_fd_sc_hd__a2bb2oi_1 _27449_ (.A1_N(_11517_),
    .A2_N(_11518_),
    .B1(_11517_),
    .B2(_11518_),
    .Y(_11519_));
 sky130_fd_sc_hd__o2bb2a_1 _27450_ (.A1_N(_11516_),
    .A2_N(_11519_),
    .B1(_11516_),
    .B2(_11519_),
    .X(_11520_));
 sky130_fd_sc_hd__a31o_1 _27451_ (.A1(_11263_),
    .A2(_13071_),
    .A3(_11450_),
    .B1(_11447_),
    .X(_11521_));
 sky130_fd_sc_hd__o22ai_2 _27452_ (.A1(_11483_),
    .A2(_11484_),
    .B1(_11485_),
    .B2(_11488_),
    .Y(_11522_));
 sky130_fd_sc_hd__o22a_2 _27453_ (.A1(_11452_),
    .A2(_11454_),
    .B1(_11401_),
    .B2(_11456_),
    .X(_11523_));
 sky130_fd_sc_hd__or2b_1 _27454_ (.A(_10923_),
    .B_N(_11474_),
    .X(_11524_));
 sky130_fd_sc_hd__a2bb2o_2 _27455_ (.A1_N(_10922_),
    .A2_N(_11474_),
    .B1(_10424_),
    .B2(_11524_),
    .X(_11525_));
 sky130_fd_sc_hd__a2bb2oi_2 _27456_ (.A1_N(_11523_),
    .A2_N(_11525_),
    .B1(_11523_),
    .B2(_11525_),
    .Y(_11526_));
 sky130_fd_sc_hd__a2bb2oi_1 _27457_ (.A1_N(_11522_),
    .A2_N(_11526_),
    .B1(_11522_),
    .B2(_11526_),
    .Y(_11527_));
 sky130_fd_sc_hd__o22a_1 _27458_ (.A1(_11374_),
    .A2(_11480_),
    .B1(_11363_),
    .B2(_11481_),
    .X(_11528_));
 sky130_fd_sc_hd__a2bb2o_1 _27459_ (.A1_N(_11487_),
    .A2_N(_11528_),
    .B1(_11487_),
    .B2(_11528_),
    .X(_11529_));
 sky130_fd_sc_hd__nor2_4 _27460_ (.A(_11723_),
    .B(_13508_),
    .Y(_11530_));
 sky130_fd_sc_hd__o2bb2a_1 _27461_ (.A1_N(_11529_),
    .A2_N(_11530_),
    .B1(_11529_),
    .B2(_11530_),
    .X(_11531_));
 sky130_fd_sc_hd__o2bb2a_1 _27462_ (.A1_N(_11527_),
    .A2_N(_11531_),
    .B1(_11527_),
    .B2(_11531_),
    .X(_11532_));
 sky130_fd_sc_hd__a2bb2o_1 _27463_ (.A1_N(_11521_),
    .A2_N(_11532_),
    .B1(_11521_),
    .B2(_11532_),
    .X(_11533_));
 sky130_fd_sc_hd__nand2_1 _27464_ (.A(_11520_),
    .B(_11533_),
    .Y(_11534_));
 sky130_fd_sc_hd__or2_1 _27465_ (.A(_11520_),
    .B(_11533_),
    .X(_11535_));
 sky130_fd_sc_hd__nand2_1 _27466_ (.A(_11534_),
    .B(_11535_),
    .Y(_11536_));
 sky130_fd_sc_hd__nand2_1 _27467_ (.A(_11497_),
    .B(_11536_),
    .Y(_11537_));
 sky130_fd_sc_hd__or2_1 _27468_ (.A(_11497_),
    .B(_11536_),
    .X(_11538_));
 sky130_fd_sc_hd__and2_1 _27469_ (.A(_11537_),
    .B(_11538_),
    .X(_02682_));
 sky130_fd_sc_hd__or2_1 _27470_ (.A(_05392_),
    .B(_05395_),
    .X(_11539_));
 sky130_fd_sc_hd__a2bb2o_1 _27471_ (.A1_N(_05418_),
    .A2_N(_11539_),
    .B1(_05418_),
    .B2(_11539_),
    .X(_02628_));
 sky130_fd_sc_hd__and2_1 _27472_ (.A(_02318_),
    .B(_00066_),
    .X(_00067_));
 sky130_fd_sc_hd__o21a_4 _27473_ (.A1(instr_sra),
    .A2(instr_srai),
    .B1(_13394_),
    .X(_00216_));
 sky130_fd_sc_hd__o21ai_1 _27474_ (.A1(_11784_),
    .A2(_11790_),
    .B1(_00321_),
    .Y(_11540_));
 sky130_vsdinv _27475_ (.A(_11540_),
    .Y(_11541_));
 sky130_fd_sc_hd__o221a_1 _27476_ (.A1(_14161_),
    .A2(_11540_),
    .B1(_11677_),
    .B2(_11541_),
    .C1(_12388_),
    .X(_04072_));
 sky130_fd_sc_hd__conb_1 _27477_ (.LO(net134));
 sky130_fd_sc_hd__conb_1 _27478_ (.LO(net145));
 sky130_fd_sc_hd__conb_1 _27479_ (.LO(net167));
 sky130_fd_sc_hd__conb_1 _27480_ (.LO(net178));
 sky130_fd_sc_hd__conb_1 _27481_ (.LO(net371));
 sky130_fd_sc_hd__conb_1 _27482_ (.LO(net382));
 sky130_fd_sc_hd__conb_1 _27483_ (.LO(net393));
 sky130_fd_sc_hd__conb_1 _27484_ (.LO(net400));
 sky130_fd_sc_hd__conb_1 _27485_ (.LO(net401));
 sky130_fd_sc_hd__conb_1 _27486_ (.LO(net402));
 sky130_fd_sc_hd__conb_1 _27487_ (.LO(net403));
 sky130_fd_sc_hd__conb_1 _27488_ (.LO(net404));
 sky130_fd_sc_hd__conb_1 _27489_ (.LO(net405));
 sky130_fd_sc_hd__conb_1 _27490_ (.LO(net406));
 sky130_fd_sc_hd__conb_1 _27491_ (.LO(net372));
 sky130_fd_sc_hd__conb_1 _27492_ (.LO(net373));
 sky130_fd_sc_hd__conb_1 _27493_ (.LO(net374));
 sky130_fd_sc_hd__conb_1 _27494_ (.LO(net375));
 sky130_fd_sc_hd__conb_1 _27495_ (.LO(net376));
 sky130_fd_sc_hd__conb_1 _27496_ (.LO(net377));
 sky130_fd_sc_hd__conb_1 _27497_ (.LO(net378));
 sky130_fd_sc_hd__conb_1 _27498_ (.LO(net379));
 sky130_fd_sc_hd__conb_1 _27499_ (.LO(net380));
 sky130_fd_sc_hd__conb_1 _27500_ (.LO(net381));
 sky130_fd_sc_hd__conb_1 _27501_ (.LO(net383));
 sky130_fd_sc_hd__conb_1 _27502_ (.LO(net384));
 sky130_fd_sc_hd__conb_1 _27503_ (.LO(net385));
 sky130_fd_sc_hd__conb_1 _27504_ (.LO(net386));
 sky130_fd_sc_hd__conb_1 _27505_ (.LO(net387));
 sky130_fd_sc_hd__conb_1 _27506_ (.LO(net388));
 sky130_fd_sc_hd__conb_1 _27507_ (.LO(net389));
 sky130_fd_sc_hd__conb_1 _27508_ (.LO(net390));
 sky130_fd_sc_hd__conb_1 _27509_ (.LO(net391));
 sky130_fd_sc_hd__conb_1 _27510_ (.LO(net392));
 sky130_fd_sc_hd__conb_1 _27511_ (.LO(net394));
 sky130_fd_sc_hd__conb_1 _27512_ (.LO(net395));
 sky130_fd_sc_hd__conb_1 _27513_ (.LO(net396));
 sky130_fd_sc_hd__conb_1 _27514_ (.LO(net397));
 sky130_fd_sc_hd__conb_1 _27515_ (.LO(net398));
 sky130_fd_sc_hd__conb_1 _27516_ (.LO(net399));
 sky130_fd_sc_hd__conb_1 _27517_ (.LO(net407));
 sky130_fd_sc_hd__conb_1 _27518_ (.LO(_00313_));
 sky130_fd_sc_hd__buf_2 _27519_ (.A(net200),
    .X(net338));
 sky130_fd_sc_hd__clkbuf_1 _27520_ (.A(net211),
    .X(net349));
 sky130_fd_sc_hd__buf_4 _27521_ (.A(net460),
    .X(net360));
 sky130_fd_sc_hd__clkbuf_2 _27522_ (.A(net225),
    .X(net363));
 sky130_fd_sc_hd__clkbuf_4 _27523_ (.A(net458),
    .X(net364));
 sky130_fd_sc_hd__buf_2 _27524_ (.A(net227),
    .X(net365));
 sky130_fd_sc_hd__clkbuf_1 _27525_ (.A(net228),
    .X(net366));
 sky130_fd_sc_hd__clkbuf_4 _27526_ (.A(net229),
    .X(net367));
 sky130_fd_sc_hd__mux2_8 _27527_ (.A0(decoder_trigger),
    .A1(_02410_),
    .S(_00309_),
    .X(_14285_));
 sky130_fd_sc_hd__mux2_2 _27528_ (.A0(\reg_out[2] ),
    .A1(\reg_next_pc[2] ),
    .S(_02183_),
    .X(_02184_));
 sky130_fd_sc_hd__mux2_8 _27529_ (.A0(_02184_),
    .A1(net328),
    .S(net416),
    .X(net189));
 sky130_fd_sc_hd__mux2_2 _27530_ (.A0(\reg_out[3] ),
    .A1(\reg_next_pc[3] ),
    .S(_02183_),
    .X(_02185_));
 sky130_fd_sc_hd__mux2_8 _27531_ (.A0(_02185_),
    .A1(net331),
    .S(net416),
    .X(net192));
 sky130_fd_sc_hd__mux2_1 _27532_ (.A0(\reg_out[4] ),
    .A1(\reg_next_pc[4] ),
    .S(_02183_),
    .X(_02186_));
 sky130_fd_sc_hd__mux2_8 _27533_ (.A0(_02186_),
    .A1(net332),
    .S(net419),
    .X(net193));
 sky130_fd_sc_hd__mux2_1 _27534_ (.A0(\reg_out[5] ),
    .A1(\reg_next_pc[5] ),
    .S(_02183_),
    .X(_02187_));
 sky130_fd_sc_hd__mux2_8 _27535_ (.A0(_02187_),
    .A1(net333),
    .S(net416),
    .X(net194));
 sky130_fd_sc_hd__mux2_2 _27536_ (.A0(\reg_out[6] ),
    .A1(\reg_next_pc[6] ),
    .S(_02183_),
    .X(_02188_));
 sky130_fd_sc_hd__mux2_8 _27537_ (.A0(_02188_),
    .A1(net334),
    .S(net416),
    .X(net195));
 sky130_fd_sc_hd__mux2_2 _27538_ (.A0(\reg_out[7] ),
    .A1(\reg_next_pc[7] ),
    .S(_02183_),
    .X(_02189_));
 sky130_fd_sc_hd__mux2_8 _27539_ (.A0(_02189_),
    .A1(net335),
    .S(net416),
    .X(net196));
 sky130_fd_sc_hd__mux2_2 _27540_ (.A0(\reg_out[8] ),
    .A1(\reg_next_pc[8] ),
    .S(_02183_),
    .X(_02190_));
 sky130_fd_sc_hd__mux2_4 _27541_ (.A0(_02190_),
    .A1(net336),
    .S(net417),
    .X(net197));
 sky130_fd_sc_hd__mux2_1 _27542_ (.A0(\reg_out[9] ),
    .A1(\reg_next_pc[9] ),
    .S(_02183_),
    .X(_02191_));
 sky130_fd_sc_hd__mux2_8 _27543_ (.A0(_02191_),
    .A1(net337),
    .S(net419),
    .X(net198));
 sky130_fd_sc_hd__mux2_1 _27544_ (.A0(\reg_out[10] ),
    .A1(\reg_next_pc[10] ),
    .S(_02183_),
    .X(_02192_));
 sky130_fd_sc_hd__mux2_8 _27545_ (.A0(_02192_),
    .A1(net307),
    .S(net419),
    .X(net168));
 sky130_fd_sc_hd__mux2_1 _27546_ (.A0(\reg_out[11] ),
    .A1(\reg_next_pc[11] ),
    .S(_02183_),
    .X(_02193_));
 sky130_fd_sc_hd__mux2_8 _27547_ (.A0(_02193_),
    .A1(net308),
    .S(net419),
    .X(net169));
 sky130_fd_sc_hd__mux2_1 _27548_ (.A0(\reg_out[12] ),
    .A1(\reg_next_pc[12] ),
    .S(_02183_),
    .X(_02194_));
 sky130_fd_sc_hd__mux2_4 _27549_ (.A0(_02194_),
    .A1(net309),
    .S(net416),
    .X(net170));
 sky130_fd_sc_hd__mux2_2 _27550_ (.A0(\reg_out[13] ),
    .A1(\reg_next_pc[13] ),
    .S(_02183_),
    .X(_02195_));
 sky130_fd_sc_hd__mux2_8 _27551_ (.A0(_02195_),
    .A1(net310),
    .S(net416),
    .X(net171));
 sky130_fd_sc_hd__mux2_1 _27552_ (.A0(\reg_out[14] ),
    .A1(\reg_next_pc[14] ),
    .S(_02183_),
    .X(_02196_));
 sky130_fd_sc_hd__mux2_8 _27553_ (.A0(_02196_),
    .A1(net311),
    .S(net418),
    .X(net172));
 sky130_fd_sc_hd__mux2_2 _27554_ (.A0(\reg_out[15] ),
    .A1(\reg_next_pc[15] ),
    .S(_02183_),
    .X(_02197_));
 sky130_fd_sc_hd__mux2_2 _27555_ (.A0(_02197_),
    .A1(net312),
    .S(net417),
    .X(net173));
 sky130_fd_sc_hd__mux2_1 _27556_ (.A0(\reg_out[16] ),
    .A1(\reg_next_pc[16] ),
    .S(_02183_),
    .X(_02198_));
 sky130_fd_sc_hd__mux2_8 _27557_ (.A0(_02198_),
    .A1(net313),
    .S(net417),
    .X(net174));
 sky130_fd_sc_hd__mux2_1 _27558_ (.A0(\reg_out[17] ),
    .A1(\reg_next_pc[17] ),
    .S(_02183_),
    .X(_02199_));
 sky130_fd_sc_hd__mux2_8 _27559_ (.A0(_02199_),
    .A1(net314),
    .S(net418),
    .X(net175));
 sky130_fd_sc_hd__mux2_1 _27560_ (.A0(\reg_out[18] ),
    .A1(\reg_next_pc[18] ),
    .S(_02183_),
    .X(_02200_));
 sky130_fd_sc_hd__mux2_4 _27561_ (.A0(_02200_),
    .A1(net315),
    .S(net417),
    .X(net176));
 sky130_fd_sc_hd__mux2_1 _27562_ (.A0(\reg_out[19] ),
    .A1(\reg_next_pc[19] ),
    .S(_02183_),
    .X(_02201_));
 sky130_fd_sc_hd__mux2_8 _27563_ (.A0(_02201_),
    .A1(net316),
    .S(net417),
    .X(net177));
 sky130_fd_sc_hd__mux2_1 _27564_ (.A0(\reg_out[20] ),
    .A1(\reg_next_pc[20] ),
    .S(_02183_),
    .X(_02202_));
 sky130_fd_sc_hd__mux2_4 _27565_ (.A0(_02202_),
    .A1(net318),
    .S(net417),
    .X(net179));
 sky130_fd_sc_hd__mux2_1 _27566_ (.A0(\reg_out[21] ),
    .A1(\reg_next_pc[21] ),
    .S(_02183_),
    .X(_02203_));
 sky130_fd_sc_hd__mux2_8 _27567_ (.A0(_02203_),
    .A1(net319),
    .S(net418),
    .X(net180));
 sky130_fd_sc_hd__mux2_1 _27568_ (.A0(\reg_out[22] ),
    .A1(\reg_next_pc[22] ),
    .S(_02183_),
    .X(_02204_));
 sky130_fd_sc_hd__mux2_8 _27569_ (.A0(_02204_),
    .A1(net320),
    .S(net417),
    .X(net181));
 sky130_fd_sc_hd__mux2_2 _27570_ (.A0(\reg_out[23] ),
    .A1(\reg_next_pc[23] ),
    .S(_02183_),
    .X(_02205_));
 sky130_fd_sc_hd__mux2_4 _27571_ (.A0(_02205_),
    .A1(net321),
    .S(net417),
    .X(net182));
 sky130_fd_sc_hd__mux2_2 _27572_ (.A0(\reg_out[24] ),
    .A1(\reg_next_pc[24] ),
    .S(_02183_),
    .X(_02206_));
 sky130_fd_sc_hd__mux2_8 _27573_ (.A0(_02206_),
    .A1(net322),
    .S(net417),
    .X(net183));
 sky130_fd_sc_hd__mux2_2 _27574_ (.A0(\reg_out[25] ),
    .A1(\reg_next_pc[25] ),
    .S(_02183_),
    .X(_02207_));
 sky130_fd_sc_hd__mux2_4 _27575_ (.A0(_02207_),
    .A1(net323),
    .S(net417),
    .X(net184));
 sky130_fd_sc_hd__mux2_1 _27576_ (.A0(\reg_out[26] ),
    .A1(\reg_next_pc[26] ),
    .S(_02183_),
    .X(_02208_));
 sky130_fd_sc_hd__mux2_4 _27577_ (.A0(_02208_),
    .A1(net324),
    .S(net418),
    .X(net185));
 sky130_fd_sc_hd__mux2_1 _27578_ (.A0(\reg_out[27] ),
    .A1(\reg_next_pc[27] ),
    .S(_02183_),
    .X(_02209_));
 sky130_fd_sc_hd__mux2_4 _27579_ (.A0(_02209_),
    .A1(net325),
    .S(net418),
    .X(net186));
 sky130_fd_sc_hd__mux2_2 _27580_ (.A0(\reg_out[28] ),
    .A1(\reg_next_pc[28] ),
    .S(_02183_),
    .X(_02210_));
 sky130_fd_sc_hd__mux2_8 _27581_ (.A0(_02210_),
    .A1(net326),
    .S(net418),
    .X(net187));
 sky130_fd_sc_hd__mux2_1 _27582_ (.A0(\reg_out[29] ),
    .A1(\reg_next_pc[29] ),
    .S(_02183_),
    .X(_02211_));
 sky130_fd_sc_hd__mux2_8 _27583_ (.A0(_02211_),
    .A1(net327),
    .S(net419),
    .X(net188));
 sky130_fd_sc_hd__mux2_1 _27584_ (.A0(\reg_out[30] ),
    .A1(\reg_next_pc[30] ),
    .S(_02183_),
    .X(_02212_));
 sky130_fd_sc_hd__mux2_8 _27585_ (.A0(_02212_),
    .A1(net329),
    .S(net419),
    .X(net190));
 sky130_fd_sc_hd__mux2_2 _27586_ (.A0(\reg_out[31] ),
    .A1(\reg_next_pc[31] ),
    .S(_02183_),
    .X(_02213_));
 sky130_fd_sc_hd__mux2_4 _27587_ (.A0(_02213_),
    .A1(net330),
    .S(net416),
    .X(net191));
 sky130_fd_sc_hd__mux2_4 _27588_ (.A0(_02167_),
    .A1(net368),
    .S(_01683_),
    .X(net230));
 sky130_fd_sc_hd__mux2_8 _27589_ (.A0(_02168_),
    .A1(net369),
    .S(net421),
    .X(net231));
 sky130_fd_sc_hd__mux2_8 _27590_ (.A0(_02169_),
    .A1(net339),
    .S(net421),
    .X(net201));
 sky130_fd_sc_hd__mux2_4 _27591_ (.A0(_02170_),
    .A1(net340),
    .S(net421),
    .X(net202));
 sky130_fd_sc_hd__mux2_4 _27592_ (.A0(_02171_),
    .A1(net341),
    .S(_01683_),
    .X(net203));
 sky130_fd_sc_hd__mux2_4 _27593_ (.A0(_02172_),
    .A1(net342),
    .S(_01683_),
    .X(net204));
 sky130_fd_sc_hd__mux2_8 _27594_ (.A0(_02173_),
    .A1(net343),
    .S(net420),
    .X(net205));
 sky130_fd_sc_hd__mux2_4 _27595_ (.A0(_02174_),
    .A1(net344),
    .S(_01683_),
    .X(net206));
 sky130_fd_sc_hd__mux2_8 _27596_ (.A0(_02175_),
    .A1(net345),
    .S(net421),
    .X(net207));
 sky130_fd_sc_hd__mux2_4 _27597_ (.A0(_02176_),
    .A1(net346),
    .S(net420),
    .X(net208));
 sky130_fd_sc_hd__mux2_8 _27598_ (.A0(_02177_),
    .A1(net347),
    .S(net420),
    .X(net209));
 sky130_fd_sc_hd__mux2_4 _27599_ (.A0(_02178_),
    .A1(net348),
    .S(net420),
    .X(net210));
 sky130_fd_sc_hd__mux2_8 _27600_ (.A0(_02179_),
    .A1(net350),
    .S(net420),
    .X(net212));
 sky130_fd_sc_hd__mux2_4 _27601_ (.A0(_02180_),
    .A1(net351),
    .S(net420),
    .X(net213));
 sky130_fd_sc_hd__mux2_8 _27602_ (.A0(_02181_),
    .A1(net352),
    .S(net420),
    .X(net214));
 sky130_fd_sc_hd__mux2_8 _27603_ (.A0(_02182_),
    .A1(net353),
    .S(net420),
    .X(net215));
 sky130_fd_sc_hd__mux2_4 _27604_ (.A0(_02167_),
    .A1(net354),
    .S(_01683_),
    .X(net216));
 sky130_fd_sc_hd__mux2_8 _27605_ (.A0(_02168_),
    .A1(net355),
    .S(net421),
    .X(net217));
 sky130_fd_sc_hd__mux2_8 _27606_ (.A0(_02169_),
    .A1(net356),
    .S(net421),
    .X(net218));
 sky130_fd_sc_hd__mux2_8 _27607_ (.A0(_02170_),
    .A1(net357),
    .S(_01683_),
    .X(net219));
 sky130_fd_sc_hd__mux2_8 _27608_ (.A0(_02171_),
    .A1(net358),
    .S(_01683_),
    .X(net220));
 sky130_fd_sc_hd__mux2_8 _27609_ (.A0(_02172_),
    .A1(net359),
    .S(_01683_),
    .X(net221));
 sky130_fd_sc_hd__mux2_8 _27610_ (.A0(_02173_),
    .A1(net361),
    .S(net420),
    .X(net223));
 sky130_fd_sc_hd__mux2_4 _27611_ (.A0(_02174_),
    .A1(net362),
    .S(_01683_),
    .X(net224));
 sky130_fd_sc_hd__mux2_1 _27612_ (.A0(\mem_rdata_q[7] ),
    .A1(net62),
    .S(mem_xfer),
    .X(\mem_rdata_latched[7] ));
 sky130_fd_sc_hd__mux2_1 _27613_ (.A0(\mem_rdata_q[8] ),
    .A1(net63),
    .S(mem_xfer),
    .X(\mem_rdata_latched[8] ));
 sky130_fd_sc_hd__mux2_1 _27614_ (.A0(\mem_rdata_q[9] ),
    .A1(net64),
    .S(mem_xfer),
    .X(\mem_rdata_latched[9] ));
 sky130_fd_sc_hd__mux2_1 _27615_ (.A0(\mem_rdata_q[10] ),
    .A1(net34),
    .S(mem_xfer),
    .X(\mem_rdata_latched[10] ));
 sky130_fd_sc_hd__mux2_1 _27616_ (.A0(\mem_rdata_q[11] ),
    .A1(net35),
    .S(net415),
    .X(\mem_rdata_latched[11] ));
 sky130_fd_sc_hd__mux2_2 _27617_ (.A0(\mem_rdata_q[12] ),
    .A1(net36),
    .S(mem_xfer),
    .X(\mem_rdata_latched[12] ));
 sky130_fd_sc_hd__mux2_2 _27618_ (.A0(\mem_rdata_q[13] ),
    .A1(net37),
    .S(mem_xfer),
    .X(\mem_rdata_latched[13] ));
 sky130_fd_sc_hd__mux2_2 _27619_ (.A0(\mem_rdata_q[14] ),
    .A1(net38),
    .S(mem_xfer),
    .X(\mem_rdata_latched[14] ));
 sky130_fd_sc_hd__mux2_2 _27620_ (.A0(\mem_rdata_q[15] ),
    .A1(net39),
    .S(mem_xfer),
    .X(\mem_rdata_latched[15] ));
 sky130_fd_sc_hd__mux2_1 _27621_ (.A0(\mem_rdata_q[16] ),
    .A1(net40),
    .S(net415),
    .X(\mem_rdata_latched[16] ));
 sky130_fd_sc_hd__mux2_1 _27622_ (.A0(\mem_rdata_q[17] ),
    .A1(net41),
    .S(net415),
    .X(\mem_rdata_latched[17] ));
 sky130_fd_sc_hd__mux2_1 _27623_ (.A0(\mem_rdata_q[18] ),
    .A1(net42),
    .S(net415),
    .X(\mem_rdata_latched[18] ));
 sky130_fd_sc_hd__mux2_1 _27624_ (.A0(\mem_rdata_q[19] ),
    .A1(net43),
    .S(net415),
    .X(\mem_rdata_latched[19] ));
 sky130_fd_sc_hd__mux2_1 _27625_ (.A0(\mem_rdata_q[20] ),
    .A1(net464),
    .S(net415),
    .X(\mem_rdata_latched[20] ));
 sky130_fd_sc_hd__mux2_1 _27626_ (.A0(\mem_rdata_q[21] ),
    .A1(net46),
    .S(mem_xfer),
    .X(\mem_rdata_latched[21] ));
 sky130_fd_sc_hd__mux2_1 _27627_ (.A0(\mem_rdata_q[22] ),
    .A1(net47),
    .S(mem_xfer),
    .X(\mem_rdata_latched[22] ));
 sky130_fd_sc_hd__mux2_1 _27628_ (.A0(\mem_rdata_q[23] ),
    .A1(net48),
    .S(net415),
    .X(\mem_rdata_latched[23] ));
 sky130_fd_sc_hd__mux2_1 _27629_ (.A0(\mem_rdata_q[24] ),
    .A1(net49),
    .S(net415),
    .X(\mem_rdata_latched[24] ));
 sky130_fd_sc_hd__mux2_1 _27630_ (.A0(\mem_rdata_q[25] ),
    .A1(net50),
    .S(net415),
    .X(\mem_rdata_latched[25] ));
 sky130_fd_sc_hd__mux2_1 _27631_ (.A0(\mem_rdata_q[26] ),
    .A1(net51),
    .S(mem_xfer),
    .X(\mem_rdata_latched[26] ));
 sky130_fd_sc_hd__mux2_2 _27632_ (.A0(\mem_rdata_q[27] ),
    .A1(net52),
    .S(net415),
    .X(\mem_rdata_latched[27] ));
 sky130_fd_sc_hd__mux2_2 _27633_ (.A0(\mem_rdata_q[28] ),
    .A1(net53),
    .S(net415),
    .X(\mem_rdata_latched[28] ));
 sky130_fd_sc_hd__mux2_1 _27634_ (.A0(\mem_rdata_q[29] ),
    .A1(net54),
    .S(net415),
    .X(\mem_rdata_latched[29] ));
 sky130_fd_sc_hd__mux2_1 _27635_ (.A0(\mem_rdata_q[30] ),
    .A1(net56),
    .S(net415),
    .X(\mem_rdata_latched[30] ));
 sky130_fd_sc_hd__mux2_1 _27636_ (.A0(\mem_rdata_q[31] ),
    .A1(net57),
    .S(net415),
    .X(\mem_rdata_latched[31] ));
 sky130_fd_sc_hd__mux2_1 _27637_ (.A0(_02134_),
    .A1(\alu_add_sub[0] ),
    .S(_02133_),
    .X(\alu_out[0] ));
 sky130_fd_sc_hd__mux2_1 _27638_ (.A0(_02135_),
    .A1(\alu_add_sub[1] ),
    .S(_02133_),
    .X(\alu_out[1] ));
 sky130_fd_sc_hd__mux2_1 _27639_ (.A0(_02136_),
    .A1(\alu_add_sub[2] ),
    .S(_02133_),
    .X(\alu_out[2] ));
 sky130_fd_sc_hd__mux2_1 _27640_ (.A0(_02137_),
    .A1(\alu_add_sub[3] ),
    .S(_02133_),
    .X(\alu_out[3] ));
 sky130_fd_sc_hd__mux2_1 _27641_ (.A0(_02138_),
    .A1(\alu_add_sub[4] ),
    .S(_02133_),
    .X(\alu_out[4] ));
 sky130_fd_sc_hd__mux2_1 _27642_ (.A0(_02139_),
    .A1(\alu_add_sub[5] ),
    .S(_02133_),
    .X(\alu_out[5] ));
 sky130_fd_sc_hd__mux2_1 _27643_ (.A0(_02140_),
    .A1(\alu_add_sub[6] ),
    .S(_02133_),
    .X(\alu_out[6] ));
 sky130_fd_sc_hd__mux2_1 _27644_ (.A0(_02141_),
    .A1(\alu_add_sub[7] ),
    .S(_02133_),
    .X(\alu_out[7] ));
 sky130_fd_sc_hd__mux2_1 _27645_ (.A0(_02142_),
    .A1(\alu_add_sub[8] ),
    .S(_02133_),
    .X(\alu_out[8] ));
 sky130_fd_sc_hd__mux2_1 _27646_ (.A0(_02143_),
    .A1(\alu_add_sub[9] ),
    .S(_02133_),
    .X(\alu_out[9] ));
 sky130_fd_sc_hd__mux2_1 _27647_ (.A0(_02144_),
    .A1(\alu_add_sub[10] ),
    .S(_02133_),
    .X(\alu_out[10] ));
 sky130_fd_sc_hd__mux2_1 _27648_ (.A0(_02145_),
    .A1(\alu_add_sub[11] ),
    .S(_02133_),
    .X(\alu_out[11] ));
 sky130_fd_sc_hd__mux2_1 _27649_ (.A0(_02146_),
    .A1(\alu_add_sub[12] ),
    .S(_02133_),
    .X(\alu_out[12] ));
 sky130_fd_sc_hd__mux2_1 _27650_ (.A0(_02147_),
    .A1(\alu_add_sub[13] ),
    .S(_02133_),
    .X(\alu_out[13] ));
 sky130_fd_sc_hd__mux2_1 _27651_ (.A0(_02148_),
    .A1(\alu_add_sub[14] ),
    .S(_02133_),
    .X(\alu_out[14] ));
 sky130_fd_sc_hd__mux2_1 _27652_ (.A0(_02149_),
    .A1(\alu_add_sub[15] ),
    .S(_02133_),
    .X(\alu_out[15] ));
 sky130_fd_sc_hd__mux2_1 _27653_ (.A0(_02150_),
    .A1(\alu_add_sub[16] ),
    .S(_02133_),
    .X(\alu_out[16] ));
 sky130_fd_sc_hd__mux2_1 _27654_ (.A0(_02151_),
    .A1(\alu_add_sub[17] ),
    .S(_02133_),
    .X(\alu_out[17] ));
 sky130_fd_sc_hd__mux2_1 _27655_ (.A0(_02152_),
    .A1(\alu_add_sub[18] ),
    .S(_02133_),
    .X(\alu_out[18] ));
 sky130_fd_sc_hd__mux2_1 _27656_ (.A0(_02153_),
    .A1(\alu_add_sub[19] ),
    .S(_02133_),
    .X(\alu_out[19] ));
 sky130_fd_sc_hd__mux2_1 _27657_ (.A0(_02154_),
    .A1(\alu_add_sub[20] ),
    .S(_02133_),
    .X(\alu_out[20] ));
 sky130_fd_sc_hd__mux2_1 _27658_ (.A0(_02155_),
    .A1(\alu_add_sub[21] ),
    .S(_02133_),
    .X(\alu_out[21] ));
 sky130_fd_sc_hd__mux2_1 _27659_ (.A0(_02156_),
    .A1(\alu_add_sub[22] ),
    .S(_02133_),
    .X(\alu_out[22] ));
 sky130_fd_sc_hd__mux2_1 _27660_ (.A0(_02157_),
    .A1(\alu_add_sub[23] ),
    .S(_02133_),
    .X(\alu_out[23] ));
 sky130_fd_sc_hd__mux2_1 _27661_ (.A0(_02158_),
    .A1(\alu_add_sub[24] ),
    .S(_02133_),
    .X(\alu_out[24] ));
 sky130_fd_sc_hd__mux2_1 _27662_ (.A0(_02159_),
    .A1(\alu_add_sub[25] ),
    .S(_02133_),
    .X(\alu_out[25] ));
 sky130_fd_sc_hd__mux2_1 _27663_ (.A0(_02160_),
    .A1(\alu_add_sub[26] ),
    .S(_02133_),
    .X(\alu_out[26] ));
 sky130_fd_sc_hd__mux2_1 _27664_ (.A0(_02161_),
    .A1(\alu_add_sub[27] ),
    .S(_02133_),
    .X(\alu_out[27] ));
 sky130_fd_sc_hd__mux2_1 _27665_ (.A0(_02162_),
    .A1(\alu_add_sub[28] ),
    .S(_02133_),
    .X(\alu_out[28] ));
 sky130_fd_sc_hd__mux2_1 _27666_ (.A0(_02163_),
    .A1(\alu_add_sub[29] ),
    .S(_02133_),
    .X(\alu_out[29] ));
 sky130_fd_sc_hd__mux2_1 _27667_ (.A0(_02164_),
    .A1(\alu_add_sub[30] ),
    .S(_02133_),
    .X(\alu_out[30] ));
 sky130_fd_sc_hd__mux2_1 _27668_ (.A0(_02165_),
    .A1(\alu_add_sub[31] ),
    .S(_02133_),
    .X(\alu_out[31] ));
 sky130_fd_sc_hd__mux2_8 _27669_ (.A0(_02071_),
    .A1(\reg_next_pc[0] ),
    .S(_02069_),
    .X(\cpuregs_wrdata[0] ));
 sky130_fd_sc_hd__mux2_8 _27670_ (.A0(_02072_),
    .A1(\reg_pc[1] ),
    .S(net414),
    .X(\cpuregs_wrdata[1] ));
 sky130_fd_sc_hd__mux2_8 _27671_ (.A0(_02074_),
    .A1(_02073_),
    .S(net414),
    .X(\cpuregs_wrdata[2] ));
 sky130_fd_sc_hd__mux2_8 _27672_ (.A0(_02076_),
    .A1(_02075_),
    .S(net414),
    .X(\cpuregs_wrdata[3] ));
 sky130_fd_sc_hd__mux2_8 _27673_ (.A0(_02078_),
    .A1(_02077_),
    .S(net414),
    .X(\cpuregs_wrdata[4] ));
 sky130_fd_sc_hd__mux2_4 _27674_ (.A0(_02080_),
    .A1(_02079_),
    .S(net414),
    .X(\cpuregs_wrdata[5] ));
 sky130_fd_sc_hd__mux2_4 _27675_ (.A0(_02082_),
    .A1(_02081_),
    .S(net414),
    .X(\cpuregs_wrdata[6] ));
 sky130_fd_sc_hd__mux2_4 _27676_ (.A0(_02084_),
    .A1(_02083_),
    .S(net414),
    .X(\cpuregs_wrdata[7] ));
 sky130_fd_sc_hd__mux2_8 _27677_ (.A0(_02086_),
    .A1(_02085_),
    .S(net414),
    .X(\cpuregs_wrdata[8] ));
 sky130_fd_sc_hd__mux2_8 _27678_ (.A0(_02088_),
    .A1(_02087_),
    .S(net414),
    .X(\cpuregs_wrdata[9] ));
 sky130_fd_sc_hd__mux2_8 _27679_ (.A0(_02090_),
    .A1(_02089_),
    .S(net414),
    .X(\cpuregs_wrdata[10] ));
 sky130_fd_sc_hd__mux2_8 _27680_ (.A0(_02092_),
    .A1(_02091_),
    .S(net414),
    .X(\cpuregs_wrdata[11] ));
 sky130_fd_sc_hd__mux2_4 _27681_ (.A0(_02094_),
    .A1(_02093_),
    .S(net414),
    .X(\cpuregs_wrdata[12] ));
 sky130_fd_sc_hd__mux2_4 _27682_ (.A0(_02096_),
    .A1(_02095_),
    .S(net414),
    .X(\cpuregs_wrdata[13] ));
 sky130_fd_sc_hd__mux2_4 _27683_ (.A0(_02098_),
    .A1(_02097_),
    .S(net414),
    .X(\cpuregs_wrdata[14] ));
 sky130_fd_sc_hd__mux2_4 _27684_ (.A0(_02100_),
    .A1(_02099_),
    .S(net414),
    .X(\cpuregs_wrdata[15] ));
 sky130_fd_sc_hd__mux2_4 _27685_ (.A0(_02102_),
    .A1(_02101_),
    .S(net414),
    .X(\cpuregs_wrdata[16] ));
 sky130_fd_sc_hd__mux2_4 _27686_ (.A0(_02104_),
    .A1(_02103_),
    .S(net414),
    .X(\cpuregs_wrdata[17] ));
 sky130_fd_sc_hd__mux2_4 _27687_ (.A0(_02106_),
    .A1(_02105_),
    .S(net414),
    .X(\cpuregs_wrdata[18] ));
 sky130_fd_sc_hd__mux2_4 _27688_ (.A0(_02108_),
    .A1(_02107_),
    .S(net414),
    .X(\cpuregs_wrdata[19] ));
 sky130_fd_sc_hd__mux2_2 _27689_ (.A0(_02110_),
    .A1(_02109_),
    .S(net414),
    .X(\cpuregs_wrdata[20] ));
 sky130_fd_sc_hd__mux2_2 _27690_ (.A0(_02112_),
    .A1(_02111_),
    .S(net414),
    .X(\cpuregs_wrdata[21] ));
 sky130_fd_sc_hd__mux2_2 _27691_ (.A0(_02114_),
    .A1(_02113_),
    .S(net414),
    .X(\cpuregs_wrdata[22] ));
 sky130_fd_sc_hd__mux2_2 _27692_ (.A0(_02116_),
    .A1(_02115_),
    .S(net414),
    .X(\cpuregs_wrdata[23] ));
 sky130_fd_sc_hd__mux2_4 _27693_ (.A0(_02118_),
    .A1(_02117_),
    .S(net414),
    .X(\cpuregs_wrdata[24] ));
 sky130_fd_sc_hd__mux2_4 _27694_ (.A0(_02120_),
    .A1(_02119_),
    .S(net414),
    .X(\cpuregs_wrdata[25] ));
 sky130_fd_sc_hd__mux2_4 _27695_ (.A0(_02122_),
    .A1(_02121_),
    .S(net414),
    .X(\cpuregs_wrdata[26] ));
 sky130_fd_sc_hd__mux2_4 _27696_ (.A0(_02124_),
    .A1(_02123_),
    .S(_02069_),
    .X(\cpuregs_wrdata[27] ));
 sky130_fd_sc_hd__mux2_2 _27697_ (.A0(_02126_),
    .A1(_02125_),
    .S(_02069_),
    .X(\cpuregs_wrdata[28] ));
 sky130_fd_sc_hd__mux2_4 _27698_ (.A0(_02128_),
    .A1(_02127_),
    .S(_02069_),
    .X(\cpuregs_wrdata[29] ));
 sky130_fd_sc_hd__mux2_4 _27699_ (.A0(_02130_),
    .A1(_02129_),
    .S(_02069_),
    .X(\cpuregs_wrdata[30] ));
 sky130_fd_sc_hd__mux2_4 _27700_ (.A0(_02132_),
    .A1(_02131_),
    .S(_02069_),
    .X(\cpuregs_wrdata[31] ));
 sky130_fd_sc_hd__mux2_1 _27701_ (.A0(_02316_),
    .A1(_02317_),
    .S(_00307_),
    .X(_00004_));
 sky130_fd_sc_hd__mux2_1 _27702_ (.A0(_00347_),
    .A1(_14286_),
    .S(_00336_),
    .X(_00348_));
 sky130_fd_sc_hd__mux2_1 _27703_ (.A0(_14286_),
    .A1(_00348_),
    .S(net101),
    .X(_00003_));
 sky130_fd_sc_hd__mux2_1 _27704_ (.A0(_02304_),
    .A1(_02305_),
    .S(\irq_state[1] ),
    .X(_02306_));
 sky130_fd_sc_hd__mux2_1 _27705_ (.A0(_02306_),
    .A1(_02304_),
    .S(_02217_),
    .X(_00008_));
 sky130_fd_sc_hd__mux2_1 _27706_ (.A0(_02214_),
    .A1(_02215_),
    .S(\irq_state[1] ),
    .X(_02216_));
 sky130_fd_sc_hd__mux2_1 _27707_ (.A0(_02216_),
    .A1(_02214_),
    .S(_02217_),
    .X(_00031_));
 sky130_fd_sc_hd__mux2_1 _27708_ (.A0(_02218_),
    .A1(_02219_),
    .S(\irq_state[1] ),
    .X(_02220_));
 sky130_fd_sc_hd__mux2_1 _27709_ (.A0(_02220_),
    .A1(_02218_),
    .S(_02217_),
    .X(_00032_));
 sky130_fd_sc_hd__mux2_1 _27710_ (.A0(_02221_),
    .A1(_02222_),
    .S(\irq_state[1] ),
    .X(_02223_));
 sky130_fd_sc_hd__mux2_1 _27711_ (.A0(_02223_),
    .A1(_02221_),
    .S(_02217_),
    .X(_00033_));
 sky130_fd_sc_hd__mux2_1 _27712_ (.A0(_02224_),
    .A1(_02225_),
    .S(\irq_state[1] ),
    .X(_02226_));
 sky130_fd_sc_hd__mux2_1 _27713_ (.A0(_02226_),
    .A1(_02224_),
    .S(_02217_),
    .X(_00034_));
 sky130_fd_sc_hd__mux2_1 _27714_ (.A0(_02227_),
    .A1(_02228_),
    .S(\irq_state[1] ),
    .X(_02229_));
 sky130_fd_sc_hd__mux2_1 _27715_ (.A0(_02229_),
    .A1(_02227_),
    .S(_02217_),
    .X(_00035_));
 sky130_fd_sc_hd__mux2_1 _27716_ (.A0(_02230_),
    .A1(_02231_),
    .S(\irq_state[1] ),
    .X(_02232_));
 sky130_fd_sc_hd__mux2_1 _27717_ (.A0(_02232_),
    .A1(_02230_),
    .S(_02217_),
    .X(_00036_));
 sky130_fd_sc_hd__mux2_1 _27718_ (.A0(_02233_),
    .A1(_02234_),
    .S(\irq_state[1] ),
    .X(_02235_));
 sky130_fd_sc_hd__mux2_1 _27719_ (.A0(_02235_),
    .A1(_02233_),
    .S(_02217_),
    .X(_00037_));
 sky130_fd_sc_hd__mux2_1 _27720_ (.A0(_02236_),
    .A1(_02237_),
    .S(\irq_state[1] ),
    .X(_02238_));
 sky130_fd_sc_hd__mux2_1 _27721_ (.A0(_02238_),
    .A1(_02236_),
    .S(_02217_),
    .X(_00009_));
 sky130_fd_sc_hd__mux2_1 _27722_ (.A0(_02239_),
    .A1(_02240_),
    .S(\irq_state[1] ),
    .X(_02241_));
 sky130_fd_sc_hd__mux2_1 _27723_ (.A0(_02241_),
    .A1(_02239_),
    .S(_02217_),
    .X(_00010_));
 sky130_fd_sc_hd__mux2_1 _27724_ (.A0(_02242_),
    .A1(_02243_),
    .S(\irq_state[1] ),
    .X(_02244_));
 sky130_fd_sc_hd__mux2_1 _27725_ (.A0(_02244_),
    .A1(_02242_),
    .S(_02217_),
    .X(_00011_));
 sky130_fd_sc_hd__mux2_1 _27726_ (.A0(_02245_),
    .A1(_02246_),
    .S(\irq_state[1] ),
    .X(_02247_));
 sky130_fd_sc_hd__mux2_1 _27727_ (.A0(_02247_),
    .A1(_02245_),
    .S(_02217_),
    .X(_00012_));
 sky130_fd_sc_hd__mux2_1 _27728_ (.A0(_02248_),
    .A1(_02249_),
    .S(\irq_state[1] ),
    .X(_02250_));
 sky130_fd_sc_hd__mux2_1 _27729_ (.A0(_02250_),
    .A1(_02248_),
    .S(_02217_),
    .X(_00013_));
 sky130_fd_sc_hd__mux2_1 _27730_ (.A0(_02251_),
    .A1(_02252_),
    .S(\irq_state[1] ),
    .X(_02253_));
 sky130_fd_sc_hd__mux2_1 _27731_ (.A0(_02253_),
    .A1(_02251_),
    .S(_02217_),
    .X(_00014_));
 sky130_fd_sc_hd__mux2_1 _27732_ (.A0(_02254_),
    .A1(_02255_),
    .S(\irq_state[1] ),
    .X(_02256_));
 sky130_fd_sc_hd__mux2_1 _27733_ (.A0(_02256_),
    .A1(_02254_),
    .S(_02217_),
    .X(_00015_));
 sky130_fd_sc_hd__mux2_1 _27734_ (.A0(_02257_),
    .A1(_02258_),
    .S(\irq_state[1] ),
    .X(_02259_));
 sky130_fd_sc_hd__mux2_1 _27735_ (.A0(_02259_),
    .A1(_02257_),
    .S(_02217_),
    .X(_00016_));
 sky130_fd_sc_hd__mux2_1 _27736_ (.A0(_02260_),
    .A1(_02261_),
    .S(\irq_state[1] ),
    .X(_02262_));
 sky130_fd_sc_hd__mux2_1 _27737_ (.A0(_02262_),
    .A1(_02260_),
    .S(_02217_),
    .X(_00017_));
 sky130_fd_sc_hd__mux2_1 _27738_ (.A0(_02263_),
    .A1(_02264_),
    .S(\irq_state[1] ),
    .X(_02265_));
 sky130_fd_sc_hd__mux2_1 _27739_ (.A0(_02265_),
    .A1(_02263_),
    .S(_02217_),
    .X(_00018_));
 sky130_fd_sc_hd__mux2_1 _27740_ (.A0(_02266_),
    .A1(_02267_),
    .S(\irq_state[1] ),
    .X(_02268_));
 sky130_fd_sc_hd__mux2_1 _27741_ (.A0(_02268_),
    .A1(_02266_),
    .S(_02217_),
    .X(_00019_));
 sky130_fd_sc_hd__mux2_1 _27742_ (.A0(_02269_),
    .A1(_02270_),
    .S(\irq_state[1] ),
    .X(_02271_));
 sky130_fd_sc_hd__mux2_1 _27743_ (.A0(_02271_),
    .A1(_02269_),
    .S(_02217_),
    .X(_00020_));
 sky130_fd_sc_hd__mux2_1 _27744_ (.A0(_02272_),
    .A1(_02273_),
    .S(\irq_state[1] ),
    .X(_02274_));
 sky130_fd_sc_hd__mux2_1 _27745_ (.A0(_02274_),
    .A1(_02272_),
    .S(_02217_),
    .X(_00021_));
 sky130_fd_sc_hd__mux2_1 _27746_ (.A0(_02275_),
    .A1(_02276_),
    .S(\irq_state[1] ),
    .X(_02277_));
 sky130_fd_sc_hd__mux2_1 _27747_ (.A0(_02277_),
    .A1(_02275_),
    .S(_02217_),
    .X(_00022_));
 sky130_fd_sc_hd__mux2_1 _27748_ (.A0(_02278_),
    .A1(_02279_),
    .S(\irq_state[1] ),
    .X(_02280_));
 sky130_fd_sc_hd__mux2_1 _27749_ (.A0(_02280_),
    .A1(_02278_),
    .S(_02217_),
    .X(_00023_));
 sky130_fd_sc_hd__mux2_1 _27750_ (.A0(_02281_),
    .A1(_02282_),
    .S(\irq_state[1] ),
    .X(_02283_));
 sky130_fd_sc_hd__mux2_1 _27751_ (.A0(_02283_),
    .A1(_02281_),
    .S(_02217_),
    .X(_00024_));
 sky130_fd_sc_hd__mux2_1 _27752_ (.A0(_02284_),
    .A1(_02285_),
    .S(\irq_state[1] ),
    .X(_02286_));
 sky130_fd_sc_hd__mux2_1 _27753_ (.A0(_02286_),
    .A1(_02284_),
    .S(_02217_),
    .X(_00025_));
 sky130_fd_sc_hd__mux2_1 _27754_ (.A0(_02287_),
    .A1(_02288_),
    .S(\irq_state[1] ),
    .X(_02289_));
 sky130_fd_sc_hd__mux2_1 _27755_ (.A0(_02289_),
    .A1(_02287_),
    .S(_02217_),
    .X(_00026_));
 sky130_fd_sc_hd__mux2_1 _27756_ (.A0(_02290_),
    .A1(_02291_),
    .S(\irq_state[1] ),
    .X(_02292_));
 sky130_fd_sc_hd__mux2_1 _27757_ (.A0(_02292_),
    .A1(_02290_),
    .S(_02217_),
    .X(_00027_));
 sky130_fd_sc_hd__mux2_1 _27758_ (.A0(_02293_),
    .A1(_02294_),
    .S(\irq_state[1] ),
    .X(_02295_));
 sky130_fd_sc_hd__mux2_1 _27759_ (.A0(_02295_),
    .A1(_02293_),
    .S(_02217_),
    .X(_00028_));
 sky130_fd_sc_hd__mux2_1 _27760_ (.A0(_02296_),
    .A1(_02297_),
    .S(\irq_state[1] ),
    .X(_02298_));
 sky130_fd_sc_hd__mux2_1 _27761_ (.A0(_02298_),
    .A1(_02296_),
    .S(_02217_),
    .X(_00029_));
 sky130_fd_sc_hd__mux2_1 _27762_ (.A0(_02299_),
    .A1(_02300_),
    .S(\irq_state[1] ),
    .X(_02301_));
 sky130_fd_sc_hd__mux2_1 _27763_ (.A0(_02301_),
    .A1(_02299_),
    .S(_02217_),
    .X(_00030_));
 sky130_fd_sc_hd__mux2_2 _27764_ (.A0(_01467_),
    .A1(\reg_next_pc[1] ),
    .S(net425),
    .X(_02590_));
 sky130_fd_sc_hd__mux2_1 _27765_ (.A0(_00295_),
    .A1(\reg_next_pc[2] ),
    .S(net425),
    .X(_02560_));
 sky130_fd_sc_hd__mux2_4 _27766_ (.A0(_01470_),
    .A1(\reg_next_pc[3] ),
    .S(net425),
    .X(_02571_));
 sky130_fd_sc_hd__mux2_2 _27767_ (.A0(_01478_),
    .A1(\reg_next_pc[5] ),
    .S(net425),
    .X(_02583_));
 sky130_fd_sc_hd__mux2_2 _27768_ (.A0(_01481_),
    .A1(\reg_next_pc[6] ),
    .S(net425),
    .X(_02584_));
 sky130_fd_sc_hd__mux2_2 _27769_ (.A0(_01484_),
    .A1(\reg_next_pc[7] ),
    .S(net425),
    .X(_02585_));
 sky130_fd_sc_hd__mux2_2 _27770_ (.A0(_01487_),
    .A1(\reg_next_pc[8] ),
    .S(net425),
    .X(_02586_));
 sky130_fd_sc_hd__mux2_2 _27771_ (.A0(_01490_),
    .A1(\reg_next_pc[9] ),
    .S(net425),
    .X(_02587_));
 sky130_fd_sc_hd__mux2_2 _27772_ (.A0(_01493_),
    .A1(\reg_next_pc[10] ),
    .S(net425),
    .X(_02588_));
 sky130_fd_sc_hd__mux2_2 _27773_ (.A0(_01496_),
    .A1(\reg_next_pc[11] ),
    .S(net425),
    .X(_02589_));
 sky130_fd_sc_hd__mux2_2 _27774_ (.A0(_01499_),
    .A1(\reg_next_pc[12] ),
    .S(net425),
    .X(_02561_));
 sky130_fd_sc_hd__mux2_2 _27775_ (.A0(_01502_),
    .A1(\reg_next_pc[13] ),
    .S(net425),
    .X(_02562_));
 sky130_fd_sc_hd__mux2_2 _27776_ (.A0(_01505_),
    .A1(\reg_next_pc[14] ),
    .S(net425),
    .X(_02563_));
 sky130_fd_sc_hd__mux2_2 _27777_ (.A0(_01508_),
    .A1(\reg_next_pc[15] ),
    .S(net425),
    .X(_02564_));
 sky130_fd_sc_hd__mux2_2 _27778_ (.A0(_01511_),
    .A1(\reg_next_pc[16] ),
    .S(net425),
    .X(_02565_));
 sky130_fd_sc_hd__mux2_2 _27779_ (.A0(_01514_),
    .A1(\reg_next_pc[17] ),
    .S(_00292_),
    .X(_02566_));
 sky130_fd_sc_hd__mux2_2 _27780_ (.A0(_01517_),
    .A1(\reg_next_pc[18] ),
    .S(_00292_),
    .X(_02567_));
 sky130_fd_sc_hd__mux2_2 _27781_ (.A0(_01520_),
    .A1(\reg_next_pc[19] ),
    .S(_00292_),
    .X(_02568_));
 sky130_fd_sc_hd__mux2_2 _27782_ (.A0(_01523_),
    .A1(\reg_next_pc[20] ),
    .S(_00292_),
    .X(_02569_));
 sky130_fd_sc_hd__mux2_2 _27783_ (.A0(_01526_),
    .A1(\reg_next_pc[21] ),
    .S(_00292_),
    .X(_02570_));
 sky130_fd_sc_hd__mux2_2 _27784_ (.A0(_01529_),
    .A1(\reg_next_pc[22] ),
    .S(_00292_),
    .X(_02572_));
 sky130_fd_sc_hd__mux2_4 _27785_ (.A0(_01532_),
    .A1(\reg_next_pc[23] ),
    .S(_00292_),
    .X(_02573_));
 sky130_fd_sc_hd__mux2_2 _27786_ (.A0(_01535_),
    .A1(\reg_next_pc[24] ),
    .S(_00292_),
    .X(_02574_));
 sky130_fd_sc_hd__mux2_2 _27787_ (.A0(_01538_),
    .A1(\reg_next_pc[25] ),
    .S(_00292_),
    .X(_02575_));
 sky130_fd_sc_hd__mux2_2 _27788_ (.A0(_01541_),
    .A1(\reg_next_pc[26] ),
    .S(_00292_),
    .X(_02576_));
 sky130_fd_sc_hd__mux2_2 _27789_ (.A0(_01544_),
    .A1(\reg_next_pc[27] ),
    .S(_00292_),
    .X(_02577_));
 sky130_fd_sc_hd__mux2_2 _27790_ (.A0(_01547_),
    .A1(\reg_next_pc[28] ),
    .S(_00292_),
    .X(_02578_));
 sky130_fd_sc_hd__mux2_2 _27791_ (.A0(_01550_),
    .A1(\reg_next_pc[29] ),
    .S(_00292_),
    .X(_02579_));
 sky130_fd_sc_hd__mux2_2 _27792_ (.A0(_01553_),
    .A1(\reg_next_pc[30] ),
    .S(_00292_),
    .X(_02580_));
 sky130_fd_sc_hd__mux2_2 _27793_ (.A0(_01556_),
    .A1(\reg_next_pc[31] ),
    .S(_00292_),
    .X(_02581_));
 sky130_fd_sc_hd__mux2_1 _27794_ (.A0(_00057_),
    .A1(_00064_),
    .S(net225),
    .X(_00065_));
 sky130_fd_sc_hd__mux2_1 _27795_ (.A0(_00065_),
    .A1(_02543_),
    .S(net458),
    .X(_14322_));
 sky130_fd_sc_hd__mux2_1 _27796_ (.A0(_00075_),
    .A1(_00082_),
    .S(net225),
    .X(_00083_));
 sky130_fd_sc_hd__mux2_2 _27797_ (.A0(_00083_),
    .A1(_02544_),
    .S(net226),
    .X(_14323_));
 sky130_fd_sc_hd__mux2_1 _27798_ (.A0(_00089_),
    .A1(_00092_),
    .S(net225),
    .X(_00093_));
 sky130_fd_sc_hd__mux2_2 _27799_ (.A0(_00093_),
    .A1(_02545_),
    .S(net458),
    .X(_14324_));
 sky130_fd_sc_hd__mux2_1 _27800_ (.A0(_00099_),
    .A1(_00102_),
    .S(net225),
    .X(_00103_));
 sky130_fd_sc_hd__mux2_1 _27801_ (.A0(_00103_),
    .A1(_02546_),
    .S(net226),
    .X(_14325_));
 sky130_fd_sc_hd__mux2_1 _27802_ (.A0(_00107_),
    .A1(_00108_),
    .S(net225),
    .X(_00109_));
 sky130_fd_sc_hd__mux2_1 _27803_ (.A0(_00109_),
    .A1(_02547_),
    .S(net458),
    .X(_14326_));
 sky130_fd_sc_hd__mux2_1 _27804_ (.A0(_00113_),
    .A1(_00114_),
    .S(net459),
    .X(_00115_));
 sky130_fd_sc_hd__mux2_2 _27805_ (.A0(_00115_),
    .A1(_02548_),
    .S(net226),
    .X(_14327_));
 sky130_fd_sc_hd__mux2_1 _27806_ (.A0(_00119_),
    .A1(_00120_),
    .S(net459),
    .X(_00121_));
 sky130_fd_sc_hd__mux2_1 _27807_ (.A0(_00121_),
    .A1(_02549_),
    .S(net226),
    .X(_14328_));
 sky130_fd_sc_hd__mux2_1 _27808_ (.A0(_00125_),
    .A1(_00126_),
    .S(net459),
    .X(_00127_));
 sky130_fd_sc_hd__mux2_2 _27809_ (.A0(_00127_),
    .A1(_02550_),
    .S(net226),
    .X(_14329_));
 sky130_fd_sc_hd__mux2_1 _27810_ (.A0(_00129_),
    .A1(_00106_),
    .S(net460),
    .X(_00130_));
 sky130_fd_sc_hd__mux2_1 _27811_ (.A0(_00130_),
    .A1(_00057_),
    .S(net459),
    .X(_00131_));
 sky130_fd_sc_hd__mux2_1 _27812_ (.A0(_00131_),
    .A1(_02551_),
    .S(net226),
    .X(_14330_));
 sky130_fd_sc_hd__mux2_1 _27813_ (.A0(_00133_),
    .A1(_00112_),
    .S(net222),
    .X(_00134_));
 sky130_fd_sc_hd__mux2_1 _27814_ (.A0(_00134_),
    .A1(_00075_),
    .S(net459),
    .X(_00135_));
 sky130_fd_sc_hd__mux2_1 _27815_ (.A0(_00135_),
    .A1(_02552_),
    .S(net226),
    .X(_14331_));
 sky130_fd_sc_hd__mux2_1 _27816_ (.A0(_00137_),
    .A1(_00118_),
    .S(net460),
    .X(_00138_));
 sky130_fd_sc_hd__mux2_1 _27817_ (.A0(_00138_),
    .A1(_00089_),
    .S(net459),
    .X(_00139_));
 sky130_fd_sc_hd__mux2_1 _27818_ (.A0(_00139_),
    .A1(_02553_),
    .S(net458),
    .X(_14332_));
 sky130_fd_sc_hd__mux2_1 _27819_ (.A0(_00141_),
    .A1(_00124_),
    .S(net222),
    .X(_00142_));
 sky130_fd_sc_hd__mux2_1 _27820_ (.A0(_00142_),
    .A1(_00099_),
    .S(net459),
    .X(_00143_));
 sky130_fd_sc_hd__mux2_1 _27821_ (.A0(_00143_),
    .A1(_02554_),
    .S(net226),
    .X(_14333_));
 sky130_fd_sc_hd__mux2_1 _27822_ (.A0(_00144_),
    .A1(_00136_),
    .S(net461),
    .X(_00145_));
 sky130_fd_sc_hd__mux2_1 _27823_ (.A0(_00145_),
    .A1(_00129_),
    .S(net460),
    .X(_00146_));
 sky130_fd_sc_hd__mux2_1 _27824_ (.A0(_00146_),
    .A1(_00107_),
    .S(net459),
    .X(_00147_));
 sky130_fd_sc_hd__mux2_1 _27825_ (.A0(_00147_),
    .A1(_02555_),
    .S(net458),
    .X(_14334_));
 sky130_fd_sc_hd__mux2_1 _27826_ (.A0(_00148_),
    .A1(_00140_),
    .S(net461),
    .X(_00149_));
 sky130_fd_sc_hd__mux2_1 _27827_ (.A0(_00149_),
    .A1(_00133_),
    .S(net222),
    .X(_00150_));
 sky130_fd_sc_hd__mux2_1 _27828_ (.A0(_00150_),
    .A1(_00113_),
    .S(net459),
    .X(_00151_));
 sky130_fd_sc_hd__mux2_1 _27829_ (.A0(_00151_),
    .A1(_02556_),
    .S(net226),
    .X(_14335_));
 sky130_fd_sc_hd__mux2_1 _27830_ (.A0(net329),
    .A1(net327),
    .S(net462),
    .X(_00152_));
 sky130_fd_sc_hd__mux2_1 _27831_ (.A0(_00152_),
    .A1(_00144_),
    .S(net461),
    .X(_00153_));
 sky130_fd_sc_hd__mux2_1 _27832_ (.A0(_00153_),
    .A1(_00137_),
    .S(net460),
    .X(_00154_));
 sky130_fd_sc_hd__mux2_1 _27833_ (.A0(_00154_),
    .A1(_00119_),
    .S(net459),
    .X(_00155_));
 sky130_fd_sc_hd__mux2_1 _27834_ (.A0(_00155_),
    .A1(_02557_),
    .S(net458),
    .X(_14336_));
 sky130_fd_sc_hd__mux2_1 _27835_ (.A0(net330),
    .A1(net329),
    .S(net200),
    .X(_00156_));
 sky130_fd_sc_hd__mux2_1 _27836_ (.A0(_00156_),
    .A1(_00148_),
    .S(net461),
    .X(_00157_));
 sky130_fd_sc_hd__mux2_1 _27837_ (.A0(_00157_),
    .A1(_00141_),
    .S(net222),
    .X(_00158_));
 sky130_fd_sc_hd__mux2_1 _27838_ (.A0(_00158_),
    .A1(_00125_),
    .S(net459),
    .X(_00159_));
 sky130_fd_sc_hd__mux2_1 _27839_ (.A0(_00159_),
    .A1(_02558_),
    .S(net226),
    .X(_14337_));
 sky130_fd_sc_hd__mux2_1 _27840_ (.A0(net306),
    .A1(net317),
    .S(net200),
    .X(_00160_));
 sky130_fd_sc_hd__mux2_1 _27841_ (.A0(_00160_),
    .A1(_00161_),
    .S(net461),
    .X(_00162_));
 sky130_fd_sc_hd__mux2_1 _27842_ (.A0(_00162_),
    .A1(_00165_),
    .S(net460),
    .X(_00166_));
 sky130_fd_sc_hd__mux2_1 _27843_ (.A0(_00166_),
    .A1(_00173_),
    .S(net459),
    .X(_00174_));
 sky130_fd_sc_hd__mux2_1 _27844_ (.A0(_00174_),
    .A1(_00189_),
    .S(net458),
    .X(_14338_));
 sky130_fd_sc_hd__mux2_1 _27845_ (.A0(net317),
    .A1(net328),
    .S(net200),
    .X(_00190_));
 sky130_fd_sc_hd__mux2_1 _27846_ (.A0(_00190_),
    .A1(_00191_),
    .S(net461),
    .X(_00192_));
 sky130_fd_sc_hd__mux2_1 _27847_ (.A0(_00192_),
    .A1(_00195_),
    .S(net222),
    .X(_00196_));
 sky130_fd_sc_hd__mux2_1 _27848_ (.A0(_00196_),
    .A1(_00203_),
    .S(net459),
    .X(_00204_));
 sky130_fd_sc_hd__mux2_1 _27849_ (.A0(_00204_),
    .A1(_00220_),
    .S(net458),
    .X(_14349_));
 sky130_fd_sc_hd__mux2_1 _27850_ (.A0(_00161_),
    .A1(_00163_),
    .S(net461),
    .X(_00221_));
 sky130_fd_sc_hd__mux2_1 _27851_ (.A0(_00221_),
    .A1(_00222_),
    .S(net460),
    .X(_00223_));
 sky130_fd_sc_hd__mux2_1 _27852_ (.A0(_00223_),
    .A1(_00226_),
    .S(net459),
    .X(_00227_));
 sky130_fd_sc_hd__mux2_1 _27853_ (.A0(_00227_),
    .A1(_00234_),
    .S(net458),
    .X(_14360_));
 sky130_fd_sc_hd__mux2_1 _27854_ (.A0(_00191_),
    .A1(_00193_),
    .S(net461),
    .X(_00235_));
 sky130_fd_sc_hd__mux2_1 _27855_ (.A0(_00235_),
    .A1(_00236_),
    .S(net222),
    .X(_00237_));
 sky130_fd_sc_hd__mux2_1 _27856_ (.A0(_00237_),
    .A1(_00240_),
    .S(net459),
    .X(_00241_));
 sky130_fd_sc_hd__mux2_1 _27857_ (.A0(_00241_),
    .A1(_00248_),
    .S(net458),
    .X(_14363_));
 sky130_fd_sc_hd__mux2_1 _27858_ (.A0(_00165_),
    .A1(_00169_),
    .S(net460),
    .X(_00249_));
 sky130_fd_sc_hd__mux2_1 _27859_ (.A0(_00249_),
    .A1(_00250_),
    .S(net459),
    .X(_00251_));
 sky130_fd_sc_hd__mux2_1 _27860_ (.A0(_00251_),
    .A1(_00254_),
    .S(net458),
    .X(_14364_));
 sky130_fd_sc_hd__mux2_1 _27861_ (.A0(_00195_),
    .A1(_00199_),
    .S(net222),
    .X(_00255_));
 sky130_fd_sc_hd__mux2_1 _27862_ (.A0(_00255_),
    .A1(_00256_),
    .S(net459),
    .X(_00257_));
 sky130_fd_sc_hd__mux2_1 _27863_ (.A0(_00257_),
    .A1(_00260_),
    .S(net458),
    .X(_14365_));
 sky130_fd_sc_hd__mux2_1 _27864_ (.A0(_00222_),
    .A1(_00224_),
    .S(net460),
    .X(_00261_));
 sky130_fd_sc_hd__mux2_1 _27865_ (.A0(_00261_),
    .A1(_00262_),
    .S(net459),
    .X(_00263_));
 sky130_fd_sc_hd__mux2_1 _27866_ (.A0(_00263_),
    .A1(_00266_),
    .S(net458),
    .X(_14366_));
 sky130_fd_sc_hd__mux2_1 _27867_ (.A0(_00236_),
    .A1(_00238_),
    .S(net222),
    .X(_00267_));
 sky130_fd_sc_hd__mux2_1 _27868_ (.A0(_00267_),
    .A1(_00268_),
    .S(net459),
    .X(_00269_));
 sky130_fd_sc_hd__mux2_1 _27869_ (.A0(_00269_),
    .A1(_00272_),
    .S(net458),
    .X(_14367_));
 sky130_fd_sc_hd__mux2_1 _27870_ (.A0(_00173_),
    .A1(_00181_),
    .S(net459),
    .X(_00273_));
 sky130_fd_sc_hd__mux2_1 _27871_ (.A0(_00273_),
    .A1(_00274_),
    .S(net458),
    .X(_14368_));
 sky130_fd_sc_hd__mux2_1 _27872_ (.A0(_00203_),
    .A1(_00211_),
    .S(net459),
    .X(_00275_));
 sky130_fd_sc_hd__mux2_1 _27873_ (.A0(_00275_),
    .A1(_00276_),
    .S(net458),
    .X(_14369_));
 sky130_fd_sc_hd__mux2_1 _27874_ (.A0(_00226_),
    .A1(_00230_),
    .S(net459),
    .X(_00277_));
 sky130_fd_sc_hd__mux2_1 _27875_ (.A0(_00277_),
    .A1(_00278_),
    .S(net458),
    .X(_14339_));
 sky130_fd_sc_hd__mux2_1 _27876_ (.A0(_00240_),
    .A1(_00244_),
    .S(net459),
    .X(_00279_));
 sky130_fd_sc_hd__mux2_1 _27877_ (.A0(_00279_),
    .A1(_00280_),
    .S(net458),
    .X(_14340_));
 sky130_fd_sc_hd__mux2_1 _27878_ (.A0(_00250_),
    .A1(_00252_),
    .S(net459),
    .X(_00281_));
 sky130_fd_sc_hd__mux2_1 _27879_ (.A0(_00281_),
    .A1(_00282_),
    .S(net458),
    .X(_14341_));
 sky130_fd_sc_hd__mux2_1 _27880_ (.A0(_00256_),
    .A1(_00258_),
    .S(net459),
    .X(_00283_));
 sky130_fd_sc_hd__mux2_1 _27881_ (.A0(_00283_),
    .A1(_00284_),
    .S(net458),
    .X(_14342_));
 sky130_fd_sc_hd__mux2_1 _27882_ (.A0(_00262_),
    .A1(_00264_),
    .S(net459),
    .X(_00285_));
 sky130_fd_sc_hd__mux2_1 _27883_ (.A0(_00285_),
    .A1(_00286_),
    .S(net458),
    .X(_14343_));
 sky130_fd_sc_hd__mux2_1 _27884_ (.A0(_00268_),
    .A1(_00270_),
    .S(net459),
    .X(_00287_));
 sky130_fd_sc_hd__mux2_1 _27885_ (.A0(_00287_),
    .A1(_00288_),
    .S(net458),
    .X(_14344_));
 sky130_fd_sc_hd__mux2_1 _27886_ (.A0(_00189_),
    .A1(_00216_),
    .S(net458),
    .X(_14345_));
 sky130_fd_sc_hd__mux2_1 _27887_ (.A0(_00220_),
    .A1(_00216_),
    .S(net458),
    .X(_14346_));
 sky130_fd_sc_hd__mux2_1 _27888_ (.A0(_00234_),
    .A1(_00216_),
    .S(net458),
    .X(_14347_));
 sky130_fd_sc_hd__mux2_1 _27889_ (.A0(_00248_),
    .A1(_00216_),
    .S(net458),
    .X(_14348_));
 sky130_fd_sc_hd__mux2_1 _27890_ (.A0(_00254_),
    .A1(_00216_),
    .S(net458),
    .X(_14350_));
 sky130_fd_sc_hd__mux2_1 _27891_ (.A0(_00260_),
    .A1(_00216_),
    .S(net458),
    .X(_14351_));
 sky130_fd_sc_hd__mux2_1 _27892_ (.A0(_00266_),
    .A1(_00216_),
    .S(net458),
    .X(_14352_));
 sky130_fd_sc_hd__mux2_1 _27893_ (.A0(_00272_),
    .A1(_00216_),
    .S(net458),
    .X(_14353_));
 sky130_fd_sc_hd__mux2_1 _27894_ (.A0(_00274_),
    .A1(_00216_),
    .S(net458),
    .X(_14354_));
 sky130_fd_sc_hd__mux2_1 _27895_ (.A0(_00276_),
    .A1(_00216_),
    .S(net458),
    .X(_14355_));
 sky130_fd_sc_hd__mux2_1 _27896_ (.A0(_00278_),
    .A1(_00216_),
    .S(net458),
    .X(_14356_));
 sky130_fd_sc_hd__mux2_1 _27897_ (.A0(_00280_),
    .A1(_00216_),
    .S(net458),
    .X(_14357_));
 sky130_fd_sc_hd__mux2_1 _27898_ (.A0(_00282_),
    .A1(_00216_),
    .S(net458),
    .X(_14358_));
 sky130_fd_sc_hd__mux2_1 _27899_ (.A0(_00284_),
    .A1(_00216_),
    .S(net458),
    .X(_14359_));
 sky130_fd_sc_hd__mux2_1 _27900_ (.A0(_00286_),
    .A1(_00216_),
    .S(net458),
    .X(_14361_));
 sky130_fd_sc_hd__mux2_1 _27901_ (.A0(_00288_),
    .A1(_00216_),
    .S(net458),
    .X(_14362_));
 sky130_fd_sc_hd__mux2_1 _27902_ (.A0(_01697_),
    .A1(_01698_),
    .S(\irq_state[1] ),
    .X(_01699_));
 sky130_fd_sc_hd__mux2_1 _27903_ (.A0(_01705_),
    .A1(_01699_),
    .S(_01700_),
    .X(_14321_));
 sky130_fd_sc_hd__mux2_1 _27904_ (.A0(_01720_),
    .A1(\irq_pending[0] ),
    .S(_01706_),
    .X(_14287_));
 sky130_fd_sc_hd__mux2_1 _27905_ (.A0(_01733_),
    .A1(\irq_pending[1] ),
    .S(_01706_),
    .X(_14298_));
 sky130_fd_sc_hd__mux2_1 _27906_ (.A0(_01746_),
    .A1(\irq_pending[2] ),
    .S(_01706_),
    .X(_14309_));
 sky130_fd_sc_hd__mux2_1 _27907_ (.A0(_01759_),
    .A1(\irq_pending[3] ),
    .S(_01706_),
    .X(_14312_));
 sky130_fd_sc_hd__mux2_1 _27908_ (.A0(_01772_),
    .A1(\irq_pending[4] ),
    .S(_01706_),
    .X(_14313_));
 sky130_fd_sc_hd__mux2_1 _27909_ (.A0(_01785_),
    .A1(\irq_pending[5] ),
    .S(_01706_),
    .X(_14314_));
 sky130_fd_sc_hd__mux2_1 _27910_ (.A0(_01798_),
    .A1(\irq_pending[6] ),
    .S(_01706_),
    .X(_14315_));
 sky130_fd_sc_hd__mux2_1 _27911_ (.A0(_01811_),
    .A1(\irq_pending[7] ),
    .S(_01706_),
    .X(_14316_));
 sky130_fd_sc_hd__mux2_1 _27912_ (.A0(_01825_),
    .A1(\irq_pending[8] ),
    .S(_01706_),
    .X(_14317_));
 sky130_fd_sc_hd__mux2_1 _27913_ (.A0(_01838_),
    .A1(\irq_pending[9] ),
    .S(_01706_),
    .X(_14318_));
 sky130_fd_sc_hd__mux2_1 _27914_ (.A0(_01851_),
    .A1(\irq_pending[10] ),
    .S(_01706_),
    .X(_14288_));
 sky130_fd_sc_hd__mux2_1 _27915_ (.A0(_01864_),
    .A1(\irq_pending[11] ),
    .S(_01706_),
    .X(_14289_));
 sky130_fd_sc_hd__mux2_1 _27916_ (.A0(_01877_),
    .A1(\irq_pending[12] ),
    .S(_01706_),
    .X(_14290_));
 sky130_fd_sc_hd__mux2_1 _27917_ (.A0(_01890_),
    .A1(\irq_pending[13] ),
    .S(_01706_),
    .X(_14291_));
 sky130_fd_sc_hd__mux2_1 _27918_ (.A0(_01903_),
    .A1(\irq_pending[14] ),
    .S(_01706_),
    .X(_14292_));
 sky130_fd_sc_hd__mux2_1 _27919_ (.A0(_01916_),
    .A1(\irq_pending[15] ),
    .S(_01706_),
    .X(_14293_));
 sky130_fd_sc_hd__mux2_1 _27920_ (.A0(_01925_),
    .A1(\irq_pending[16] ),
    .S(_01706_),
    .X(_14294_));
 sky130_fd_sc_hd__mux2_1 _27921_ (.A0(_01934_),
    .A1(\irq_pending[17] ),
    .S(_01706_),
    .X(_14295_));
 sky130_fd_sc_hd__mux2_1 _27922_ (.A0(_01943_),
    .A1(\irq_pending[18] ),
    .S(_01706_),
    .X(_14296_));
 sky130_fd_sc_hd__mux2_1 _27923_ (.A0(_01952_),
    .A1(\irq_pending[19] ),
    .S(_01706_),
    .X(_14297_));
 sky130_fd_sc_hd__mux2_1 _27924_ (.A0(_01961_),
    .A1(\irq_pending[20] ),
    .S(_01706_),
    .X(_14299_));
 sky130_fd_sc_hd__mux2_1 _27925_ (.A0(_01970_),
    .A1(\irq_pending[21] ),
    .S(_01706_),
    .X(_14300_));
 sky130_fd_sc_hd__mux2_1 _27926_ (.A0(_01979_),
    .A1(\irq_pending[22] ),
    .S(_01706_),
    .X(_14301_));
 sky130_fd_sc_hd__mux2_1 _27927_ (.A0(_01988_),
    .A1(\irq_pending[23] ),
    .S(_01706_),
    .X(_14302_));
 sky130_fd_sc_hd__mux2_1 _27928_ (.A0(_01997_),
    .A1(\irq_pending[24] ),
    .S(_01706_),
    .X(_14303_));
 sky130_fd_sc_hd__mux2_1 _27929_ (.A0(_02006_),
    .A1(\irq_pending[25] ),
    .S(_01706_),
    .X(_14304_));
 sky130_fd_sc_hd__mux2_1 _27930_ (.A0(_02015_),
    .A1(\irq_pending[26] ),
    .S(_01706_),
    .X(_14305_));
 sky130_fd_sc_hd__mux2_1 _27931_ (.A0(_02024_),
    .A1(\irq_pending[27] ),
    .S(_01706_),
    .X(_14306_));
 sky130_fd_sc_hd__mux2_1 _27932_ (.A0(_02033_),
    .A1(\irq_pending[28] ),
    .S(_01706_),
    .X(_14307_));
 sky130_fd_sc_hd__mux2_1 _27933_ (.A0(_02042_),
    .A1(\irq_pending[29] ),
    .S(_01706_),
    .X(_14308_));
 sky130_fd_sc_hd__mux2_1 _27934_ (.A0(_02051_),
    .A1(\irq_pending[30] ),
    .S(_01706_),
    .X(_14310_));
 sky130_fd_sc_hd__mux2_1 _27935_ (.A0(_02060_),
    .A1(\irq_pending[31] ),
    .S(_01706_),
    .X(_14311_));
 sky130_fd_sc_hd__mux2_4 _27936_ (.A0(_02061_),
    .A1(\cpu_state[2] ),
    .S(_02542_),
    .X(_14282_));
 sky130_fd_sc_hd__mux2_2 _27937_ (.A0(\decoded_rd[0] ),
    .A1(\irq_state[0] ),
    .S(net410),
    .X(_14281_));
 sky130_fd_sc_hd__mux2_1 _27938_ (.A0(_02062_),
    .A1(_02065_),
    .S(_02542_),
    .X(_14319_));
 sky130_fd_sc_hd__mux2_1 _27939_ (.A0(_02068_),
    .A1(_02066_),
    .S(_02067_),
    .X(_14320_));
 sky130_fd_sc_hd__mux2_1 _27940_ (.A0(_02166_),
    .A1(_00291_),
    .S(_00290_),
    .X(_14283_));
 sky130_fd_sc_hd__mux2_1 _27941_ (.A0(_02166_),
    .A1(mem_do_wdata),
    .S(_00290_),
    .X(_14284_));
 sky130_fd_sc_hd__mux2_1 _27942_ (.A0(_00271_),
    .A1(_00216_),
    .S(net459),
    .X(_00288_));
 sky130_fd_sc_hd__mux2_1 _27943_ (.A0(_00265_),
    .A1(_00216_),
    .S(net459),
    .X(_00286_));
 sky130_fd_sc_hd__mux2_1 _27944_ (.A0(_00259_),
    .A1(_00216_),
    .S(net459),
    .X(_00284_));
 sky130_fd_sc_hd__mux2_1 _27945_ (.A0(_00253_),
    .A1(_00216_),
    .S(net459),
    .X(_00282_));
 sky130_fd_sc_hd__mux2_1 _27946_ (.A0(_00247_),
    .A1(_00216_),
    .S(net459),
    .X(_00280_));
 sky130_fd_sc_hd__mux2_1 _27947_ (.A0(_00233_),
    .A1(_00216_),
    .S(net459),
    .X(_00278_));
 sky130_fd_sc_hd__mux2_1 _27948_ (.A0(_00219_),
    .A1(_00216_),
    .S(net459),
    .X(_00276_));
 sky130_fd_sc_hd__mux2_1 _27949_ (.A0(_00188_),
    .A1(_00216_),
    .S(net459),
    .X(_00274_));
 sky130_fd_sc_hd__mux2_1 _27950_ (.A0(_00270_),
    .A1(_00271_),
    .S(net459),
    .X(_00272_));
 sky130_fd_sc_hd__mux2_1 _27951_ (.A0(_00246_),
    .A1(_00216_),
    .S(net222),
    .X(_00271_));
 sky130_fd_sc_hd__mux2_1 _27952_ (.A0(_00243_),
    .A1(_00245_),
    .S(net222),
    .X(_00270_));
 sky130_fd_sc_hd__mux2_1 _27953_ (.A0(_00239_),
    .A1(_00242_),
    .S(net222),
    .X(_00268_));
 sky130_fd_sc_hd__mux2_2 _27954_ (.A0(_00264_),
    .A1(_00265_),
    .S(net459),
    .X(_00266_));
 sky130_fd_sc_hd__mux2_1 _27955_ (.A0(_00232_),
    .A1(_00216_),
    .S(net460),
    .X(_00265_));
 sky130_fd_sc_hd__mux2_1 _27956_ (.A0(_00229_),
    .A1(_00231_),
    .S(net460),
    .X(_00264_));
 sky130_fd_sc_hd__mux2_1 _27957_ (.A0(_00225_),
    .A1(_00228_),
    .S(net460),
    .X(_00262_));
 sky130_fd_sc_hd__mux2_1 _27958_ (.A0(_00258_),
    .A1(_00259_),
    .S(net459),
    .X(_00260_));
 sky130_fd_sc_hd__mux2_1 _27959_ (.A0(_00218_),
    .A1(_00216_),
    .S(net222),
    .X(_00259_));
 sky130_fd_sc_hd__mux2_1 _27960_ (.A0(_00210_),
    .A1(_00214_),
    .S(net222),
    .X(_00258_));
 sky130_fd_sc_hd__mux2_1 _27961_ (.A0(_00202_),
    .A1(_00207_),
    .S(net222),
    .X(_00256_));
 sky130_fd_sc_hd__mux2_2 _27962_ (.A0(_00252_),
    .A1(_00253_),
    .S(net459),
    .X(_00254_));
 sky130_fd_sc_hd__mux2_1 _27963_ (.A0(_00187_),
    .A1(_00216_),
    .S(net460),
    .X(_00253_));
 sky130_fd_sc_hd__mux2_1 _27964_ (.A0(_00180_),
    .A1(_00184_),
    .S(net460),
    .X(_00252_));
 sky130_fd_sc_hd__mux2_1 _27965_ (.A0(_00172_),
    .A1(_00177_),
    .S(net460),
    .X(_00250_));
 sky130_fd_sc_hd__mux2_1 _27966_ (.A0(_00244_),
    .A1(_00247_),
    .S(net459),
    .X(_00248_));
 sky130_fd_sc_hd__mux2_1 _27967_ (.A0(_00245_),
    .A1(_00246_),
    .S(net222),
    .X(_00247_));
 sky130_fd_sc_hd__mux2_1 _27968_ (.A0(_00217_),
    .A1(_00216_),
    .S(net461),
    .X(_00246_));
 sky130_fd_sc_hd__mux2_1 _27969_ (.A0(_00213_),
    .A1(_00215_),
    .S(net461),
    .X(_00245_));
 sky130_fd_sc_hd__mux2_1 _27970_ (.A0(_00242_),
    .A1(_00243_),
    .S(net222),
    .X(_00244_));
 sky130_fd_sc_hd__mux2_1 _27971_ (.A0(_00209_),
    .A1(_00212_),
    .S(net461),
    .X(_00243_));
 sky130_fd_sc_hd__mux2_1 _27972_ (.A0(_00206_),
    .A1(_00208_),
    .S(net461),
    .X(_00242_));
 sky130_fd_sc_hd__mux2_1 _27973_ (.A0(_00238_),
    .A1(_00239_),
    .S(net222),
    .X(_00240_));
 sky130_fd_sc_hd__mux2_1 _27974_ (.A0(_00201_),
    .A1(_00205_),
    .S(net461),
    .X(_00239_));
 sky130_fd_sc_hd__mux2_1 _27975_ (.A0(_00198_),
    .A1(_00200_),
    .S(net461),
    .X(_00238_));
 sky130_fd_sc_hd__mux2_1 _27976_ (.A0(_00194_),
    .A1(_00197_),
    .S(net461),
    .X(_00236_));
 sky130_fd_sc_hd__mux2_2 _27977_ (.A0(_00230_),
    .A1(_00233_),
    .S(net459),
    .X(_00234_));
 sky130_fd_sc_hd__mux2_1 _27978_ (.A0(_00231_),
    .A1(_00232_),
    .S(net460),
    .X(_00233_));
 sky130_fd_sc_hd__mux2_1 _27979_ (.A0(_00186_),
    .A1(_00216_),
    .S(net461),
    .X(_00232_));
 sky130_fd_sc_hd__mux2_1 _27980_ (.A0(_00183_),
    .A1(_00185_),
    .S(net461),
    .X(_00231_));
 sky130_fd_sc_hd__mux2_1 _27981_ (.A0(_00228_),
    .A1(_00229_),
    .S(net460),
    .X(_00230_));
 sky130_fd_sc_hd__mux2_1 _27982_ (.A0(_00179_),
    .A1(_00182_),
    .S(net461),
    .X(_00229_));
 sky130_fd_sc_hd__mux2_1 _27983_ (.A0(_00176_),
    .A1(_00178_),
    .S(net461),
    .X(_00228_));
 sky130_fd_sc_hd__mux2_1 _27984_ (.A0(_00224_),
    .A1(_00225_),
    .S(net460),
    .X(_00226_));
 sky130_fd_sc_hd__mux2_1 _27985_ (.A0(_00171_),
    .A1(_00175_),
    .S(net461),
    .X(_00225_));
 sky130_fd_sc_hd__mux2_1 _27986_ (.A0(_00168_),
    .A1(_00170_),
    .S(net461),
    .X(_00224_));
 sky130_fd_sc_hd__mux2_1 _27987_ (.A0(_00164_),
    .A1(_00167_),
    .S(net461),
    .X(_00222_));
 sky130_fd_sc_hd__mux2_1 _27988_ (.A0(_00211_),
    .A1(_00219_),
    .S(net459),
    .X(_00220_));
 sky130_fd_sc_hd__mux2_1 _27989_ (.A0(_00214_),
    .A1(_00218_),
    .S(net222),
    .X(_00219_));
 sky130_fd_sc_hd__mux2_1 _27990_ (.A0(_00215_),
    .A1(_00217_),
    .S(net461),
    .X(_00218_));
 sky130_fd_sc_hd__mux2_1 _27991_ (.A0(net330),
    .A1(_00216_),
    .S(net200),
    .X(_00217_));
 sky130_fd_sc_hd__mux2_1 _27992_ (.A0(net327),
    .A1(net329),
    .S(net200),
    .X(_00215_));
 sky130_fd_sc_hd__mux2_1 _27993_ (.A0(_00212_),
    .A1(_00213_),
    .S(net461),
    .X(_00214_));
 sky130_fd_sc_hd__mux2_1 _27994_ (.A0(net325),
    .A1(net326),
    .S(net200),
    .X(_00213_));
 sky130_fd_sc_hd__mux2_1 _27995_ (.A0(net323),
    .A1(net324),
    .S(net200),
    .X(_00212_));
 sky130_fd_sc_hd__mux2_1 _27996_ (.A0(_00207_),
    .A1(_00210_),
    .S(net222),
    .X(_00211_));
 sky130_fd_sc_hd__mux2_1 _27997_ (.A0(_00208_),
    .A1(_00209_),
    .S(net461),
    .X(_00210_));
 sky130_fd_sc_hd__mux2_1 _27998_ (.A0(net321),
    .A1(net322),
    .S(net200),
    .X(_00209_));
 sky130_fd_sc_hd__mux2_1 _27999_ (.A0(net319),
    .A1(net320),
    .S(net200),
    .X(_00208_));
 sky130_fd_sc_hd__mux2_1 _28000_ (.A0(_00205_),
    .A1(_00206_),
    .S(net461),
    .X(_00207_));
 sky130_fd_sc_hd__mux2_1 _28001_ (.A0(net316),
    .A1(net318),
    .S(net200),
    .X(_00206_));
 sky130_fd_sc_hd__mux2_1 _28002_ (.A0(net314),
    .A1(net315),
    .S(net200),
    .X(_00205_));
 sky130_fd_sc_hd__mux2_1 _28003_ (.A0(_00199_),
    .A1(_00202_),
    .S(net222),
    .X(_00203_));
 sky130_fd_sc_hd__mux2_1 _28004_ (.A0(_00200_),
    .A1(_00201_),
    .S(net461),
    .X(_00202_));
 sky130_fd_sc_hd__mux2_1 _28005_ (.A0(net312),
    .A1(net313),
    .S(net200),
    .X(_00201_));
 sky130_fd_sc_hd__mux2_1 _28006_ (.A0(net310),
    .A1(net311),
    .S(net200),
    .X(_00200_));
 sky130_fd_sc_hd__mux2_1 _28007_ (.A0(_00197_),
    .A1(_00198_),
    .S(net461),
    .X(_00199_));
 sky130_fd_sc_hd__mux2_1 _28008_ (.A0(net308),
    .A1(net309),
    .S(net200),
    .X(_00198_));
 sky130_fd_sc_hd__mux2_1 _28009_ (.A0(net337),
    .A1(net307),
    .S(net200),
    .X(_00197_));
 sky130_fd_sc_hd__mux2_1 _28010_ (.A0(_00193_),
    .A1(_00194_),
    .S(net461),
    .X(_00195_));
 sky130_fd_sc_hd__mux2_1 _28011_ (.A0(net335),
    .A1(net336),
    .S(net200),
    .X(_00194_));
 sky130_fd_sc_hd__mux2_1 _28012_ (.A0(net333),
    .A1(net334),
    .S(net200),
    .X(_00193_));
 sky130_fd_sc_hd__mux2_1 _28013_ (.A0(net331),
    .A1(net332),
    .S(net200),
    .X(_00191_));
 sky130_fd_sc_hd__mux2_1 _28014_ (.A0(_00181_),
    .A1(_00188_),
    .S(net459),
    .X(_00189_));
 sky130_fd_sc_hd__mux2_1 _28015_ (.A0(_00184_),
    .A1(_00187_),
    .S(net460),
    .X(_00188_));
 sky130_fd_sc_hd__mux2_1 _28016_ (.A0(_00185_),
    .A1(_00186_),
    .S(net461),
    .X(_00187_));
 sky130_fd_sc_hd__mux2_1 _28017_ (.A0(net329),
    .A1(net330),
    .S(net462),
    .X(_00186_));
 sky130_fd_sc_hd__mux2_1 _28018_ (.A0(net326),
    .A1(net327),
    .S(net462),
    .X(_00185_));
 sky130_fd_sc_hd__mux2_1 _28019_ (.A0(_00182_),
    .A1(_00183_),
    .S(net461),
    .X(_00184_));
 sky130_fd_sc_hd__mux2_1 _28020_ (.A0(net324),
    .A1(net325),
    .S(net462),
    .X(_00183_));
 sky130_fd_sc_hd__mux2_1 _28021_ (.A0(net322),
    .A1(net323),
    .S(net462),
    .X(_00182_));
 sky130_fd_sc_hd__mux2_1 _28022_ (.A0(_00177_),
    .A1(_00180_),
    .S(net460),
    .X(_00181_));
 sky130_fd_sc_hd__mux2_1 _28023_ (.A0(_00178_),
    .A1(_00179_),
    .S(net461),
    .X(_00180_));
 sky130_fd_sc_hd__mux2_1 _28024_ (.A0(net320),
    .A1(net321),
    .S(net462),
    .X(_00179_));
 sky130_fd_sc_hd__mux2_1 _28025_ (.A0(net318),
    .A1(net319),
    .S(net462),
    .X(_00178_));
 sky130_fd_sc_hd__mux2_1 _28026_ (.A0(_00175_),
    .A1(_00176_),
    .S(net461),
    .X(_00177_));
 sky130_fd_sc_hd__mux2_1 _28027_ (.A0(net315),
    .A1(net316),
    .S(net462),
    .X(_00176_));
 sky130_fd_sc_hd__mux2_1 _28028_ (.A0(net313),
    .A1(net314),
    .S(net462),
    .X(_00175_));
 sky130_fd_sc_hd__mux2_1 _28029_ (.A0(_00169_),
    .A1(_00172_),
    .S(net460),
    .X(_00173_));
 sky130_fd_sc_hd__mux2_1 _28030_ (.A0(_00170_),
    .A1(_00171_),
    .S(net461),
    .X(_00172_));
 sky130_fd_sc_hd__mux2_1 _28031_ (.A0(net311),
    .A1(net312),
    .S(net462),
    .X(_00171_));
 sky130_fd_sc_hd__mux2_1 _28032_ (.A0(net309),
    .A1(net310),
    .S(net462),
    .X(_00170_));
 sky130_fd_sc_hd__mux2_1 _28033_ (.A0(_00167_),
    .A1(_00168_),
    .S(net461),
    .X(_00169_));
 sky130_fd_sc_hd__mux2_1 _28034_ (.A0(net307),
    .A1(net308),
    .S(net462),
    .X(_00168_));
 sky130_fd_sc_hd__mux2_1 _28035_ (.A0(net336),
    .A1(net337),
    .S(net462),
    .X(_00167_));
 sky130_fd_sc_hd__mux2_1 _28036_ (.A0(_00163_),
    .A1(_00164_),
    .S(net461),
    .X(_00165_));
 sky130_fd_sc_hd__mux2_1 _28037_ (.A0(net334),
    .A1(net335),
    .S(net462),
    .X(_00164_));
 sky130_fd_sc_hd__mux2_1 _28038_ (.A0(net332),
    .A1(net333),
    .S(net462),
    .X(_00163_));
 sky130_fd_sc_hd__mux2_1 _28039_ (.A0(net328),
    .A1(net331),
    .S(net462),
    .X(_00161_));
 sky130_fd_sc_hd__mux2_1 _28040_ (.A0(net327),
    .A1(net326),
    .S(net200),
    .X(_00148_));
 sky130_fd_sc_hd__mux2_1 _28041_ (.A0(net326),
    .A1(net325),
    .S(net462),
    .X(_00144_));
 sky130_fd_sc_hd__mux2_1 _28042_ (.A0(_00140_),
    .A1(_00132_),
    .S(net461),
    .X(_00141_));
 sky130_fd_sc_hd__mux2_1 _28043_ (.A0(net325),
    .A1(net324),
    .S(net200),
    .X(_00140_));
 sky130_fd_sc_hd__mux2_1 _28044_ (.A0(_00136_),
    .A1(_00128_),
    .S(net461),
    .X(_00137_));
 sky130_fd_sc_hd__mux2_1 _28045_ (.A0(net324),
    .A1(net323),
    .S(net462),
    .X(_00136_));
 sky130_fd_sc_hd__mux2_1 _28046_ (.A0(_00132_),
    .A1(_00123_),
    .S(net461),
    .X(_00133_));
 sky130_fd_sc_hd__mux2_1 _28047_ (.A0(net323),
    .A1(net322),
    .S(net200),
    .X(_00132_));
 sky130_fd_sc_hd__mux2_1 _28048_ (.A0(_00128_),
    .A1(_00117_),
    .S(net461),
    .X(_00129_));
 sky130_fd_sc_hd__mux2_1 _28049_ (.A0(net322),
    .A1(net321),
    .S(net462),
    .X(_00128_));
 sky130_fd_sc_hd__mux2_1 _28050_ (.A0(_00098_),
    .A1(_00100_),
    .S(net222),
    .X(_00126_));
 sky130_fd_sc_hd__mux2_1 _28051_ (.A0(_00124_),
    .A1(_00097_),
    .S(net222),
    .X(_00125_));
 sky130_fd_sc_hd__mux2_1 _28052_ (.A0(_00123_),
    .A1(_00111_),
    .S(net461),
    .X(_00124_));
 sky130_fd_sc_hd__mux2_1 _28053_ (.A0(net321),
    .A1(net320),
    .S(net200),
    .X(_00123_));
 sky130_fd_sc_hd__mux2_1 _28054_ (.A0(_00101_),
    .A1(_00094_),
    .S(net222),
    .X(_00122_));
 sky130_fd_sc_hd__mux2_1 _28055_ (.A0(_00088_),
    .A1(_00090_),
    .S(net460),
    .X(_00120_));
 sky130_fd_sc_hd__mux2_1 _28056_ (.A0(_00118_),
    .A1(_00087_),
    .S(net460),
    .X(_00119_));
 sky130_fd_sc_hd__mux2_1 _28057_ (.A0(_00117_),
    .A1(_00105_),
    .S(net461),
    .X(_00118_));
 sky130_fd_sc_hd__mux2_1 _28058_ (.A0(net320),
    .A1(net319),
    .S(net462),
    .X(_00117_));
 sky130_fd_sc_hd__mux2_2 _28059_ (.A0(_00091_),
    .A1(_00084_),
    .S(net460),
    .X(_00116_));
 sky130_fd_sc_hd__mux2_1 _28060_ (.A0(_00074_),
    .A1(_00078_),
    .S(net222),
    .X(_00114_));
 sky130_fd_sc_hd__mux2_1 _28061_ (.A0(_00112_),
    .A1(_00071_),
    .S(net222),
    .X(_00113_));
 sky130_fd_sc_hd__mux2_1 _28062_ (.A0(_00111_),
    .A1(_00096_),
    .S(net461),
    .X(_00112_));
 sky130_fd_sc_hd__mux2_1 _28063_ (.A0(net319),
    .A1(net318),
    .S(net200),
    .X(_00111_));
 sky130_fd_sc_hd__mux2_1 _28064_ (.A0(_00081_),
    .A1(_00067_),
    .S(net222),
    .X(_00110_));
 sky130_fd_sc_hd__mux2_1 _28065_ (.A0(_00056_),
    .A1(_00060_),
    .S(net460),
    .X(_00108_));
 sky130_fd_sc_hd__mux2_1 _28066_ (.A0(_00106_),
    .A1(_00053_),
    .S(net460),
    .X(_00107_));
 sky130_fd_sc_hd__mux2_1 _28067_ (.A0(_00105_),
    .A1(_00086_),
    .S(net461),
    .X(_00106_));
 sky130_fd_sc_hd__mux2_1 _28068_ (.A0(net318),
    .A1(net316),
    .S(net462),
    .X(_00105_));
 sky130_fd_sc_hd__mux2_2 _28069_ (.A0(_00063_),
    .A1(_00049_),
    .S(net460),
    .X(_00104_));
 sky130_fd_sc_hd__mux2_1 _28070_ (.A0(_00100_),
    .A1(_00101_),
    .S(net222),
    .X(_00102_));
 sky130_fd_sc_hd__mux2_1 _28071_ (.A0(_00077_),
    .A1(_00079_),
    .S(net211),
    .X(_00101_));
 sky130_fd_sc_hd__mux2_1 _28072_ (.A0(_00073_),
    .A1(_00076_),
    .S(net211),
    .X(_00100_));
 sky130_fd_sc_hd__mux2_1 _28073_ (.A0(_00097_),
    .A1(_00098_),
    .S(net222),
    .X(_00099_));
 sky130_fd_sc_hd__mux2_1 _28074_ (.A0(_00070_),
    .A1(_00072_),
    .S(net461),
    .X(_00098_));
 sky130_fd_sc_hd__mux2_1 _28075_ (.A0(_00096_),
    .A1(_00069_),
    .S(net461),
    .X(_00097_));
 sky130_fd_sc_hd__mux2_1 _28076_ (.A0(net316),
    .A1(net315),
    .S(net462),
    .X(_00096_));
 sky130_fd_sc_hd__mux2_1 _28077_ (.A0(_00080_),
    .A1(_00066_),
    .S(net211),
    .X(_00094_));
 sky130_fd_sc_hd__mux2_1 _28078_ (.A0(_00090_),
    .A1(_00091_),
    .S(net460),
    .X(_00092_));
 sky130_fd_sc_hd__mux2_1 _28079_ (.A0(_00059_),
    .A1(_00061_),
    .S(net211),
    .X(_00091_));
 sky130_fd_sc_hd__mux2_1 _28080_ (.A0(_00055_),
    .A1(_00058_),
    .S(net211),
    .X(_00090_));
 sky130_fd_sc_hd__mux2_1 _28081_ (.A0(_00087_),
    .A1(_00088_),
    .S(net460),
    .X(_00089_));
 sky130_fd_sc_hd__mux2_1 _28082_ (.A0(_00052_),
    .A1(_00054_),
    .S(net211),
    .X(_00088_));
 sky130_fd_sc_hd__mux2_1 _28083_ (.A0(_00086_),
    .A1(_00051_),
    .S(net461),
    .X(_00087_));
 sky130_fd_sc_hd__mux2_1 _28084_ (.A0(net315),
    .A1(net314),
    .S(net462),
    .X(_00086_));
 sky130_fd_sc_hd__mux2_1 _28085_ (.A0(_00062_),
    .A1(_00048_),
    .S(net211),
    .X(_00084_));
 sky130_fd_sc_hd__mux2_1 _28086_ (.A0(_00078_),
    .A1(_00081_),
    .S(net222),
    .X(_00082_));
 sky130_fd_sc_hd__mux2_1 _28087_ (.A0(_00079_),
    .A1(_00080_),
    .S(net211),
    .X(_00081_));
 sky130_fd_sc_hd__mux2_1 _28088_ (.A0(net331),
    .A1(net328),
    .S(net200),
    .X(_00080_));
 sky130_fd_sc_hd__mux2_1 _28089_ (.A0(net333),
    .A1(net332),
    .S(net200),
    .X(_00079_));
 sky130_fd_sc_hd__mux2_1 _28090_ (.A0(_00076_),
    .A1(_00077_),
    .S(net211),
    .X(_00078_));
 sky130_fd_sc_hd__mux2_1 _28091_ (.A0(net335),
    .A1(net334),
    .S(net200),
    .X(_00077_));
 sky130_fd_sc_hd__mux2_1 _28092_ (.A0(net337),
    .A1(net336),
    .S(net200),
    .X(_00076_));
 sky130_fd_sc_hd__mux2_1 _28093_ (.A0(_00071_),
    .A1(_00074_),
    .S(net222),
    .X(_00075_));
 sky130_fd_sc_hd__mux2_1 _28094_ (.A0(_00072_),
    .A1(_00073_),
    .S(net211),
    .X(_00074_));
 sky130_fd_sc_hd__mux2_1 _28095_ (.A0(net308),
    .A1(net307),
    .S(net200),
    .X(_00073_));
 sky130_fd_sc_hd__mux2_1 _28096_ (.A0(net310),
    .A1(net309),
    .S(net200),
    .X(_00072_));
 sky130_fd_sc_hd__mux2_1 _28097_ (.A0(_00069_),
    .A1(_00070_),
    .S(net461),
    .X(_00071_));
 sky130_fd_sc_hd__mux2_1 _28098_ (.A0(net312),
    .A1(net311),
    .S(net200),
    .X(_00070_));
 sky130_fd_sc_hd__mux2_1 _28099_ (.A0(net314),
    .A1(net313),
    .S(net462),
    .X(_00069_));
 sky130_fd_sc_hd__mux2_1 _28100_ (.A0(net317),
    .A1(net306),
    .S(net200),
    .X(_00066_));
 sky130_fd_sc_hd__mux2_1 _28101_ (.A0(_00060_),
    .A1(_00063_),
    .S(net460),
    .X(_00064_));
 sky130_fd_sc_hd__mux2_1 _28102_ (.A0(_00061_),
    .A1(_00062_),
    .S(net211),
    .X(_00063_));
 sky130_fd_sc_hd__mux2_1 _28103_ (.A0(net328),
    .A1(net317),
    .S(net200),
    .X(_00062_));
 sky130_fd_sc_hd__mux2_1 _28104_ (.A0(net332),
    .A1(net331),
    .S(net462),
    .X(_00061_));
 sky130_fd_sc_hd__mux2_1 _28105_ (.A0(_00058_),
    .A1(_00059_),
    .S(net211),
    .X(_00060_));
 sky130_fd_sc_hd__mux2_1 _28106_ (.A0(net334),
    .A1(net333),
    .S(net462),
    .X(_00059_));
 sky130_fd_sc_hd__mux2_1 _28107_ (.A0(net336),
    .A1(net335),
    .S(net462),
    .X(_00058_));
 sky130_fd_sc_hd__mux2_1 _28108_ (.A0(_00053_),
    .A1(_00056_),
    .S(net460),
    .X(_00057_));
 sky130_fd_sc_hd__mux2_1 _28109_ (.A0(_00054_),
    .A1(_00055_),
    .S(net211),
    .X(_00056_));
 sky130_fd_sc_hd__mux2_1 _28110_ (.A0(net307),
    .A1(net337),
    .S(net462),
    .X(_00055_));
 sky130_fd_sc_hd__mux2_1 _28111_ (.A0(net309),
    .A1(net308),
    .S(net462),
    .X(_00054_));
 sky130_fd_sc_hd__mux2_1 _28112_ (.A0(_00051_),
    .A1(_00052_),
    .S(net211),
    .X(_00053_));
 sky130_fd_sc_hd__mux2_1 _28113_ (.A0(net311),
    .A1(net310),
    .S(net462),
    .X(_00052_));
 sky130_fd_sc_hd__mux2_1 _28114_ (.A0(net313),
    .A1(net312),
    .S(net462),
    .X(_00051_));
 sky130_fd_sc_hd__mux2_1 _28115_ (.A0(_02408_),
    .A1(net362),
    .S(instr_sub),
    .X(_02409_));
 sky130_fd_sc_hd__mux2_1 _28116_ (.A0(_02406_),
    .A1(_02405_),
    .S(instr_sub),
    .X(_02407_));
 sky130_fd_sc_hd__mux2_1 _28117_ (.A0(_02403_),
    .A1(_02402_),
    .S(instr_sub),
    .X(_02404_));
 sky130_fd_sc_hd__mux2_1 _28118_ (.A0(_02400_),
    .A1(_02399_),
    .S(instr_sub),
    .X(_02401_));
 sky130_fd_sc_hd__mux2_1 _28119_ (.A0(_02397_),
    .A1(_02396_),
    .S(instr_sub),
    .X(_02398_));
 sky130_fd_sc_hd__mux2_1 _28120_ (.A0(_02394_),
    .A1(_02393_),
    .S(instr_sub),
    .X(_02395_));
 sky130_fd_sc_hd__mux2_1 _28121_ (.A0(_02391_),
    .A1(_02390_),
    .S(instr_sub),
    .X(_02392_));
 sky130_fd_sc_hd__mux2_2 _28122_ (.A0(_02388_),
    .A1(_02387_),
    .S(instr_sub),
    .X(_02389_));
 sky130_fd_sc_hd__mux2_1 _28123_ (.A0(_02385_),
    .A1(_02384_),
    .S(instr_sub),
    .X(_02386_));
 sky130_fd_sc_hd__mux2_1 _28124_ (.A0(_02382_),
    .A1(_02381_),
    .S(instr_sub),
    .X(_02383_));
 sky130_fd_sc_hd__mux2_1 _28125_ (.A0(_02379_),
    .A1(_02378_),
    .S(instr_sub),
    .X(_02380_));
 sky130_fd_sc_hd__mux2_1 _28126_ (.A0(_02376_),
    .A1(_02375_),
    .S(instr_sub),
    .X(_02377_));
 sky130_fd_sc_hd__mux2_1 _28127_ (.A0(_02373_),
    .A1(_02372_),
    .S(instr_sub),
    .X(_02374_));
 sky130_fd_sc_hd__mux2_1 _28128_ (.A0(_02370_),
    .A1(_02369_),
    .S(instr_sub),
    .X(_02371_));
 sky130_fd_sc_hd__mux2_1 _28129_ (.A0(_02367_),
    .A1(_02366_),
    .S(instr_sub),
    .X(_02368_));
 sky130_fd_sc_hd__mux2_2 _28130_ (.A0(_02364_),
    .A1(_02363_),
    .S(instr_sub),
    .X(_02365_));
 sky130_fd_sc_hd__mux2_1 _28131_ (.A0(_02361_),
    .A1(_02360_),
    .S(instr_sub),
    .X(_02362_));
 sky130_fd_sc_hd__mux2_1 _28132_ (.A0(_02358_),
    .A1(_02357_),
    .S(instr_sub),
    .X(_02359_));
 sky130_fd_sc_hd__mux2_1 _28133_ (.A0(_02355_),
    .A1(_02354_),
    .S(instr_sub),
    .X(_02356_));
 sky130_fd_sc_hd__mux2_1 _28134_ (.A0(_02352_),
    .A1(_02351_),
    .S(instr_sub),
    .X(_02353_));
 sky130_fd_sc_hd__mux2_1 _28135_ (.A0(_02349_),
    .A1(_02348_),
    .S(instr_sub),
    .X(_02350_));
 sky130_fd_sc_hd__mux2_1 _28136_ (.A0(_02346_),
    .A1(_02345_),
    .S(instr_sub),
    .X(_02347_));
 sky130_fd_sc_hd__mux2_1 _28137_ (.A0(_02343_),
    .A1(_02342_),
    .S(instr_sub),
    .X(_02344_));
 sky130_fd_sc_hd__mux2_2 _28138_ (.A0(_02340_),
    .A1(_02339_),
    .S(instr_sub),
    .X(_02341_));
 sky130_fd_sc_hd__mux2_1 _28139_ (.A0(_02337_),
    .A1(_02336_),
    .S(instr_sub),
    .X(_02338_));
 sky130_fd_sc_hd__mux2_2 _28140_ (.A0(_02334_),
    .A1(_02333_),
    .S(instr_sub),
    .X(_02335_));
 sky130_fd_sc_hd__mux2_2 _28141_ (.A0(_02331_),
    .A1(_02330_),
    .S(instr_sub),
    .X(_02332_));
 sky130_fd_sc_hd__mux2_1 _28142_ (.A0(_02328_),
    .A1(_02327_),
    .S(instr_sub),
    .X(_02329_));
 sky130_fd_sc_hd__mux2_1 _28143_ (.A0(_02325_),
    .A1(_02324_),
    .S(instr_sub),
    .X(_02326_));
 sky130_fd_sc_hd__mux2_1 _28144_ (.A0(_02322_),
    .A1(_02321_),
    .S(instr_sub),
    .X(_02323_));
 sky130_fd_sc_hd__mux2_1 _28145_ (.A0(_02319_),
    .A1(_02318_),
    .S(instr_sub),
    .X(_02320_));
 sky130_fd_sc_hd__mux2_1 _28146_ (.A0(_02313_),
    .A1(_02314_),
    .S(_00306_),
    .X(_02315_));
 sky130_fd_sc_hd__mux2_1 _28147_ (.A0(_02311_),
    .A1(_02315_),
    .S(_00303_),
    .X(_02316_));
 sky130_fd_sc_hd__mux2_1 _28148_ (.A0(_02311_),
    .A1(_02312_),
    .S(_00305_),
    .X(_02313_));
 sky130_fd_sc_hd__mux2_1 _28149_ (.A0(_02307_),
    .A1(_02308_),
    .S(\irq_state[1] ),
    .X(_02309_));
 sky130_fd_sc_hd__mux2_1 _28150_ (.A0(_02309_),
    .A1(_02307_),
    .S(_02217_),
    .X(_02310_));
 sky130_fd_sc_hd__mux2_1 _28151_ (.A0(_02302_),
    .A1(\irq_pending[0] ),
    .S(_01208_),
    .X(_02303_));
 sky130_fd_sc_hd__mux2_1 _28152_ (.A0(\reg_out[0] ),
    .A1(\alu_out_q[0] ),
    .S(latched_stalu),
    .X(_02070_));
 sky130_fd_sc_hd__mux2_1 _28153_ (.A0(_02063_),
    .A1(_00343_),
    .S(is_beq_bne_blt_bge_bltu_bgeu),
    .X(_02064_));
 sky130_fd_sc_hd__mux2_1 _28154_ (.A0(_02056_),
    .A1(_02055_),
    .S(net426),
    .X(_02057_));
 sky130_fd_sc_hd__mux2_1 _28155_ (.A0(_02058_),
    .A1(_02057_),
    .S(_01717_),
    .X(_02059_));
 sky130_fd_sc_hd__mux2_1 _28156_ (.A0(\pcpi_mul.rd[31] ),
    .A1(\pcpi_mul.rd[63] ),
    .S(\pcpi_mul.shift_out ),
    .X(_02054_));
 sky130_fd_sc_hd__mux2_2 _28157_ (.A0(_01908_),
    .A1(_02052_),
    .S(net455),
    .X(_02053_));
 sky130_fd_sc_hd__mux2_1 _28158_ (.A0(_02047_),
    .A1(_02046_),
    .S(net426),
    .X(_02048_));
 sky130_fd_sc_hd__mux2_1 _28159_ (.A0(_02049_),
    .A1(_02048_),
    .S(_01717_),
    .X(_02050_));
 sky130_fd_sc_hd__mux2_1 _28160_ (.A0(\pcpi_mul.rd[30] ),
    .A1(\pcpi_mul.rd[62] ),
    .S(\pcpi_mul.shift_out ),
    .X(_02045_));
 sky130_fd_sc_hd__mux2_2 _28161_ (.A0(_01908_),
    .A1(_02043_),
    .S(net455),
    .X(_02044_));
 sky130_fd_sc_hd__mux2_2 _28162_ (.A0(_02038_),
    .A1(_02037_),
    .S(net426),
    .X(_02039_));
 sky130_fd_sc_hd__mux2_2 _28163_ (.A0(_02040_),
    .A1(_02039_),
    .S(net429),
    .X(_02041_));
 sky130_fd_sc_hd__mux2_1 _28164_ (.A0(\pcpi_mul.rd[29] ),
    .A1(\pcpi_mul.rd[61] ),
    .S(\pcpi_mul.shift_out ),
    .X(_02036_));
 sky130_fd_sc_hd__mux2_2 _28165_ (.A0(_01908_),
    .A1(_02034_),
    .S(net455),
    .X(_02035_));
 sky130_fd_sc_hd__mux2_2 _28166_ (.A0(_02029_),
    .A1(_02028_),
    .S(net426),
    .X(_02030_));
 sky130_fd_sc_hd__mux2_1 _28167_ (.A0(_02031_),
    .A1(_02030_),
    .S(net429),
    .X(_02032_));
 sky130_fd_sc_hd__mux2_1 _28168_ (.A0(\pcpi_mul.rd[28] ),
    .A1(\pcpi_mul.rd[60] ),
    .S(\pcpi_mul.shift_out ),
    .X(_02027_));
 sky130_fd_sc_hd__mux2_2 _28169_ (.A0(_01908_),
    .A1(_02025_),
    .S(net455),
    .X(_02026_));
 sky130_fd_sc_hd__mux2_2 _28170_ (.A0(_02020_),
    .A1(_02019_),
    .S(net426),
    .X(_02021_));
 sky130_fd_sc_hd__mux2_4 _28171_ (.A0(_02022_),
    .A1(_02021_),
    .S(net429),
    .X(_02023_));
 sky130_fd_sc_hd__mux2_2 _28172_ (.A0(\pcpi_mul.rd[27] ),
    .A1(\pcpi_mul.rd[59] ),
    .S(\pcpi_mul.shift_out ),
    .X(_02018_));
 sky130_fd_sc_hd__mux2_2 _28173_ (.A0(_01908_),
    .A1(_02016_),
    .S(net455),
    .X(_02017_));
 sky130_fd_sc_hd__mux2_1 _28174_ (.A0(_02011_),
    .A1(_02010_),
    .S(net426),
    .X(_02012_));
 sky130_fd_sc_hd__mux2_2 _28175_ (.A0(_02013_),
    .A1(_02012_),
    .S(_01717_),
    .X(_02014_));
 sky130_fd_sc_hd__mux2_1 _28176_ (.A0(\pcpi_mul.rd[26] ),
    .A1(\pcpi_mul.rd[58] ),
    .S(\pcpi_mul.shift_out ),
    .X(_02009_));
 sky130_fd_sc_hd__mux2_2 _28177_ (.A0(_01908_),
    .A1(_02007_),
    .S(net455),
    .X(_02008_));
 sky130_fd_sc_hd__mux2_2 _28178_ (.A0(_02002_),
    .A1(_02001_),
    .S(_01714_),
    .X(_02003_));
 sky130_fd_sc_hd__mux2_4 _28179_ (.A0(_02004_),
    .A1(_02003_),
    .S(net429),
    .X(_02005_));
 sky130_fd_sc_hd__mux2_2 _28180_ (.A0(\pcpi_mul.rd[25] ),
    .A1(\pcpi_mul.rd[57] ),
    .S(\pcpi_mul.shift_out ),
    .X(_02000_));
 sky130_fd_sc_hd__mux2_2 _28181_ (.A0(_01908_),
    .A1(_01998_),
    .S(net455),
    .X(_01999_));
 sky130_fd_sc_hd__mux2_2 _28182_ (.A0(_01993_),
    .A1(_01992_),
    .S(_01714_),
    .X(_01994_));
 sky130_fd_sc_hd__mux2_2 _28183_ (.A0(_01995_),
    .A1(_01994_),
    .S(_01717_),
    .X(_01996_));
 sky130_fd_sc_hd__mux2_1 _28184_ (.A0(\pcpi_mul.rd[24] ),
    .A1(\pcpi_mul.rd[56] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01991_));
 sky130_fd_sc_hd__mux2_1 _28185_ (.A0(_01908_),
    .A1(_01989_),
    .S(net455),
    .X(_01990_));
 sky130_fd_sc_hd__mux2_2 _28186_ (.A0(_01984_),
    .A1(_01983_),
    .S(_01714_),
    .X(_01985_));
 sky130_fd_sc_hd__mux2_2 _28187_ (.A0(_01986_),
    .A1(_01985_),
    .S(_01717_),
    .X(_01987_));
 sky130_fd_sc_hd__mux2_1 _28188_ (.A0(\pcpi_mul.rd[23] ),
    .A1(\pcpi_mul.rd[55] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01982_));
 sky130_fd_sc_hd__mux2_1 _28189_ (.A0(_01908_),
    .A1(_01980_),
    .S(net455),
    .X(_01981_));
 sky130_fd_sc_hd__mux2_2 _28190_ (.A0(_01975_),
    .A1(_01974_),
    .S(_01714_),
    .X(_01976_));
 sky130_fd_sc_hd__mux2_2 _28191_ (.A0(_01977_),
    .A1(_01976_),
    .S(_01717_),
    .X(_01978_));
 sky130_fd_sc_hd__mux2_1 _28192_ (.A0(\pcpi_mul.rd[22] ),
    .A1(\pcpi_mul.rd[54] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01973_));
 sky130_fd_sc_hd__mux2_1 _28193_ (.A0(_01908_),
    .A1(_01971_),
    .S(net455),
    .X(_01972_));
 sky130_fd_sc_hd__mux2_2 _28194_ (.A0(_01966_),
    .A1(_01965_),
    .S(_01714_),
    .X(_01967_));
 sky130_fd_sc_hd__mux2_2 _28195_ (.A0(_01968_),
    .A1(_01967_),
    .S(_01717_),
    .X(_01969_));
 sky130_fd_sc_hd__mux2_1 _28196_ (.A0(\pcpi_mul.rd[21] ),
    .A1(\pcpi_mul.rd[53] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01964_));
 sky130_fd_sc_hd__mux2_1 _28197_ (.A0(_01908_),
    .A1(_01962_),
    .S(net455),
    .X(_01963_));
 sky130_fd_sc_hd__mux2_2 _28198_ (.A0(_01957_),
    .A1(_01956_),
    .S(_01714_),
    .X(_01958_));
 sky130_fd_sc_hd__mux2_2 _28199_ (.A0(_01959_),
    .A1(_01958_),
    .S(_01717_),
    .X(_01960_));
 sky130_fd_sc_hd__mux2_1 _28200_ (.A0(\pcpi_mul.rd[20] ),
    .A1(\pcpi_mul.rd[52] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01955_));
 sky130_fd_sc_hd__mux2_1 _28201_ (.A0(_01908_),
    .A1(_01953_),
    .S(net455),
    .X(_01954_));
 sky130_fd_sc_hd__mux2_2 _28202_ (.A0(_01948_),
    .A1(_01947_),
    .S(_01714_),
    .X(_01949_));
 sky130_fd_sc_hd__mux2_2 _28203_ (.A0(_01950_),
    .A1(_01949_),
    .S(_01717_),
    .X(_01951_));
 sky130_fd_sc_hd__mux2_1 _28204_ (.A0(\pcpi_mul.rd[19] ),
    .A1(\pcpi_mul.rd[51] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01946_));
 sky130_fd_sc_hd__mux2_1 _28205_ (.A0(_01908_),
    .A1(_01944_),
    .S(_01816_),
    .X(_01945_));
 sky130_fd_sc_hd__mux2_2 _28206_ (.A0(_01939_),
    .A1(_01938_),
    .S(_01714_),
    .X(_01940_));
 sky130_fd_sc_hd__mux2_2 _28207_ (.A0(_01941_),
    .A1(_01940_),
    .S(_01717_),
    .X(_01942_));
 sky130_fd_sc_hd__mux2_1 _28208_ (.A0(\pcpi_mul.rd[18] ),
    .A1(\pcpi_mul.rd[50] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01937_));
 sky130_fd_sc_hd__mux2_1 _28209_ (.A0(_01908_),
    .A1(_01935_),
    .S(_01816_),
    .X(_01936_));
 sky130_fd_sc_hd__mux2_2 _28210_ (.A0(_01930_),
    .A1(_01929_),
    .S(_01714_),
    .X(_01931_));
 sky130_fd_sc_hd__mux2_2 _28211_ (.A0(_01932_),
    .A1(_01931_),
    .S(net429),
    .X(_01933_));
 sky130_fd_sc_hd__mux2_1 _28212_ (.A0(\pcpi_mul.rd[17] ),
    .A1(\pcpi_mul.rd[49] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01928_));
 sky130_fd_sc_hd__mux2_1 _28213_ (.A0(_01908_),
    .A1(_01926_),
    .S(net455),
    .X(_01927_));
 sky130_fd_sc_hd__mux2_2 _28214_ (.A0(_01921_),
    .A1(_01920_),
    .S(_01714_),
    .X(_01922_));
 sky130_fd_sc_hd__mux2_2 _28215_ (.A0(_01923_),
    .A1(_01922_),
    .S(net430),
    .X(_01924_));
 sky130_fd_sc_hd__mux2_1 _28216_ (.A0(\pcpi_mul.rd[16] ),
    .A1(\pcpi_mul.rd[48] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01919_));
 sky130_fd_sc_hd__mux2_1 _28217_ (.A0(_01908_),
    .A1(_01917_),
    .S(_01816_),
    .X(_01918_));
 sky130_fd_sc_hd__mux2_2 _28218_ (.A0(_01912_),
    .A1(_01911_),
    .S(_01714_),
    .X(_01913_));
 sky130_fd_sc_hd__mux2_2 _28219_ (.A0(_01914_),
    .A1(_01913_),
    .S(net430),
    .X(_01915_));
 sky130_fd_sc_hd__mux2_1 _28220_ (.A0(\pcpi_mul.rd[15] ),
    .A1(\pcpi_mul.rd[47] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01910_));
 sky130_fd_sc_hd__mux2_2 _28221_ (.A0(_01908_),
    .A1(_01907_),
    .S(net455),
    .X(_01909_));
 sky130_fd_sc_hd__mux2_1 _28222_ (.A0(_01906_),
    .A1(_01904_),
    .S(net422),
    .X(_01907_));
 sky130_fd_sc_hd__mux2_1 _28223_ (.A0(net39),
    .A1(net57),
    .S(net317),
    .X(_01905_));
 sky130_fd_sc_hd__mux2_2 _28224_ (.A0(_01899_),
    .A1(_01898_),
    .S(_01714_),
    .X(_01900_));
 sky130_fd_sc_hd__mux2_2 _28225_ (.A0(_01901_),
    .A1(_01900_),
    .S(net430),
    .X(_01902_));
 sky130_fd_sc_hd__mux2_1 _28226_ (.A0(\pcpi_mul.rd[14] ),
    .A1(\pcpi_mul.rd[46] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01897_));
 sky130_fd_sc_hd__mux2_1 _28227_ (.A0(_01895_),
    .A1(_01894_),
    .S(net455),
    .X(_01896_));
 sky130_fd_sc_hd__mux2_1 _28228_ (.A0(_01893_),
    .A1(_01891_),
    .S(net422),
    .X(_01894_));
 sky130_fd_sc_hd__mux2_1 _28229_ (.A0(net38),
    .A1(net56),
    .S(net317),
    .X(_01892_));
 sky130_fd_sc_hd__mux2_2 _28230_ (.A0(_01886_),
    .A1(_01885_),
    .S(_01714_),
    .X(_01887_));
 sky130_fd_sc_hd__mux2_2 _28231_ (.A0(_01888_),
    .A1(_01887_),
    .S(net430),
    .X(_01889_));
 sky130_fd_sc_hd__mux2_1 _28232_ (.A0(\pcpi_mul.rd[13] ),
    .A1(\pcpi_mul.rd[45] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01884_));
 sky130_fd_sc_hd__mux2_1 _28233_ (.A0(_01882_),
    .A1(_01881_),
    .S(net455),
    .X(_01883_));
 sky130_fd_sc_hd__mux2_1 _28234_ (.A0(_01880_),
    .A1(_01878_),
    .S(net422),
    .X(_01881_));
 sky130_fd_sc_hd__mux2_1 _28235_ (.A0(net37),
    .A1(net54),
    .S(net317),
    .X(_01879_));
 sky130_fd_sc_hd__mux2_2 _28236_ (.A0(_01873_),
    .A1(_01872_),
    .S(_01714_),
    .X(_01874_));
 sky130_fd_sc_hd__mux2_2 _28237_ (.A0(_01875_),
    .A1(_01874_),
    .S(net430),
    .X(_01876_));
 sky130_fd_sc_hd__mux2_1 _28238_ (.A0(\pcpi_mul.rd[12] ),
    .A1(\pcpi_mul.rd[44] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01871_));
 sky130_fd_sc_hd__mux2_1 _28239_ (.A0(_01869_),
    .A1(_01868_),
    .S(net455),
    .X(_01870_));
 sky130_fd_sc_hd__mux2_1 _28240_ (.A0(_01867_),
    .A1(_01865_),
    .S(net422),
    .X(_01868_));
 sky130_fd_sc_hd__mux2_1 _28241_ (.A0(net36),
    .A1(net53),
    .S(net317),
    .X(_01866_));
 sky130_fd_sc_hd__mux2_2 _28242_ (.A0(_01860_),
    .A1(_01859_),
    .S(_01714_),
    .X(_01861_));
 sky130_fd_sc_hd__mux2_2 _28243_ (.A0(_01862_),
    .A1(_01861_),
    .S(net430),
    .X(_01863_));
 sky130_fd_sc_hd__mux2_2 _28244_ (.A0(\pcpi_mul.rd[11] ),
    .A1(\pcpi_mul.rd[43] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01858_));
 sky130_fd_sc_hd__mux2_1 _28245_ (.A0(_01856_),
    .A1(_01855_),
    .S(net455),
    .X(_01857_));
 sky130_fd_sc_hd__mux2_1 _28246_ (.A0(_01854_),
    .A1(_01852_),
    .S(net422),
    .X(_01855_));
 sky130_fd_sc_hd__mux2_1 _28247_ (.A0(net35),
    .A1(net52),
    .S(net317),
    .X(_01853_));
 sky130_fd_sc_hd__mux2_2 _28248_ (.A0(_01847_),
    .A1(_01846_),
    .S(_01714_),
    .X(_01848_));
 sky130_fd_sc_hd__mux2_2 _28249_ (.A0(_01849_),
    .A1(_01848_),
    .S(net430),
    .X(_01850_));
 sky130_fd_sc_hd__mux2_2 _28250_ (.A0(\pcpi_mul.rd[10] ),
    .A1(\pcpi_mul.rd[42] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01845_));
 sky130_fd_sc_hd__mux2_1 _28251_ (.A0(_01843_),
    .A1(_01842_),
    .S(net455),
    .X(_01844_));
 sky130_fd_sc_hd__mux2_1 _28252_ (.A0(_01841_),
    .A1(_01839_),
    .S(net422),
    .X(_01842_));
 sky130_fd_sc_hd__mux2_1 _28253_ (.A0(net34),
    .A1(net51),
    .S(net317),
    .X(_01840_));
 sky130_fd_sc_hd__mux2_1 _28254_ (.A0(_01834_),
    .A1(_01833_),
    .S(net426),
    .X(_01835_));
 sky130_fd_sc_hd__mux2_4 _28255_ (.A0(_01836_),
    .A1(_01835_),
    .S(net430),
    .X(_01837_));
 sky130_fd_sc_hd__mux2_2 _28256_ (.A0(\pcpi_mul.rd[9] ),
    .A1(\pcpi_mul.rd[41] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01832_));
 sky130_fd_sc_hd__mux2_2 _28257_ (.A0(_01830_),
    .A1(_01829_),
    .S(_01816_),
    .X(_01831_));
 sky130_fd_sc_hd__mux2_1 _28258_ (.A0(_01828_),
    .A1(_01826_),
    .S(net422),
    .X(_01829_));
 sky130_fd_sc_hd__mux2_1 _28259_ (.A0(net64),
    .A1(net50),
    .S(net317),
    .X(_01827_));
 sky130_fd_sc_hd__mux2_1 _28260_ (.A0(_01821_),
    .A1(_01820_),
    .S(net426),
    .X(_01822_));
 sky130_fd_sc_hd__mux2_2 _28261_ (.A0(_01823_),
    .A1(_01822_),
    .S(net430),
    .X(_01824_));
 sky130_fd_sc_hd__mux2_2 _28262_ (.A0(\pcpi_mul.rd[8] ),
    .A1(\pcpi_mul.rd[40] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01819_));
 sky130_fd_sc_hd__mux2_1 _28263_ (.A0(_01817_),
    .A1(_01815_),
    .S(net455),
    .X(_01818_));
 sky130_fd_sc_hd__mux2_1 _28264_ (.A0(_01814_),
    .A1(_01812_),
    .S(net422),
    .X(_01815_));
 sky130_fd_sc_hd__mux2_1 _28265_ (.A0(net63),
    .A1(net49),
    .S(net317),
    .X(_01813_));
 sky130_fd_sc_hd__mux2_1 _28266_ (.A0(_01807_),
    .A1(_01806_),
    .S(net426),
    .X(_01808_));
 sky130_fd_sc_hd__mux2_4 _28267_ (.A0(_01809_),
    .A1(_01808_),
    .S(net429),
    .X(_01810_));
 sky130_fd_sc_hd__mux2_2 _28268_ (.A0(\pcpi_mul.rd[7] ),
    .A1(\pcpi_mul.rd[39] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01805_));
 sky130_fd_sc_hd__mux2_4 _28269_ (.A0(_01803_),
    .A1(_01799_),
    .S(net422),
    .X(_01804_));
 sky130_fd_sc_hd__mux2_1 _28270_ (.A0(net62),
    .A1(net48),
    .S(net317),
    .X(_01802_));
 sky130_fd_sc_hd__mux2_1 _28271_ (.A0(_01800_),
    .A1(_01799_),
    .S(_00304_),
    .X(_01801_));
 sky130_fd_sc_hd__mux2_1 _28272_ (.A0(_01794_),
    .A1(_01793_),
    .S(net426),
    .X(_01795_));
 sky130_fd_sc_hd__mux2_2 _28273_ (.A0(_01796_),
    .A1(_01795_),
    .S(net429),
    .X(_01797_));
 sky130_fd_sc_hd__mux2_2 _28274_ (.A0(\pcpi_mul.rd[6] ),
    .A1(\pcpi_mul.rd[38] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01792_));
 sky130_fd_sc_hd__mux2_1 _28275_ (.A0(_01790_),
    .A1(_01786_),
    .S(net422),
    .X(_01791_));
 sky130_fd_sc_hd__mux2_1 _28276_ (.A0(net61),
    .A1(net47),
    .S(net317),
    .X(_01789_));
 sky130_fd_sc_hd__mux2_1 _28277_ (.A0(_01787_),
    .A1(_01786_),
    .S(_00304_),
    .X(_01788_));
 sky130_fd_sc_hd__mux2_1 _28278_ (.A0(_01781_),
    .A1(_01780_),
    .S(net426),
    .X(_01782_));
 sky130_fd_sc_hd__mux2_2 _28279_ (.A0(_01783_),
    .A1(_01782_),
    .S(net429),
    .X(_01784_));
 sky130_fd_sc_hd__mux2_2 _28280_ (.A0(\pcpi_mul.rd[5] ),
    .A1(\pcpi_mul.rd[37] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01779_));
 sky130_fd_sc_hd__mux2_2 _28281_ (.A0(_01777_),
    .A1(_01773_),
    .S(net422),
    .X(_01778_));
 sky130_fd_sc_hd__mux2_1 _28282_ (.A0(net60),
    .A1(net46),
    .S(net317),
    .X(_01776_));
 sky130_fd_sc_hd__mux2_1 _28283_ (.A0(_01774_),
    .A1(_01773_),
    .S(_00304_),
    .X(_01775_));
 sky130_fd_sc_hd__mux2_1 _28284_ (.A0(_01768_),
    .A1(_01767_),
    .S(net426),
    .X(_01769_));
 sky130_fd_sc_hd__mux2_2 _28285_ (.A0(_01770_),
    .A1(_01769_),
    .S(net429),
    .X(_01771_));
 sky130_fd_sc_hd__mux2_2 _28286_ (.A0(\pcpi_mul.rd[4] ),
    .A1(\pcpi_mul.rd[36] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01766_));
 sky130_fd_sc_hd__mux2_1 _28287_ (.A0(_01764_),
    .A1(_01760_),
    .S(net422),
    .X(_01765_));
 sky130_fd_sc_hd__mux2_1 _28288_ (.A0(net59),
    .A1(net464),
    .S(net317),
    .X(_01763_));
 sky130_fd_sc_hd__mux2_1 _28289_ (.A0(_01761_),
    .A1(_01760_),
    .S(_00304_),
    .X(_01762_));
 sky130_fd_sc_hd__mux2_1 _28290_ (.A0(_01755_),
    .A1(_01754_),
    .S(net426),
    .X(_01756_));
 sky130_fd_sc_hd__mux2_1 _28291_ (.A0(_01757_),
    .A1(_01756_),
    .S(net429),
    .X(_01758_));
 sky130_fd_sc_hd__mux2_4 _28292_ (.A0(\pcpi_mul.rd[3] ),
    .A1(\pcpi_mul.rd[35] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01753_));
 sky130_fd_sc_hd__mux2_1 _28293_ (.A0(_01751_),
    .A1(_01747_),
    .S(net422),
    .X(_01752_));
 sky130_fd_sc_hd__mux2_1 _28294_ (.A0(net58),
    .A1(net43),
    .S(net317),
    .X(_01750_));
 sky130_fd_sc_hd__mux2_1 _28295_ (.A0(_01748_),
    .A1(_01747_),
    .S(_00304_),
    .X(_01749_));
 sky130_fd_sc_hd__mux2_1 _28296_ (.A0(_01742_),
    .A1(_01741_),
    .S(net426),
    .X(_01743_));
 sky130_fd_sc_hd__mux2_1 _28297_ (.A0(_01744_),
    .A1(_01743_),
    .S(net429),
    .X(_01745_));
 sky130_fd_sc_hd__mux2_4 _28298_ (.A0(\pcpi_mul.rd[2] ),
    .A1(\pcpi_mul.rd[34] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01740_));
 sky130_fd_sc_hd__mux2_2 _28299_ (.A0(_01738_),
    .A1(_01734_),
    .S(net422),
    .X(_01739_));
 sky130_fd_sc_hd__mux2_1 _28300_ (.A0(net55),
    .A1(net42),
    .S(net317),
    .X(_01737_));
 sky130_fd_sc_hd__mux2_1 _28301_ (.A0(_01735_),
    .A1(_01734_),
    .S(_00304_),
    .X(_01736_));
 sky130_fd_sc_hd__mux2_1 _28302_ (.A0(_01729_),
    .A1(_01728_),
    .S(net426),
    .X(_01730_));
 sky130_fd_sc_hd__mux2_2 _28303_ (.A0(_01731_),
    .A1(_01730_),
    .S(net429),
    .X(_01732_));
 sky130_fd_sc_hd__mux2_2 _28304_ (.A0(\pcpi_mul.rd[1] ),
    .A1(\pcpi_mul.rd[33] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01727_));
 sky130_fd_sc_hd__mux2_1 _28305_ (.A0(_01725_),
    .A1(_01721_),
    .S(net422),
    .X(_01726_));
 sky130_fd_sc_hd__mux2_1 _28306_ (.A0(net44),
    .A1(net41),
    .S(net317),
    .X(_01724_));
 sky130_fd_sc_hd__mux2_1 _28307_ (.A0(_01722_),
    .A1(_01721_),
    .S(_00304_),
    .X(_01723_));
 sky130_fd_sc_hd__mux2_1 _28308_ (.A0(_01715_),
    .A1(_02559_),
    .S(net426),
    .X(_01716_));
 sky130_fd_sc_hd__mux2_2 _28309_ (.A0(_01718_),
    .A1(_01716_),
    .S(net429),
    .X(_01719_));
 sky130_fd_sc_hd__mux2_4 _28310_ (.A0(\pcpi_mul.rd[0] ),
    .A1(\pcpi_mul.rd[32] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01713_));
 sky130_fd_sc_hd__mux2_2 _28311_ (.A0(_01711_),
    .A1(_01707_),
    .S(net422),
    .X(_01712_));
 sky130_fd_sc_hd__mux2_1 _28312_ (.A0(net33),
    .A1(net40),
    .S(net317),
    .X(_01710_));
 sky130_fd_sc_hd__mux2_1 _28313_ (.A0(_01708_),
    .A1(_01707_),
    .S(_00304_),
    .X(_01709_));
 sky130_fd_sc_hd__mux2_1 _28314_ (.A0(_01701_),
    .A1(_01696_),
    .S(_00311_),
    .X(_01702_));
 sky130_fd_sc_hd__mux2_1 _28315_ (.A0(_01702_),
    .A1(_01696_),
    .S(\pcpi_mul.active[1] ),
    .X(_01703_));
 sky130_fd_sc_hd__mux2_1 _28316_ (.A0(_01696_),
    .A1(_01703_),
    .S(_00310_),
    .X(_01704_));
 sky130_fd_sc_hd__mux2_1 _28317_ (.A0(_01693_),
    .A1(net273),
    .S(_00316_),
    .X(_01694_));
 sky130_fd_sc_hd__mux2_1 _28318_ (.A0(_01690_),
    .A1(net272),
    .S(_00316_),
    .X(_01691_));
 sky130_fd_sc_hd__mux2_1 _28319_ (.A0(_01687_),
    .A1(net271),
    .S(_00316_),
    .X(_01688_));
 sky130_fd_sc_hd__mux2_1 _28320_ (.A0(_01684_),
    .A1(net270),
    .S(_00316_),
    .X(_01685_));
 sky130_fd_sc_hd__mux2_1 _28321_ (.A0(\reg_next_pc[31] ),
    .A1(_01554_),
    .S(latched_store),
    .X(_01555_));
 sky130_fd_sc_hd__mux2_1 _28322_ (.A0(\reg_out[31] ),
    .A1(\alu_out_q[31] ),
    .S(latched_stalu),
    .X(_01554_));
 sky130_fd_sc_hd__mux2_1 _28323_ (.A0(\reg_next_pc[30] ),
    .A1(_01551_),
    .S(latched_store),
    .X(_01552_));
 sky130_fd_sc_hd__mux2_1 _28324_ (.A0(\reg_out[30] ),
    .A1(\alu_out_q[30] ),
    .S(latched_stalu),
    .X(_01551_));
 sky130_fd_sc_hd__mux2_1 _28325_ (.A0(\reg_next_pc[29] ),
    .A1(_01548_),
    .S(latched_store),
    .X(_01549_));
 sky130_fd_sc_hd__mux2_1 _28326_ (.A0(\reg_out[29] ),
    .A1(\alu_out_q[29] ),
    .S(latched_stalu),
    .X(_01548_));
 sky130_fd_sc_hd__mux2_1 _28327_ (.A0(\reg_next_pc[28] ),
    .A1(_01545_),
    .S(latched_store),
    .X(_01546_));
 sky130_fd_sc_hd__mux2_1 _28328_ (.A0(\reg_out[28] ),
    .A1(\alu_out_q[28] ),
    .S(latched_stalu),
    .X(_01545_));
 sky130_fd_sc_hd__mux2_1 _28329_ (.A0(\reg_next_pc[27] ),
    .A1(_01542_),
    .S(latched_store),
    .X(_01543_));
 sky130_fd_sc_hd__mux2_1 _28330_ (.A0(\reg_out[27] ),
    .A1(\alu_out_q[27] ),
    .S(latched_stalu),
    .X(_01542_));
 sky130_fd_sc_hd__mux2_1 _28331_ (.A0(\reg_next_pc[26] ),
    .A1(_01539_),
    .S(latched_store),
    .X(_01540_));
 sky130_fd_sc_hd__mux2_1 _28332_ (.A0(\reg_out[26] ),
    .A1(\alu_out_q[26] ),
    .S(latched_stalu),
    .X(_01539_));
 sky130_fd_sc_hd__mux2_1 _28333_ (.A0(\reg_next_pc[25] ),
    .A1(_01536_),
    .S(latched_store),
    .X(_01537_));
 sky130_fd_sc_hd__mux2_1 _28334_ (.A0(\reg_out[25] ),
    .A1(\alu_out_q[25] ),
    .S(latched_stalu),
    .X(_01536_));
 sky130_fd_sc_hd__mux2_1 _28335_ (.A0(\reg_next_pc[24] ),
    .A1(_01533_),
    .S(latched_store),
    .X(_01534_));
 sky130_fd_sc_hd__mux2_1 _28336_ (.A0(\reg_out[24] ),
    .A1(\alu_out_q[24] ),
    .S(latched_stalu),
    .X(_01533_));
 sky130_fd_sc_hd__mux2_1 _28337_ (.A0(\reg_next_pc[23] ),
    .A1(_01530_),
    .S(latched_store),
    .X(_01531_));
 sky130_fd_sc_hd__mux2_1 _28338_ (.A0(\reg_out[23] ),
    .A1(\alu_out_q[23] ),
    .S(latched_stalu),
    .X(_01530_));
 sky130_fd_sc_hd__mux2_1 _28339_ (.A0(\reg_next_pc[22] ),
    .A1(_01527_),
    .S(latched_store),
    .X(_01528_));
 sky130_fd_sc_hd__mux2_1 _28340_ (.A0(\reg_out[22] ),
    .A1(\alu_out_q[22] ),
    .S(latched_stalu),
    .X(_01527_));
 sky130_fd_sc_hd__mux2_1 _28341_ (.A0(\reg_next_pc[21] ),
    .A1(_01524_),
    .S(latched_store),
    .X(_01525_));
 sky130_fd_sc_hd__mux2_1 _28342_ (.A0(\reg_out[21] ),
    .A1(\alu_out_q[21] ),
    .S(latched_stalu),
    .X(_01524_));
 sky130_fd_sc_hd__mux2_1 _28343_ (.A0(\reg_next_pc[20] ),
    .A1(_01521_),
    .S(latched_store),
    .X(_01522_));
 sky130_fd_sc_hd__mux2_1 _28344_ (.A0(\reg_out[20] ),
    .A1(\alu_out_q[20] ),
    .S(latched_stalu),
    .X(_01521_));
 sky130_fd_sc_hd__mux2_1 _28345_ (.A0(\reg_next_pc[19] ),
    .A1(_01518_),
    .S(latched_store),
    .X(_01519_));
 sky130_fd_sc_hd__mux2_1 _28346_ (.A0(\reg_out[19] ),
    .A1(\alu_out_q[19] ),
    .S(latched_stalu),
    .X(_01518_));
 sky130_fd_sc_hd__mux2_1 _28347_ (.A0(\reg_next_pc[18] ),
    .A1(_01515_),
    .S(latched_store),
    .X(_01516_));
 sky130_fd_sc_hd__mux2_1 _28348_ (.A0(\reg_out[18] ),
    .A1(\alu_out_q[18] ),
    .S(latched_stalu),
    .X(_01515_));
 sky130_fd_sc_hd__mux2_1 _28349_ (.A0(\reg_next_pc[17] ),
    .A1(_01512_),
    .S(latched_store),
    .X(_01513_));
 sky130_fd_sc_hd__mux2_1 _28350_ (.A0(\reg_out[17] ),
    .A1(\alu_out_q[17] ),
    .S(latched_stalu),
    .X(_01512_));
 sky130_fd_sc_hd__mux2_1 _28351_ (.A0(\reg_next_pc[16] ),
    .A1(_01509_),
    .S(latched_store),
    .X(_01510_));
 sky130_fd_sc_hd__mux2_1 _28352_ (.A0(\reg_out[16] ),
    .A1(\alu_out_q[16] ),
    .S(latched_stalu),
    .X(_01509_));
 sky130_fd_sc_hd__mux2_1 _28353_ (.A0(\reg_next_pc[15] ),
    .A1(_01506_),
    .S(latched_store),
    .X(_01507_));
 sky130_fd_sc_hd__mux2_1 _28354_ (.A0(\reg_out[15] ),
    .A1(\alu_out_q[15] ),
    .S(latched_stalu),
    .X(_01506_));
 sky130_fd_sc_hd__mux2_1 _28355_ (.A0(\reg_next_pc[14] ),
    .A1(_01503_),
    .S(latched_store),
    .X(_01504_));
 sky130_fd_sc_hd__mux2_1 _28356_ (.A0(\reg_out[14] ),
    .A1(\alu_out_q[14] ),
    .S(latched_stalu),
    .X(_01503_));
 sky130_fd_sc_hd__mux2_1 _28357_ (.A0(\reg_next_pc[13] ),
    .A1(_01500_),
    .S(latched_store),
    .X(_01501_));
 sky130_fd_sc_hd__mux2_1 _28358_ (.A0(\reg_out[13] ),
    .A1(\alu_out_q[13] ),
    .S(latched_stalu),
    .X(_01500_));
 sky130_fd_sc_hd__mux2_1 _28359_ (.A0(\reg_next_pc[12] ),
    .A1(_01497_),
    .S(latched_store),
    .X(_01498_));
 sky130_fd_sc_hd__mux2_1 _28360_ (.A0(\reg_out[12] ),
    .A1(\alu_out_q[12] ),
    .S(latched_stalu),
    .X(_01497_));
 sky130_fd_sc_hd__mux2_1 _28361_ (.A0(\reg_next_pc[11] ),
    .A1(_01494_),
    .S(latched_store),
    .X(_01495_));
 sky130_fd_sc_hd__mux2_1 _28362_ (.A0(\reg_out[11] ),
    .A1(\alu_out_q[11] ),
    .S(latched_stalu),
    .X(_01494_));
 sky130_fd_sc_hd__mux2_1 _28363_ (.A0(\reg_next_pc[10] ),
    .A1(_01491_),
    .S(latched_store),
    .X(_01492_));
 sky130_fd_sc_hd__mux2_1 _28364_ (.A0(\reg_out[10] ),
    .A1(\alu_out_q[10] ),
    .S(latched_stalu),
    .X(_01491_));
 sky130_fd_sc_hd__mux2_1 _28365_ (.A0(\reg_next_pc[9] ),
    .A1(_01488_),
    .S(latched_store),
    .X(_01489_));
 sky130_fd_sc_hd__mux2_1 _28366_ (.A0(\reg_out[9] ),
    .A1(\alu_out_q[9] ),
    .S(latched_stalu),
    .X(_01488_));
 sky130_fd_sc_hd__mux2_1 _28367_ (.A0(\reg_next_pc[8] ),
    .A1(_01485_),
    .S(latched_store),
    .X(_01486_));
 sky130_fd_sc_hd__mux2_1 _28368_ (.A0(\reg_out[8] ),
    .A1(\alu_out_q[8] ),
    .S(latched_stalu),
    .X(_01485_));
 sky130_fd_sc_hd__mux2_1 _28369_ (.A0(\reg_next_pc[7] ),
    .A1(_01482_),
    .S(latched_store),
    .X(_01483_));
 sky130_fd_sc_hd__mux2_1 _28370_ (.A0(\reg_out[7] ),
    .A1(\alu_out_q[7] ),
    .S(latched_stalu),
    .X(_01482_));
 sky130_fd_sc_hd__mux2_1 _28371_ (.A0(\reg_next_pc[6] ),
    .A1(_01479_),
    .S(latched_store),
    .X(_01480_));
 sky130_fd_sc_hd__mux2_1 _28372_ (.A0(\reg_out[6] ),
    .A1(\alu_out_q[6] ),
    .S(latched_stalu),
    .X(_01479_));
 sky130_fd_sc_hd__mux2_1 _28373_ (.A0(\reg_next_pc[5] ),
    .A1(_01476_),
    .S(latched_store),
    .X(_01477_));
 sky130_fd_sc_hd__mux2_1 _28374_ (.A0(\reg_out[5] ),
    .A1(\alu_out_q[5] ),
    .S(latched_stalu),
    .X(_01476_));
 sky130_fd_sc_hd__mux2_1 _28375_ (.A0(_01474_),
    .A1(_01471_),
    .S(net425),
    .X(_01475_));
 sky130_fd_sc_hd__mux2_1 _28376_ (.A0(\reg_next_pc[4] ),
    .A1(_01472_),
    .S(latched_store),
    .X(_01473_));
 sky130_fd_sc_hd__mux2_1 _28377_ (.A0(\reg_out[4] ),
    .A1(\alu_out_q[4] ),
    .S(latched_stalu),
    .X(_01472_));
 sky130_fd_sc_hd__mux2_1 _28378_ (.A0(\reg_next_pc[3] ),
    .A1(_01468_),
    .S(latched_store),
    .X(_01469_));
 sky130_fd_sc_hd__mux2_1 _28379_ (.A0(\reg_out[3] ),
    .A1(\alu_out_q[3] ),
    .S(latched_stalu),
    .X(_01468_));
 sky130_fd_sc_hd__mux2_1 _28380_ (.A0(\reg_next_pc[1] ),
    .A1(_01465_),
    .S(latched_store),
    .X(_01466_));
 sky130_fd_sc_hd__mux2_2 _28381_ (.A0(\reg_out[1] ),
    .A1(\alu_out_q[1] ),
    .S(latched_stalu),
    .X(_01465_));
 sky130_fd_sc_hd__mux2_1 _28382_ (.A0(_01301_),
    .A1(\timer[31] ),
    .S(_01208_),
    .X(_01302_));
 sky130_fd_sc_hd__mux2_1 _28383_ (.A0(_01298_),
    .A1(\timer[30] ),
    .S(_01208_),
    .X(_01299_));
 sky130_fd_sc_hd__mux2_1 _28384_ (.A0(_01295_),
    .A1(\timer[29] ),
    .S(_01208_),
    .X(_01296_));
 sky130_fd_sc_hd__mux2_1 _28385_ (.A0(_01292_),
    .A1(\timer[28] ),
    .S(net409),
    .X(_01293_));
 sky130_fd_sc_hd__mux2_1 _28386_ (.A0(_01289_),
    .A1(\timer[27] ),
    .S(net409),
    .X(_01290_));
 sky130_fd_sc_hd__mux2_1 _28387_ (.A0(_01286_),
    .A1(\timer[26] ),
    .S(net409),
    .X(_01287_));
 sky130_fd_sc_hd__mux2_1 _28388_ (.A0(_01283_),
    .A1(\timer[25] ),
    .S(net409),
    .X(_01284_));
 sky130_fd_sc_hd__mux2_1 _28389_ (.A0(_01280_),
    .A1(\timer[24] ),
    .S(net409),
    .X(_01281_));
 sky130_fd_sc_hd__mux2_1 _28390_ (.A0(_01277_),
    .A1(\timer[23] ),
    .S(net409),
    .X(_01278_));
 sky130_fd_sc_hd__mux2_1 _28391_ (.A0(_01274_),
    .A1(\timer[22] ),
    .S(net409),
    .X(_01275_));
 sky130_fd_sc_hd__mux2_1 _28392_ (.A0(_01271_),
    .A1(\timer[21] ),
    .S(net409),
    .X(_01272_));
 sky130_fd_sc_hd__mux2_1 _28393_ (.A0(_01268_),
    .A1(\timer[20] ),
    .S(net409),
    .X(_01269_));
 sky130_fd_sc_hd__mux2_1 _28394_ (.A0(_01265_),
    .A1(\timer[19] ),
    .S(net409),
    .X(_01266_));
 sky130_fd_sc_hd__mux2_1 _28395_ (.A0(_01262_),
    .A1(\timer[18] ),
    .S(net409),
    .X(_01263_));
 sky130_fd_sc_hd__mux2_1 _28396_ (.A0(_01259_),
    .A1(\timer[17] ),
    .S(net409),
    .X(_01260_));
 sky130_fd_sc_hd__mux2_1 _28397_ (.A0(_01256_),
    .A1(\timer[16] ),
    .S(net409),
    .X(_01257_));
 sky130_fd_sc_hd__mux2_1 _28398_ (.A0(_01253_),
    .A1(\timer[15] ),
    .S(net409),
    .X(_01254_));
 sky130_fd_sc_hd__mux2_1 _28399_ (.A0(_01250_),
    .A1(\timer[14] ),
    .S(net409),
    .X(_01251_));
 sky130_fd_sc_hd__mux2_1 _28400_ (.A0(_01247_),
    .A1(\timer[13] ),
    .S(net409),
    .X(_01248_));
 sky130_fd_sc_hd__mux2_1 _28401_ (.A0(_01244_),
    .A1(\timer[12] ),
    .S(_01208_),
    .X(_01245_));
 sky130_fd_sc_hd__mux2_1 _28402_ (.A0(_01241_),
    .A1(\timer[11] ),
    .S(_01208_),
    .X(_01242_));
 sky130_fd_sc_hd__mux2_1 _28403_ (.A0(_01238_),
    .A1(\timer[10] ),
    .S(_01208_),
    .X(_01239_));
 sky130_fd_sc_hd__mux2_1 _28404_ (.A0(_01235_),
    .A1(\timer[9] ),
    .S(_01208_),
    .X(_01236_));
 sky130_fd_sc_hd__mux2_1 _28405_ (.A0(_01232_),
    .A1(\timer[8] ),
    .S(_01208_),
    .X(_01233_));
 sky130_fd_sc_hd__mux2_1 _28406_ (.A0(_01229_),
    .A1(\timer[7] ),
    .S(_01208_),
    .X(_01230_));
 sky130_fd_sc_hd__mux2_1 _28407_ (.A0(_01226_),
    .A1(\timer[6] ),
    .S(_01208_),
    .X(_01227_));
 sky130_fd_sc_hd__mux2_1 _28408_ (.A0(_01223_),
    .A1(\timer[5] ),
    .S(_01208_),
    .X(_01224_));
 sky130_fd_sc_hd__mux2_1 _28409_ (.A0(_01220_),
    .A1(\timer[4] ),
    .S(_01208_),
    .X(_01221_));
 sky130_fd_sc_hd__mux2_1 _28410_ (.A0(_01217_),
    .A1(\timer[3] ),
    .S(_01208_),
    .X(_01218_));
 sky130_fd_sc_hd__mux2_1 _28411_ (.A0(_01214_),
    .A1(\timer[2] ),
    .S(_01208_),
    .X(_01215_));
 sky130_fd_sc_hd__mux2_1 _28412_ (.A0(_01211_),
    .A1(\timer[1] ),
    .S(_01208_),
    .X(_01212_));
 sky130_fd_sc_hd__mux2_4 _28413_ (.A0(_01206_),
    .A1(_01201_),
    .S(_00368_),
    .X(_01207_));
 sky130_fd_sc_hd__mux2_2 _28414_ (.A0(_01179_),
    .A1(_01174_),
    .S(_00368_),
    .X(_01180_));
 sky130_fd_sc_hd__mux2_4 _28415_ (.A0(_01152_),
    .A1(_01147_),
    .S(_00368_),
    .X(_01153_));
 sky130_fd_sc_hd__mux2_2 _28416_ (.A0(_01125_),
    .A1(_01120_),
    .S(_00368_),
    .X(_01126_));
 sky130_fd_sc_hd__mux2_4 _28417_ (.A0(_01098_),
    .A1(_01093_),
    .S(_00368_),
    .X(_01099_));
 sky130_fd_sc_hd__mux2_4 _28418_ (.A0(_01071_),
    .A1(_01066_),
    .S(_00368_),
    .X(_01072_));
 sky130_fd_sc_hd__mux2_4 _28419_ (.A0(_01044_),
    .A1(_01039_),
    .S(_00368_),
    .X(_01045_));
 sky130_fd_sc_hd__mux2_2 _28420_ (.A0(_01017_),
    .A1(_01012_),
    .S(_00368_),
    .X(_01018_));
 sky130_fd_sc_hd__mux2_2 _28421_ (.A0(_00990_),
    .A1(_00985_),
    .S(net428),
    .X(_00991_));
 sky130_fd_sc_hd__mux2_2 _28422_ (.A0(_00963_),
    .A1(_00958_),
    .S(net428),
    .X(_00964_));
 sky130_fd_sc_hd__mux2_2 _28423_ (.A0(_00936_),
    .A1(_00931_),
    .S(net428),
    .X(_00937_));
 sky130_fd_sc_hd__mux2_2 _28424_ (.A0(_00909_),
    .A1(_00904_),
    .S(net428),
    .X(_00910_));
 sky130_fd_sc_hd__mux2_4 _28425_ (.A0(_00882_),
    .A1(_00877_),
    .S(net428),
    .X(_00883_));
 sky130_fd_sc_hd__mux2_2 _28426_ (.A0(_00855_),
    .A1(_00850_),
    .S(net428),
    .X(_00856_));
 sky130_fd_sc_hd__mux2_4 _28427_ (.A0(_00828_),
    .A1(_00823_),
    .S(net428),
    .X(_00829_));
 sky130_fd_sc_hd__mux2_4 _28428_ (.A0(_00801_),
    .A1(_00796_),
    .S(net428),
    .X(_00802_));
 sky130_fd_sc_hd__mux2_4 _28429_ (.A0(_00774_),
    .A1(_00769_),
    .S(net427),
    .X(_00775_));
 sky130_fd_sc_hd__mux2_4 _28430_ (.A0(_00747_),
    .A1(_00742_),
    .S(net427),
    .X(_00748_));
 sky130_fd_sc_hd__mux2_4 _28431_ (.A0(_00720_),
    .A1(_00715_),
    .S(net427),
    .X(_00721_));
 sky130_fd_sc_hd__mux2_4 _28432_ (.A0(_00693_),
    .A1(_00688_),
    .S(net427),
    .X(_00694_));
 sky130_fd_sc_hd__mux2_8 _28433_ (.A0(_00666_),
    .A1(_00661_),
    .S(net427),
    .X(_00667_));
 sky130_fd_sc_hd__mux2_4 _28434_ (.A0(_00639_),
    .A1(_00634_),
    .S(net427),
    .X(_00640_));
 sky130_fd_sc_hd__mux2_4 _28435_ (.A0(_00612_),
    .A1(_00607_),
    .S(net427),
    .X(_00613_));
 sky130_fd_sc_hd__mux2_8 _28436_ (.A0(_00585_),
    .A1(_00580_),
    .S(net427),
    .X(_00586_));
 sky130_fd_sc_hd__mux2_4 _28437_ (.A0(_00558_),
    .A1(_00553_),
    .S(net427),
    .X(_00559_));
 sky130_fd_sc_hd__mux2_4 _28438_ (.A0(_00531_),
    .A1(_00526_),
    .S(net427),
    .X(_00532_));
 sky130_fd_sc_hd__mux2_4 _28439_ (.A0(_00504_),
    .A1(_00499_),
    .S(net427),
    .X(_00505_));
 sky130_fd_sc_hd__mux2_4 _28440_ (.A0(_00477_),
    .A1(_00472_),
    .S(net427),
    .X(_00478_));
 sky130_fd_sc_hd__mux2_4 _28441_ (.A0(_00450_),
    .A1(_00445_),
    .S(net427),
    .X(_00451_));
 sky130_fd_sc_hd__mux2_4 _28442_ (.A0(_00423_),
    .A1(_00418_),
    .S(net427),
    .X(_00424_));
 sky130_fd_sc_hd__mux2_4 _28443_ (.A0(_00396_),
    .A1(_00391_),
    .S(net428),
    .X(_00397_));
 sky130_fd_sc_hd__mux2_2 _28444_ (.A0(_00369_),
    .A1(_00365_),
    .S(net428),
    .X(_00370_));
 sky130_fd_sc_hd__mux2_8 _28445_ (.A0(_00366_),
    .A1(_00367_),
    .S(\cpu_state[3] ),
    .X(_00368_));
 sky130_fd_sc_hd__mux2_2 _28446_ (.A0(\decoded_rs1[3] ),
    .A1(\decoded_imm_uj[3] ),
    .S(net463),
    .X(_00362_));
 sky130_fd_sc_hd__mux2_8 _28447_ (.A0(\decoded_rs1[2] ),
    .A1(\decoded_imm_uj[2] ),
    .S(net463),
    .X(_00360_));
 sky130_fd_sc_hd__mux2_8 _28448_ (.A0(\decoded_rs1[1] ),
    .A1(\decoded_imm_uj[1] ),
    .S(net463),
    .X(_00358_));
 sky130_fd_sc_hd__mux2_2 _28449_ (.A0(\decoded_rs1[0] ),
    .A1(\decoded_imm_uj[11] ),
    .S(net463),
    .X(_00357_));
 sky130_fd_sc_hd__mux2_1 _28450_ (.A0(_00349_),
    .A1(_00323_),
    .S(decoder_trigger),
    .X(_00350_));
 sky130_fd_sc_hd__mux2_1 _28451_ (.A0(_00350_),
    .A1(_00351_),
    .S(_00309_),
    .X(_00352_));
 sky130_fd_sc_hd__mux2_1 _28452_ (.A0(_00352_),
    .A1(_00349_),
    .S(_00308_),
    .X(_00353_));
 sky130_fd_sc_hd__mux2_1 _28453_ (.A0(_00355_),
    .A1(_00353_),
    .S(_00354_),
    .X(_00356_));
 sky130_fd_sc_hd__mux2_1 _28454_ (.A0(_00337_),
    .A1(_00344_),
    .S(is_beq_bne_blt_bge_bltu_bgeu),
    .X(_00345_));
 sky130_fd_sc_hd__mux2_1 _28455_ (.A0(_00345_),
    .A1(_00337_),
    .S(alu_wait),
    .X(_00346_));
 sky130_fd_sc_hd__mux2_8 _28456_ (.A0(_00342_),
    .A1(_00340_),
    .S(_00341_),
    .X(_00343_));
 sky130_fd_sc_hd__mux2_1 _28457_ (.A0(_00338_),
    .A1(_00337_),
    .S(_00296_),
    .X(_00339_));
 sky130_fd_sc_hd__mux2_1 _28458_ (.A0(\mem_rdata_q[12] ),
    .A1(_00334_),
    .S(\mem_rdata_q[13] ),
    .X(_00335_));
 sky130_fd_sc_hd__mux2_1 _28459_ (.A0(\cpu_state[1] ),
    .A1(_00302_),
    .S(\cpu_state[4] ),
    .X(_00333_));
 sky130_fd_sc_hd__mux2_1 _28460_ (.A0(_00322_),
    .A1(_00296_),
    .S(\cpu_state[6] ),
    .X(_00332_));
 sky130_fd_sc_hd__mux2_1 _28461_ (.A0(_00315_),
    .A1(alu_wait),
    .S(\cpu_state[4] ),
    .X(_00331_));
 sky130_fd_sc_hd__mux2_2 _28462_ (.A0(\mem_rdata_q[6] ),
    .A1(net61),
    .S(mem_xfer),
    .X(_00330_));
 sky130_fd_sc_hd__mux2_1 _28463_ (.A0(\mem_rdata_q[5] ),
    .A1(net60),
    .S(mem_xfer),
    .X(_00329_));
 sky130_fd_sc_hd__mux2_2 _28464_ (.A0(\mem_rdata_q[4] ),
    .A1(net59),
    .S(mem_xfer),
    .X(_00328_));
 sky130_fd_sc_hd__mux2_2 _28465_ (.A0(\mem_rdata_q[3] ),
    .A1(net58),
    .S(mem_xfer),
    .X(_00327_));
 sky130_fd_sc_hd__mux2_1 _28466_ (.A0(\mem_rdata_q[2] ),
    .A1(net55),
    .S(mem_xfer),
    .X(_00326_));
 sky130_fd_sc_hd__mux2_1 _28467_ (.A0(\mem_rdata_q[1] ),
    .A1(net44),
    .S(mem_xfer),
    .X(_00325_));
 sky130_fd_sc_hd__mux2_1 _28468_ (.A0(\mem_rdata_q[0] ),
    .A1(net33),
    .S(mem_xfer),
    .X(_00324_));
 sky130_fd_sc_hd__mux2_1 _28469_ (.A0(\cpu_state[1] ),
    .A1(instr_retirq),
    .S(\cpu_state[2] ),
    .X(_00321_));
 sky130_fd_sc_hd__mux2_1 _28470_ (.A0(_00319_),
    .A1(\cpu_state[5] ),
    .S(_00296_),
    .X(_00320_));
 sky130_fd_sc_hd__mux2_1 _28471_ (.A0(_00317_),
    .A1(\cpu_state[6] ),
    .S(_00296_),
    .X(_00318_));
 sky130_fd_sc_hd__mux2_1 _28472_ (.A0(_00313_),
    .A1(_00312_),
    .S(_00307_),
    .X(_00314_));
 sky130_fd_sc_hd__mux2_1 _28473_ (.A0(_00298_),
    .A1(_00299_),
    .S(_00289_),
    .X(_00300_));
 sky130_fd_sc_hd__mux2_1 _28474_ (.A0(\reg_next_pc[2] ),
    .A1(_00293_),
    .S(latched_store),
    .X(_00294_));
 sky130_fd_sc_hd__mux2_1 _28475_ (.A0(\reg_out[2] ),
    .A1(\alu_out_q[2] ),
    .S(latched_stalu),
    .X(_00293_));
 sky130_fd_sc_hd__mux2_1 _28476_ (.A0(_00126_),
    .A1(_00122_),
    .S(net459),
    .X(_02558_));
 sky130_fd_sc_hd__mux2_1 _28477_ (.A0(_00120_),
    .A1(_00116_),
    .S(net459),
    .X(_02557_));
 sky130_fd_sc_hd__mux2_1 _28478_ (.A0(_00114_),
    .A1(_00110_),
    .S(net459),
    .X(_02556_));
 sky130_fd_sc_hd__mux2_1 _28479_ (.A0(_00108_),
    .A1(_00104_),
    .S(net225),
    .X(_02555_));
 sky130_fd_sc_hd__mux2_1 _28480_ (.A0(_00102_),
    .A1(_00095_),
    .S(net225),
    .X(_02554_));
 sky130_fd_sc_hd__mux2_1 _28481_ (.A0(_00092_),
    .A1(_00085_),
    .S(net225),
    .X(_02553_));
 sky130_fd_sc_hd__mux2_1 _28482_ (.A0(_00082_),
    .A1(_00068_),
    .S(net225),
    .X(_02552_));
 sky130_fd_sc_hd__mux2_1 _28483_ (.A0(_00064_),
    .A1(_00050_),
    .S(net225),
    .X(_02551_));
 sky130_fd_sc_hd__mux2_1 _28484_ (.A0(_01694_),
    .A1(_01695_),
    .S(_00290_),
    .X(_02541_));
 sky130_fd_sc_hd__mux2_1 _28485_ (.A0(_01691_),
    .A1(_01692_),
    .S(_00290_),
    .X(_02540_));
 sky130_fd_sc_hd__mux2_1 _28486_ (.A0(_01688_),
    .A1(_01689_),
    .S(_00290_),
    .X(_02539_));
 sky130_fd_sc_hd__mux2_1 _28487_ (.A0(_01685_),
    .A1(_01686_),
    .S(_00290_),
    .X(_02538_));
 sky130_fd_sc_hd__mux2_1 _28488_ (.A0(_01679_),
    .A1(_01680_),
    .S(instr_jal),
    .X(_01681_));
 sky130_fd_sc_hd__mux2_1 _28489_ (.A0(_01682_),
    .A1(_02581_),
    .S(net411),
    .X(_02530_));
 sky130_fd_sc_hd__mux2_1 _28490_ (.A0(_01675_),
    .A1(_01676_),
    .S(instr_jal),
    .X(_01677_));
 sky130_fd_sc_hd__mux2_1 _28491_ (.A0(_01678_),
    .A1(_02580_),
    .S(net411),
    .X(_02529_));
 sky130_fd_sc_hd__mux2_1 _28492_ (.A0(_01671_),
    .A1(_01672_),
    .S(instr_jal),
    .X(_01673_));
 sky130_fd_sc_hd__mux2_1 _28493_ (.A0(_01674_),
    .A1(_02579_),
    .S(net411),
    .X(_02527_));
 sky130_fd_sc_hd__mux2_1 _28494_ (.A0(_01667_),
    .A1(_01668_),
    .S(instr_jal),
    .X(_01669_));
 sky130_fd_sc_hd__mux2_1 _28495_ (.A0(_01670_),
    .A1(_02578_),
    .S(net411),
    .X(_02526_));
 sky130_fd_sc_hd__mux2_1 _28496_ (.A0(_01663_),
    .A1(_01664_),
    .S(instr_jal),
    .X(_01665_));
 sky130_fd_sc_hd__mux2_1 _28497_ (.A0(_01666_),
    .A1(_02577_),
    .S(net411),
    .X(_02525_));
 sky130_fd_sc_hd__mux2_1 _28498_ (.A0(_01659_),
    .A1(_01660_),
    .S(instr_jal),
    .X(_01661_));
 sky130_fd_sc_hd__mux2_1 _28499_ (.A0(_01662_),
    .A1(_02576_),
    .S(net411),
    .X(_02524_));
 sky130_fd_sc_hd__mux2_1 _28500_ (.A0(_01655_),
    .A1(_01656_),
    .S(instr_jal),
    .X(_01657_));
 sky130_fd_sc_hd__mux2_1 _28501_ (.A0(_01658_),
    .A1(_02575_),
    .S(net411),
    .X(_02523_));
 sky130_fd_sc_hd__mux2_1 _28502_ (.A0(_01651_),
    .A1(_01652_),
    .S(instr_jal),
    .X(_01653_));
 sky130_fd_sc_hd__mux2_1 _28503_ (.A0(_01654_),
    .A1(_02574_),
    .S(net411),
    .X(_02522_));
 sky130_fd_sc_hd__mux2_1 _28504_ (.A0(_01647_),
    .A1(_01648_),
    .S(instr_jal),
    .X(_01649_));
 sky130_fd_sc_hd__mux2_1 _28505_ (.A0(_01650_),
    .A1(_02573_),
    .S(net411),
    .X(_02521_));
 sky130_fd_sc_hd__mux2_1 _28506_ (.A0(_01643_),
    .A1(_01644_),
    .S(instr_jal),
    .X(_01645_));
 sky130_fd_sc_hd__mux2_1 _28507_ (.A0(_01646_),
    .A1(_02572_),
    .S(net411),
    .X(_02520_));
 sky130_fd_sc_hd__mux2_1 _28508_ (.A0(_01639_),
    .A1(_01640_),
    .S(instr_jal),
    .X(_01641_));
 sky130_fd_sc_hd__mux2_1 _28509_ (.A0(_01642_),
    .A1(_02570_),
    .S(net411),
    .X(_02519_));
 sky130_fd_sc_hd__mux2_1 _28510_ (.A0(_01635_),
    .A1(_01636_),
    .S(instr_jal),
    .X(_01637_));
 sky130_fd_sc_hd__mux2_1 _28511_ (.A0(_01638_),
    .A1(_02569_),
    .S(net411),
    .X(_02518_));
 sky130_fd_sc_hd__mux2_1 _28512_ (.A0(_01631_),
    .A1(_01632_),
    .S(instr_jal),
    .X(_01633_));
 sky130_fd_sc_hd__mux2_1 _28513_ (.A0(_01634_),
    .A1(_02568_),
    .S(net410),
    .X(_02516_));
 sky130_fd_sc_hd__mux2_1 _28514_ (.A0(_01627_),
    .A1(_01628_),
    .S(instr_jal),
    .X(_01629_));
 sky130_fd_sc_hd__mux2_1 _28515_ (.A0(_01630_),
    .A1(_02567_),
    .S(net410),
    .X(_02515_));
 sky130_fd_sc_hd__mux2_1 _28516_ (.A0(_01623_),
    .A1(_01624_),
    .S(instr_jal),
    .X(_01625_));
 sky130_fd_sc_hd__mux2_1 _28517_ (.A0(_01626_),
    .A1(_02566_),
    .S(net410),
    .X(_02514_));
 sky130_fd_sc_hd__mux2_1 _28518_ (.A0(_01619_),
    .A1(_01620_),
    .S(instr_jal),
    .X(_01621_));
 sky130_fd_sc_hd__mux2_1 _28519_ (.A0(_01622_),
    .A1(_02565_),
    .S(net410),
    .X(_02513_));
 sky130_fd_sc_hd__mux2_1 _28520_ (.A0(_01615_),
    .A1(_01616_),
    .S(instr_jal),
    .X(_01617_));
 sky130_fd_sc_hd__mux2_1 _28521_ (.A0(_01618_),
    .A1(_02564_),
    .S(net410),
    .X(_02512_));
 sky130_fd_sc_hd__mux2_1 _28522_ (.A0(_01611_),
    .A1(_01612_),
    .S(instr_jal),
    .X(_01613_));
 sky130_fd_sc_hd__mux2_1 _28523_ (.A0(_01614_),
    .A1(_02563_),
    .S(net410),
    .X(_02511_));
 sky130_fd_sc_hd__mux2_1 _28524_ (.A0(_01607_),
    .A1(_01608_),
    .S(instr_jal),
    .X(_01609_));
 sky130_fd_sc_hd__mux2_1 _28525_ (.A0(_01610_),
    .A1(_02562_),
    .S(net410),
    .X(_02510_));
 sky130_fd_sc_hd__mux2_1 _28526_ (.A0(_01603_),
    .A1(_01604_),
    .S(instr_jal),
    .X(_01605_));
 sky130_fd_sc_hd__mux2_1 _28527_ (.A0(_01606_),
    .A1(_02561_),
    .S(net410),
    .X(_02509_));
 sky130_fd_sc_hd__mux2_1 _28528_ (.A0(_01599_),
    .A1(_01600_),
    .S(instr_jal),
    .X(_01601_));
 sky130_fd_sc_hd__mux2_1 _28529_ (.A0(_01602_),
    .A1(_02589_),
    .S(net410),
    .X(_02508_));
 sky130_fd_sc_hd__mux2_1 _28530_ (.A0(_01595_),
    .A1(_01596_),
    .S(instr_jal),
    .X(_01597_));
 sky130_fd_sc_hd__mux2_1 _28531_ (.A0(_01598_),
    .A1(_02588_),
    .S(net410),
    .X(_02507_));
 sky130_fd_sc_hd__mux2_1 _28532_ (.A0(_01591_),
    .A1(_01592_),
    .S(instr_jal),
    .X(_01593_));
 sky130_fd_sc_hd__mux2_1 _28533_ (.A0(_01594_),
    .A1(_02587_),
    .S(net410),
    .X(_02537_));
 sky130_fd_sc_hd__mux2_1 _28534_ (.A0(_01587_),
    .A1(_01588_),
    .S(instr_jal),
    .X(_01589_));
 sky130_fd_sc_hd__mux2_1 _28535_ (.A0(_01590_),
    .A1(_02586_),
    .S(net410),
    .X(_02536_));
 sky130_fd_sc_hd__mux2_1 _28536_ (.A0(_01583_),
    .A1(_01584_),
    .S(instr_jal),
    .X(_01585_));
 sky130_fd_sc_hd__mux2_1 _28537_ (.A0(_01586_),
    .A1(_02585_),
    .S(net410),
    .X(_02535_));
 sky130_fd_sc_hd__mux2_1 _28538_ (.A0(_01579_),
    .A1(_01580_),
    .S(instr_jal),
    .X(_01581_));
 sky130_fd_sc_hd__mux2_1 _28539_ (.A0(_01582_),
    .A1(_02584_),
    .S(net410),
    .X(_02534_));
 sky130_fd_sc_hd__mux2_1 _28540_ (.A0(_01575_),
    .A1(_01576_),
    .S(instr_jal),
    .X(_01577_));
 sky130_fd_sc_hd__mux2_1 _28541_ (.A0(_01578_),
    .A1(_02583_),
    .S(net410),
    .X(_02533_));
 sky130_fd_sc_hd__mux2_1 _28542_ (.A0(_01571_),
    .A1(_01572_),
    .S(instr_jal),
    .X(_01573_));
 sky130_fd_sc_hd__mux2_1 _28543_ (.A0(_01574_),
    .A1(_02582_),
    .S(net410),
    .X(_02532_));
 sky130_fd_sc_hd__mux2_1 _28544_ (.A0(_01567_),
    .A1(_01568_),
    .S(instr_jal),
    .X(_01569_));
 sky130_fd_sc_hd__mux2_1 _28545_ (.A0(_01570_),
    .A1(_02571_),
    .S(_00308_),
    .X(_02531_));
 sky130_fd_sc_hd__mux2_1 _28546_ (.A0(_01561_),
    .A1(_01562_),
    .S(instr_jal),
    .X(_01563_));
 sky130_fd_sc_hd__mux2_1 _28547_ (.A0(_02560_),
    .A1(_01563_),
    .S(decoder_trigger),
    .X(_01564_));
 sky130_fd_sc_hd__mux2_1 _28548_ (.A0(_01564_),
    .A1(_01565_),
    .S(_00309_),
    .X(_01566_));
 sky130_fd_sc_hd__mux2_1 _28549_ (.A0(_01566_),
    .A1(_02560_),
    .S(_00308_),
    .X(_02528_));
 sky130_fd_sc_hd__mux2_1 _28550_ (.A0(_02590_),
    .A1(_01557_),
    .S(instr_jal),
    .X(_01558_));
 sky130_fd_sc_hd__mux2_1 _28551_ (.A0(_02590_),
    .A1(_01558_),
    .S(decoder_trigger),
    .X(_01559_));
 sky130_fd_sc_hd__mux2_1 _28552_ (.A0(_01559_),
    .A1(_02590_),
    .S(_00309_),
    .X(_01560_));
 sky130_fd_sc_hd__mux2_1 _28553_ (.A0(_01560_),
    .A1(_02590_),
    .S(_00308_),
    .X(_02517_));
 sky130_fd_sc_hd__mux2_1 _28554_ (.A0(\cpuregs_rs1[31] ),
    .A1(_01462_),
    .S(is_lui_auipc_jal),
    .X(_01463_));
 sky130_fd_sc_hd__mux2_1 _28555_ (.A0(_01464_),
    .A1(_01463_),
    .S(net424),
    .X(_02499_));
 sky130_fd_sc_hd__mux2_2 _28556_ (.A0(\cpuregs_rs1[30] ),
    .A1(_01459_),
    .S(is_lui_auipc_jal),
    .X(_01460_));
 sky130_fd_sc_hd__mux2_1 _28557_ (.A0(_01461_),
    .A1(_01460_),
    .S(net424),
    .X(_02498_));
 sky130_fd_sc_hd__mux2_2 _28558_ (.A0(\cpuregs_rs1[29] ),
    .A1(_01456_),
    .S(is_lui_auipc_jal),
    .X(_01457_));
 sky130_fd_sc_hd__mux2_1 _28559_ (.A0(_01458_),
    .A1(_01457_),
    .S(net424),
    .X(_02496_));
 sky130_fd_sc_hd__mux2_2 _28560_ (.A0(\cpuregs_rs1[28] ),
    .A1(_01453_),
    .S(is_lui_auipc_jal),
    .X(_01454_));
 sky130_fd_sc_hd__mux2_1 _28561_ (.A0(_01455_),
    .A1(_01454_),
    .S(net424),
    .X(_02495_));
 sky130_fd_sc_hd__mux2_2 _28562_ (.A0(\cpuregs_rs1[27] ),
    .A1(_01450_),
    .S(is_lui_auipc_jal),
    .X(_01451_));
 sky130_fd_sc_hd__mux2_1 _28563_ (.A0(_01452_),
    .A1(_01451_),
    .S(net423),
    .X(_02494_));
 sky130_fd_sc_hd__mux2_2 _28564_ (.A0(\cpuregs_rs1[26] ),
    .A1(_01447_),
    .S(is_lui_auipc_jal),
    .X(_01448_));
 sky130_fd_sc_hd__mux2_1 _28565_ (.A0(_01449_),
    .A1(_01448_),
    .S(net423),
    .X(_02493_));
 sky130_fd_sc_hd__mux2_2 _28566_ (.A0(\cpuregs_rs1[25] ),
    .A1(_01444_),
    .S(is_lui_auipc_jal),
    .X(_01445_));
 sky130_fd_sc_hd__mux2_1 _28567_ (.A0(_01446_),
    .A1(_01445_),
    .S(net423),
    .X(_02492_));
 sky130_fd_sc_hd__mux2_1 _28568_ (.A0(\cpuregs_rs1[24] ),
    .A1(_01441_),
    .S(is_lui_auipc_jal),
    .X(_01442_));
 sky130_fd_sc_hd__mux2_1 _28569_ (.A0(_01443_),
    .A1(_01442_),
    .S(net423),
    .X(_02491_));
 sky130_fd_sc_hd__mux2_1 _28570_ (.A0(\cpuregs_rs1[23] ),
    .A1(_01438_),
    .S(is_lui_auipc_jal),
    .X(_01439_));
 sky130_fd_sc_hd__mux2_1 _28571_ (.A0(_01440_),
    .A1(_01439_),
    .S(net423),
    .X(_02490_));
 sky130_fd_sc_hd__mux2_1 _28572_ (.A0(\cpuregs_rs1[22] ),
    .A1(_01435_),
    .S(is_lui_auipc_jal),
    .X(_01436_));
 sky130_fd_sc_hd__mux2_1 _28573_ (.A0(_01437_),
    .A1(_01436_),
    .S(net423),
    .X(_02489_));
 sky130_fd_sc_hd__mux2_1 _28574_ (.A0(\cpuregs_rs1[21] ),
    .A1(_01432_),
    .S(is_lui_auipc_jal),
    .X(_01433_));
 sky130_fd_sc_hd__mux2_1 _28575_ (.A0(_01434_),
    .A1(_01433_),
    .S(net423),
    .X(_02488_));
 sky130_fd_sc_hd__mux2_1 _28576_ (.A0(\cpuregs_rs1[20] ),
    .A1(_01429_),
    .S(is_lui_auipc_jal),
    .X(_01430_));
 sky130_fd_sc_hd__mux2_1 _28577_ (.A0(_01431_),
    .A1(_01430_),
    .S(net423),
    .X(_02487_));
 sky130_fd_sc_hd__mux2_1 _28578_ (.A0(\cpuregs_rs1[19] ),
    .A1(_01426_),
    .S(is_lui_auipc_jal),
    .X(_01427_));
 sky130_fd_sc_hd__mux2_1 _28579_ (.A0(_01428_),
    .A1(_01427_),
    .S(net423),
    .X(_02485_));
 sky130_fd_sc_hd__mux2_1 _28580_ (.A0(\cpuregs_rs1[18] ),
    .A1(_01423_),
    .S(is_lui_auipc_jal),
    .X(_01424_));
 sky130_fd_sc_hd__mux2_1 _28581_ (.A0(_01425_),
    .A1(_01424_),
    .S(net423),
    .X(_02484_));
 sky130_fd_sc_hd__mux2_1 _28582_ (.A0(\cpuregs_rs1[17] ),
    .A1(_01420_),
    .S(is_lui_auipc_jal),
    .X(_01421_));
 sky130_fd_sc_hd__mux2_1 _28583_ (.A0(_01422_),
    .A1(_01421_),
    .S(net423),
    .X(_02483_));
 sky130_fd_sc_hd__mux2_1 _28584_ (.A0(\cpuregs_rs1[16] ),
    .A1(_01417_),
    .S(is_lui_auipc_jal),
    .X(_01418_));
 sky130_fd_sc_hd__mux2_1 _28585_ (.A0(_01419_),
    .A1(_01418_),
    .S(net423),
    .X(_02482_));
 sky130_fd_sc_hd__mux2_1 _28586_ (.A0(\cpuregs_rs1[15] ),
    .A1(_01414_),
    .S(is_lui_auipc_jal),
    .X(_01415_));
 sky130_fd_sc_hd__mux2_1 _28587_ (.A0(_01416_),
    .A1(_01415_),
    .S(net423),
    .X(_02481_));
 sky130_fd_sc_hd__mux2_1 _28588_ (.A0(\cpuregs_rs1[14] ),
    .A1(_01411_),
    .S(is_lui_auipc_jal),
    .X(_01412_));
 sky130_fd_sc_hd__mux2_1 _28589_ (.A0(_01413_),
    .A1(_01412_),
    .S(net423),
    .X(_02480_));
 sky130_fd_sc_hd__mux2_1 _28590_ (.A0(\cpuregs_rs1[13] ),
    .A1(_01408_),
    .S(is_lui_auipc_jal),
    .X(_01409_));
 sky130_fd_sc_hd__mux2_1 _28591_ (.A0(_01410_),
    .A1(_01409_),
    .S(net423),
    .X(_02479_));
 sky130_fd_sc_hd__mux2_1 _28592_ (.A0(\cpuregs_rs1[12] ),
    .A1(_01405_),
    .S(is_lui_auipc_jal),
    .X(_01406_));
 sky130_fd_sc_hd__mux2_1 _28593_ (.A0(_01407_),
    .A1(_01406_),
    .S(net423),
    .X(_02478_));
 sky130_fd_sc_hd__mux2_1 _28594_ (.A0(\cpuregs_rs1[11] ),
    .A1(_01402_),
    .S(is_lui_auipc_jal),
    .X(_01403_));
 sky130_fd_sc_hd__mux2_1 _28595_ (.A0(_01404_),
    .A1(_01403_),
    .S(net423),
    .X(_02477_));
 sky130_fd_sc_hd__mux2_1 _28596_ (.A0(\cpuregs_rs1[10] ),
    .A1(_01399_),
    .S(is_lui_auipc_jal),
    .X(_01400_));
 sky130_fd_sc_hd__mux2_1 _28597_ (.A0(_01401_),
    .A1(_01400_),
    .S(net424),
    .X(_02476_));
 sky130_fd_sc_hd__mux2_1 _28598_ (.A0(\cpuregs_rs1[9] ),
    .A1(_01396_),
    .S(is_lui_auipc_jal),
    .X(_01397_));
 sky130_fd_sc_hd__mux2_1 _28599_ (.A0(_01398_),
    .A1(_01397_),
    .S(net424),
    .X(_02506_));
 sky130_fd_sc_hd__mux2_1 _28600_ (.A0(\cpuregs_rs1[8] ),
    .A1(_01393_),
    .S(is_lui_auipc_jal),
    .X(_01394_));
 sky130_fd_sc_hd__mux2_1 _28601_ (.A0(_01395_),
    .A1(_01394_),
    .S(net424),
    .X(_02505_));
 sky130_fd_sc_hd__mux2_1 _28602_ (.A0(\cpuregs_rs1[7] ),
    .A1(_01390_),
    .S(is_lui_auipc_jal),
    .X(_01391_));
 sky130_fd_sc_hd__mux2_1 _28603_ (.A0(_01392_),
    .A1(_01391_),
    .S(net424),
    .X(_02504_));
 sky130_fd_sc_hd__mux2_1 _28604_ (.A0(\cpuregs_rs1[6] ),
    .A1(_01387_),
    .S(is_lui_auipc_jal),
    .X(_01388_));
 sky130_fd_sc_hd__mux2_1 _28605_ (.A0(_01389_),
    .A1(_01388_),
    .S(net424),
    .X(_02503_));
 sky130_fd_sc_hd__mux2_1 _28606_ (.A0(\cpuregs_rs1[5] ),
    .A1(_01384_),
    .S(is_lui_auipc_jal),
    .X(_01385_));
 sky130_fd_sc_hd__mux2_1 _28607_ (.A0(_01386_),
    .A1(_01385_),
    .S(net424),
    .X(_02502_));
 sky130_fd_sc_hd__mux2_1 _28608_ (.A0(\cpuregs_rs1[4] ),
    .A1(_01381_),
    .S(is_lui_auipc_jal),
    .X(_01382_));
 sky130_fd_sc_hd__mux2_1 _28609_ (.A0(_01383_),
    .A1(_01382_),
    .S(net424),
    .X(_02501_));
 sky130_fd_sc_hd__mux2_1 _28610_ (.A0(\cpuregs_rs1[3] ),
    .A1(_01378_),
    .S(is_lui_auipc_jal),
    .X(_01379_));
 sky130_fd_sc_hd__mux2_1 _28611_ (.A0(_01380_),
    .A1(_01379_),
    .S(net424),
    .X(_02500_));
 sky130_fd_sc_hd__mux2_1 _28612_ (.A0(\cpuregs_rs1[2] ),
    .A1(_01375_),
    .S(is_lui_auipc_jal),
    .X(_01376_));
 sky130_fd_sc_hd__mux2_1 _28613_ (.A0(_01377_),
    .A1(_01376_),
    .S(net424),
    .X(_02497_));
 sky130_fd_sc_hd__mux2_1 _28614_ (.A0(\cpuregs_rs1[1] ),
    .A1(_01372_),
    .S(is_lui_auipc_jal),
    .X(_01373_));
 sky130_fd_sc_hd__mux2_1 _28615_ (.A0(_01374_),
    .A1(_01373_),
    .S(net424),
    .X(_02486_));
 sky130_fd_sc_hd__mux2_1 _28616_ (.A0(\cpuregs_rs1[0] ),
    .A1(_01369_),
    .S(is_lui_auipc_jal),
    .X(_01370_));
 sky130_fd_sc_hd__mux2_1 _28617_ (.A0(_01371_),
    .A1(_01370_),
    .S(_00297_),
    .X(_02475_));
 sky130_fd_sc_hd__mux2_1 _28618_ (.A0(_01367_),
    .A1(\decoded_imm[31] ),
    .S(net457),
    .X(_01368_));
 sky130_fd_sc_hd__mux2_1 _28619_ (.A0(_01368_),
    .A1(\cpuregs_rs1[31] ),
    .S(net463),
    .X(_02467_));
 sky130_fd_sc_hd__mux2_1 _28620_ (.A0(_01365_),
    .A1(\decoded_imm[30] ),
    .S(net457),
    .X(_01366_));
 sky130_fd_sc_hd__mux2_1 _28621_ (.A0(_01366_),
    .A1(\cpuregs_rs1[30] ),
    .S(net463),
    .X(_02466_));
 sky130_fd_sc_hd__mux2_1 _28622_ (.A0(_01363_),
    .A1(\decoded_imm[29] ),
    .S(net457),
    .X(_01364_));
 sky130_fd_sc_hd__mux2_2 _28623_ (.A0(_01364_),
    .A1(\cpuregs_rs1[29] ),
    .S(net463),
    .X(_02464_));
 sky130_fd_sc_hd__mux2_1 _28624_ (.A0(_01361_),
    .A1(\decoded_imm[28] ),
    .S(net457),
    .X(_01362_));
 sky130_fd_sc_hd__mux2_2 _28625_ (.A0(_01362_),
    .A1(\cpuregs_rs1[28] ),
    .S(net463),
    .X(_02463_));
 sky130_fd_sc_hd__mux2_1 _28626_ (.A0(_01359_),
    .A1(\decoded_imm[27] ),
    .S(net457),
    .X(_01360_));
 sky130_fd_sc_hd__mux2_2 _28627_ (.A0(_01360_),
    .A1(\cpuregs_rs1[27] ),
    .S(net463),
    .X(_02462_));
 sky130_fd_sc_hd__mux2_1 _28628_ (.A0(_01357_),
    .A1(\decoded_imm[26] ),
    .S(net457),
    .X(_01358_));
 sky130_fd_sc_hd__mux2_2 _28629_ (.A0(_01358_),
    .A1(\cpuregs_rs1[26] ),
    .S(net463),
    .X(_02461_));
 sky130_fd_sc_hd__mux2_1 _28630_ (.A0(_01355_),
    .A1(\decoded_imm[25] ),
    .S(net457),
    .X(_01356_));
 sky130_fd_sc_hd__mux2_2 _28631_ (.A0(_01356_),
    .A1(\cpuregs_rs1[25] ),
    .S(net463),
    .X(_02460_));
 sky130_fd_sc_hd__mux2_1 _28632_ (.A0(_01353_),
    .A1(\decoded_imm[24] ),
    .S(net457),
    .X(_01354_));
 sky130_fd_sc_hd__mux2_1 _28633_ (.A0(_01354_),
    .A1(\cpuregs_rs1[24] ),
    .S(net463),
    .X(_02459_));
 sky130_fd_sc_hd__mux2_1 _28634_ (.A0(_01351_),
    .A1(\decoded_imm[23] ),
    .S(net456),
    .X(_01352_));
 sky130_fd_sc_hd__mux2_1 _28635_ (.A0(_01352_),
    .A1(\cpuregs_rs1[23] ),
    .S(net463),
    .X(_02458_));
 sky130_fd_sc_hd__mux2_1 _28636_ (.A0(_01349_),
    .A1(\decoded_imm[22] ),
    .S(net456),
    .X(_01350_));
 sky130_fd_sc_hd__mux2_1 _28637_ (.A0(_01350_),
    .A1(\cpuregs_rs1[22] ),
    .S(net463),
    .X(_02457_));
 sky130_fd_sc_hd__mux2_1 _28638_ (.A0(_01347_),
    .A1(\decoded_imm[21] ),
    .S(net456),
    .X(_01348_));
 sky130_fd_sc_hd__mux2_1 _28639_ (.A0(_01348_),
    .A1(\cpuregs_rs1[21] ),
    .S(net463),
    .X(_02456_));
 sky130_fd_sc_hd__mux2_1 _28640_ (.A0(_01345_),
    .A1(\decoded_imm[20] ),
    .S(net456),
    .X(_01346_));
 sky130_fd_sc_hd__mux2_1 _28641_ (.A0(_01346_),
    .A1(\cpuregs_rs1[20] ),
    .S(net463),
    .X(_02455_));
 sky130_fd_sc_hd__mux2_1 _28642_ (.A0(_01343_),
    .A1(\decoded_imm[19] ),
    .S(net456),
    .X(_01344_));
 sky130_fd_sc_hd__mux2_1 _28643_ (.A0(_01344_),
    .A1(\cpuregs_rs1[19] ),
    .S(net463),
    .X(_02453_));
 sky130_fd_sc_hd__mux2_1 _28644_ (.A0(_01341_),
    .A1(\decoded_imm[18] ),
    .S(net456),
    .X(_01342_));
 sky130_fd_sc_hd__mux2_1 _28645_ (.A0(_01342_),
    .A1(\cpuregs_rs1[18] ),
    .S(net463),
    .X(_02452_));
 sky130_fd_sc_hd__mux2_1 _28646_ (.A0(_01339_),
    .A1(\decoded_imm[17] ),
    .S(net456),
    .X(_01340_));
 sky130_fd_sc_hd__mux2_1 _28647_ (.A0(_01340_),
    .A1(\cpuregs_rs1[17] ),
    .S(net463),
    .X(_02451_));
 sky130_fd_sc_hd__mux2_1 _28648_ (.A0(_01337_),
    .A1(\decoded_imm[16] ),
    .S(net456),
    .X(_01338_));
 sky130_fd_sc_hd__mux2_1 _28649_ (.A0(_01338_),
    .A1(\cpuregs_rs1[16] ),
    .S(net463),
    .X(_02450_));
 sky130_fd_sc_hd__mux2_1 _28650_ (.A0(_01335_),
    .A1(\decoded_imm[15] ),
    .S(net456),
    .X(_01336_));
 sky130_fd_sc_hd__mux2_1 _28651_ (.A0(_01336_),
    .A1(\cpuregs_rs1[15] ),
    .S(net463),
    .X(_02449_));
 sky130_fd_sc_hd__mux2_1 _28652_ (.A0(_01333_),
    .A1(\decoded_imm[14] ),
    .S(net456),
    .X(_01334_));
 sky130_fd_sc_hd__mux2_1 _28653_ (.A0(_01334_),
    .A1(\cpuregs_rs1[14] ),
    .S(net463),
    .X(_02448_));
 sky130_fd_sc_hd__mux2_1 _28654_ (.A0(_01331_),
    .A1(\decoded_imm[13] ),
    .S(net456),
    .X(_01332_));
 sky130_fd_sc_hd__mux2_1 _28655_ (.A0(_01332_),
    .A1(\cpuregs_rs1[13] ),
    .S(net463),
    .X(_02447_));
 sky130_fd_sc_hd__mux2_1 _28656_ (.A0(_01329_),
    .A1(\decoded_imm[12] ),
    .S(net456),
    .X(_01330_));
 sky130_fd_sc_hd__mux2_1 _28657_ (.A0(_01330_),
    .A1(\cpuregs_rs1[12] ),
    .S(net463),
    .X(_02446_));
 sky130_fd_sc_hd__mux2_1 _28658_ (.A0(_01327_),
    .A1(\decoded_imm[11] ),
    .S(net456),
    .X(_01328_));
 sky130_fd_sc_hd__mux2_1 _28659_ (.A0(_01328_),
    .A1(\cpuregs_rs1[11] ),
    .S(net463),
    .X(_02445_));
 sky130_fd_sc_hd__mux2_1 _28660_ (.A0(_01325_),
    .A1(\decoded_imm[10] ),
    .S(net456),
    .X(_01326_));
 sky130_fd_sc_hd__mux2_1 _28661_ (.A0(_01326_),
    .A1(\cpuregs_rs1[10] ),
    .S(net463),
    .X(_02444_));
 sky130_fd_sc_hd__mux2_1 _28662_ (.A0(_01323_),
    .A1(\decoded_imm[9] ),
    .S(net456),
    .X(_01324_));
 sky130_fd_sc_hd__mux2_1 _28663_ (.A0(_01324_),
    .A1(\cpuregs_rs1[9] ),
    .S(net463),
    .X(_02474_));
 sky130_fd_sc_hd__mux2_1 _28664_ (.A0(_01321_),
    .A1(\decoded_imm[8] ),
    .S(net456),
    .X(_01322_));
 sky130_fd_sc_hd__mux2_1 _28665_ (.A0(_01322_),
    .A1(\cpuregs_rs1[8] ),
    .S(net463),
    .X(_02473_));
 sky130_fd_sc_hd__mux2_1 _28666_ (.A0(_01319_),
    .A1(\decoded_imm[7] ),
    .S(net456),
    .X(_01320_));
 sky130_fd_sc_hd__mux2_1 _28667_ (.A0(_01320_),
    .A1(\cpuregs_rs1[7] ),
    .S(net463),
    .X(_02472_));
 sky130_fd_sc_hd__mux2_1 _28668_ (.A0(_01317_),
    .A1(\decoded_imm[6] ),
    .S(_01304_),
    .X(_01318_));
 sky130_fd_sc_hd__mux2_1 _28669_ (.A0(_01318_),
    .A1(\cpuregs_rs1[6] ),
    .S(net463),
    .X(_02471_));
 sky130_fd_sc_hd__mux2_1 _28670_ (.A0(_01315_),
    .A1(\decoded_imm[5] ),
    .S(_01304_),
    .X(_01316_));
 sky130_fd_sc_hd__mux2_1 _28671_ (.A0(_01316_),
    .A1(\cpuregs_rs1[5] ),
    .S(net463),
    .X(_02470_));
 sky130_fd_sc_hd__mux2_1 _28672_ (.A0(\decoded_imm[4] ),
    .A1(\decoded_imm_uj[4] ),
    .S(is_slli_srli_srai),
    .X(_01313_));
 sky130_fd_sc_hd__mux2_1 _28673_ (.A0(_01313_),
    .A1(\decoded_imm[4] ),
    .S(_01304_),
    .X(_01314_));
 sky130_fd_sc_hd__mux2_1 _28674_ (.A0(_01314_),
    .A1(\cpuregs_rs1[4] ),
    .S(net463),
    .X(_02469_));
 sky130_fd_sc_hd__mux2_1 _28675_ (.A0(\decoded_imm[3] ),
    .A1(\decoded_imm_uj[3] ),
    .S(is_slli_srli_srai),
    .X(_01311_));
 sky130_fd_sc_hd__mux2_1 _28676_ (.A0(_01311_),
    .A1(\decoded_imm[3] ),
    .S(_01304_),
    .X(_01312_));
 sky130_fd_sc_hd__mux2_1 _28677_ (.A0(_01312_),
    .A1(\cpuregs_rs1[3] ),
    .S(net463),
    .X(_02468_));
 sky130_fd_sc_hd__mux2_1 _28678_ (.A0(\decoded_imm[2] ),
    .A1(\decoded_imm_uj[2] ),
    .S(is_slli_srli_srai),
    .X(_01309_));
 sky130_fd_sc_hd__mux2_1 _28679_ (.A0(_01309_),
    .A1(\decoded_imm[2] ),
    .S(_01304_),
    .X(_01310_));
 sky130_fd_sc_hd__mux2_1 _28680_ (.A0(_01310_),
    .A1(\cpuregs_rs1[2] ),
    .S(net463),
    .X(_02465_));
 sky130_fd_sc_hd__mux2_1 _28681_ (.A0(\decoded_imm[1] ),
    .A1(\decoded_imm_uj[1] ),
    .S(is_slli_srli_srai),
    .X(_01307_));
 sky130_fd_sc_hd__mux2_1 _28682_ (.A0(_01307_),
    .A1(\decoded_imm[1] ),
    .S(_01304_),
    .X(_01308_));
 sky130_fd_sc_hd__mux2_1 _28683_ (.A0(_01308_),
    .A1(\cpuregs_rs1[1] ),
    .S(net463),
    .X(_02454_));
 sky130_fd_sc_hd__mux2_1 _28684_ (.A0(\decoded_imm[0] ),
    .A1(\decoded_imm_uj[11] ),
    .S(is_slli_srli_srai),
    .X(_01305_));
 sky130_fd_sc_hd__mux2_1 _28685_ (.A0(_01305_),
    .A1(\decoded_imm[0] ),
    .S(_01304_),
    .X(_01306_));
 sky130_fd_sc_hd__mux2_1 _28686_ (.A0(_01306_),
    .A1(\cpuregs_rs1[0] ),
    .S(net463),
    .X(_02443_));
 sky130_fd_sc_hd__mux2_1 _28687_ (.A0(_01302_),
    .A1(\cpuregs_rs1[31] ),
    .S(instr_timer),
    .X(_01303_));
 sky130_fd_sc_hd__mux2_1 _28688_ (.A0(_01302_),
    .A1(_01303_),
    .S(\cpu_state[2] ),
    .X(_02435_));
 sky130_fd_sc_hd__mux2_1 _28689_ (.A0(_01299_),
    .A1(\cpuregs_rs1[30] ),
    .S(instr_timer),
    .X(_01300_));
 sky130_fd_sc_hd__mux2_1 _28690_ (.A0(_01299_),
    .A1(_01300_),
    .S(\cpu_state[2] ),
    .X(_02434_));
 sky130_fd_sc_hd__mux2_1 _28691_ (.A0(_01296_),
    .A1(\cpuregs_rs1[29] ),
    .S(instr_timer),
    .X(_01297_));
 sky130_fd_sc_hd__mux2_1 _28692_ (.A0(_01296_),
    .A1(_01297_),
    .S(\cpu_state[2] ),
    .X(_02432_));
 sky130_fd_sc_hd__mux2_1 _28693_ (.A0(_01293_),
    .A1(\cpuregs_rs1[28] ),
    .S(instr_timer),
    .X(_01294_));
 sky130_fd_sc_hd__mux2_1 _28694_ (.A0(_01293_),
    .A1(_01294_),
    .S(\cpu_state[2] ),
    .X(_02431_));
 sky130_fd_sc_hd__mux2_1 _28695_ (.A0(_01290_),
    .A1(\cpuregs_rs1[27] ),
    .S(instr_timer),
    .X(_01291_));
 sky130_fd_sc_hd__mux2_1 _28696_ (.A0(_01290_),
    .A1(_01291_),
    .S(\cpu_state[2] ),
    .X(_02430_));
 sky130_fd_sc_hd__mux2_1 _28697_ (.A0(_01287_),
    .A1(\cpuregs_rs1[26] ),
    .S(instr_timer),
    .X(_01288_));
 sky130_fd_sc_hd__mux2_1 _28698_ (.A0(_01287_),
    .A1(_01288_),
    .S(\cpu_state[2] ),
    .X(_02429_));
 sky130_fd_sc_hd__mux2_1 _28699_ (.A0(_01284_),
    .A1(\cpuregs_rs1[25] ),
    .S(instr_timer),
    .X(_01285_));
 sky130_fd_sc_hd__mux2_1 _28700_ (.A0(_01284_),
    .A1(_01285_),
    .S(\cpu_state[2] ),
    .X(_02428_));
 sky130_fd_sc_hd__mux2_1 _28701_ (.A0(_01281_),
    .A1(\cpuregs_rs1[24] ),
    .S(instr_timer),
    .X(_01282_));
 sky130_fd_sc_hd__mux2_1 _28702_ (.A0(_01281_),
    .A1(_01282_),
    .S(\cpu_state[2] ),
    .X(_02427_));
 sky130_fd_sc_hd__mux2_1 _28703_ (.A0(_01278_),
    .A1(\cpuregs_rs1[23] ),
    .S(instr_timer),
    .X(_01279_));
 sky130_fd_sc_hd__mux2_1 _28704_ (.A0(_01278_),
    .A1(_01279_),
    .S(\cpu_state[2] ),
    .X(_02426_));
 sky130_fd_sc_hd__mux2_1 _28705_ (.A0(_01275_),
    .A1(\cpuregs_rs1[22] ),
    .S(instr_timer),
    .X(_01276_));
 sky130_fd_sc_hd__mux2_1 _28706_ (.A0(_01275_),
    .A1(_01276_),
    .S(\cpu_state[2] ),
    .X(_02425_));
 sky130_fd_sc_hd__mux2_1 _28707_ (.A0(_01272_),
    .A1(\cpuregs_rs1[21] ),
    .S(instr_timer),
    .X(_01273_));
 sky130_fd_sc_hd__mux2_1 _28708_ (.A0(_01272_),
    .A1(_01273_),
    .S(\cpu_state[2] ),
    .X(_02424_));
 sky130_fd_sc_hd__mux2_1 _28709_ (.A0(_01269_),
    .A1(\cpuregs_rs1[20] ),
    .S(instr_timer),
    .X(_01270_));
 sky130_fd_sc_hd__mux2_1 _28710_ (.A0(_01269_),
    .A1(_01270_),
    .S(\cpu_state[2] ),
    .X(_02423_));
 sky130_fd_sc_hd__mux2_1 _28711_ (.A0(_01266_),
    .A1(\cpuregs_rs1[19] ),
    .S(instr_timer),
    .X(_01267_));
 sky130_fd_sc_hd__mux2_1 _28712_ (.A0(_01266_),
    .A1(_01267_),
    .S(\cpu_state[2] ),
    .X(_02421_));
 sky130_fd_sc_hd__mux2_1 _28713_ (.A0(_01263_),
    .A1(\cpuregs_rs1[18] ),
    .S(instr_timer),
    .X(_01264_));
 sky130_fd_sc_hd__mux2_1 _28714_ (.A0(_01263_),
    .A1(_01264_),
    .S(\cpu_state[2] ),
    .X(_02420_));
 sky130_fd_sc_hd__mux2_1 _28715_ (.A0(_01260_),
    .A1(\cpuregs_rs1[17] ),
    .S(instr_timer),
    .X(_01261_));
 sky130_fd_sc_hd__mux2_1 _28716_ (.A0(_01260_),
    .A1(_01261_),
    .S(\cpu_state[2] ),
    .X(_02419_));
 sky130_fd_sc_hd__mux2_1 _28717_ (.A0(_01257_),
    .A1(\cpuregs_rs1[16] ),
    .S(instr_timer),
    .X(_01258_));
 sky130_fd_sc_hd__mux2_1 _28718_ (.A0(_01257_),
    .A1(_01258_),
    .S(\cpu_state[2] ),
    .X(_02418_));
 sky130_fd_sc_hd__mux2_1 _28719_ (.A0(_01254_),
    .A1(\cpuregs_rs1[15] ),
    .S(instr_timer),
    .X(_01255_));
 sky130_fd_sc_hd__mux2_1 _28720_ (.A0(_01254_),
    .A1(_01255_),
    .S(\cpu_state[2] ),
    .X(_02417_));
 sky130_fd_sc_hd__mux2_1 _28721_ (.A0(_01251_),
    .A1(\cpuregs_rs1[14] ),
    .S(instr_timer),
    .X(_01252_));
 sky130_fd_sc_hd__mux2_1 _28722_ (.A0(_01251_),
    .A1(_01252_),
    .S(\cpu_state[2] ),
    .X(_02416_));
 sky130_fd_sc_hd__mux2_1 _28723_ (.A0(_01248_),
    .A1(\cpuregs_rs1[13] ),
    .S(instr_timer),
    .X(_01249_));
 sky130_fd_sc_hd__mux2_1 _28724_ (.A0(_01248_),
    .A1(_01249_),
    .S(\cpu_state[2] ),
    .X(_02415_));
 sky130_fd_sc_hd__mux2_1 _28725_ (.A0(_01245_),
    .A1(\cpuregs_rs1[12] ),
    .S(instr_timer),
    .X(_01246_));
 sky130_fd_sc_hd__mux2_1 _28726_ (.A0(_01245_),
    .A1(_01246_),
    .S(\cpu_state[2] ),
    .X(_02414_));
 sky130_fd_sc_hd__mux2_1 _28727_ (.A0(_01242_),
    .A1(\cpuregs_rs1[11] ),
    .S(instr_timer),
    .X(_01243_));
 sky130_fd_sc_hd__mux2_1 _28728_ (.A0(_01242_),
    .A1(_01243_),
    .S(\cpu_state[2] ),
    .X(_02413_));
 sky130_fd_sc_hd__mux2_1 _28729_ (.A0(_01239_),
    .A1(\cpuregs_rs1[10] ),
    .S(instr_timer),
    .X(_01240_));
 sky130_fd_sc_hd__mux2_1 _28730_ (.A0(_01239_),
    .A1(_01240_),
    .S(\cpu_state[2] ),
    .X(_02412_));
 sky130_fd_sc_hd__mux2_1 _28731_ (.A0(_01236_),
    .A1(\cpuregs_rs1[9] ),
    .S(instr_timer),
    .X(_01237_));
 sky130_fd_sc_hd__mux2_1 _28732_ (.A0(_01236_),
    .A1(_01237_),
    .S(\cpu_state[2] ),
    .X(_02442_));
 sky130_fd_sc_hd__mux2_1 _28733_ (.A0(_01233_),
    .A1(\cpuregs_rs1[8] ),
    .S(instr_timer),
    .X(_01234_));
 sky130_fd_sc_hd__mux2_1 _28734_ (.A0(_01233_),
    .A1(_01234_),
    .S(\cpu_state[2] ),
    .X(_02441_));
 sky130_fd_sc_hd__mux2_1 _28735_ (.A0(_01230_),
    .A1(\cpuregs_rs1[7] ),
    .S(instr_timer),
    .X(_01231_));
 sky130_fd_sc_hd__mux2_1 _28736_ (.A0(_01230_),
    .A1(_01231_),
    .S(\cpu_state[2] ),
    .X(_02440_));
 sky130_fd_sc_hd__mux2_1 _28737_ (.A0(_01227_),
    .A1(\cpuregs_rs1[6] ),
    .S(instr_timer),
    .X(_01228_));
 sky130_fd_sc_hd__mux2_1 _28738_ (.A0(_01227_),
    .A1(_01228_),
    .S(\cpu_state[2] ),
    .X(_02439_));
 sky130_fd_sc_hd__mux2_1 _28739_ (.A0(_01224_),
    .A1(\cpuregs_rs1[5] ),
    .S(instr_timer),
    .X(_01225_));
 sky130_fd_sc_hd__mux2_1 _28740_ (.A0(_01224_),
    .A1(_01225_),
    .S(\cpu_state[2] ),
    .X(_02438_));
 sky130_fd_sc_hd__mux2_1 _28741_ (.A0(_01221_),
    .A1(\cpuregs_rs1[4] ),
    .S(instr_timer),
    .X(_01222_));
 sky130_fd_sc_hd__mux2_1 _28742_ (.A0(_01221_),
    .A1(_01222_),
    .S(\cpu_state[2] ),
    .X(_02437_));
 sky130_fd_sc_hd__mux2_1 _28743_ (.A0(_01218_),
    .A1(\cpuregs_rs1[3] ),
    .S(instr_timer),
    .X(_01219_));
 sky130_fd_sc_hd__mux2_1 _28744_ (.A0(_01218_),
    .A1(_01219_),
    .S(\cpu_state[2] ),
    .X(_02436_));
 sky130_fd_sc_hd__mux2_1 _28745_ (.A0(_01215_),
    .A1(\cpuregs_rs1[2] ),
    .S(instr_timer),
    .X(_01216_));
 sky130_fd_sc_hd__mux2_1 _28746_ (.A0(_01215_),
    .A1(_01216_),
    .S(\cpu_state[2] ),
    .X(_02433_));
 sky130_fd_sc_hd__mux2_1 _28747_ (.A0(_01212_),
    .A1(\cpuregs_rs1[1] ),
    .S(instr_timer),
    .X(_01213_));
 sky130_fd_sc_hd__mux2_1 _28748_ (.A0(_01212_),
    .A1(_01213_),
    .S(\cpu_state[2] ),
    .X(_02422_));
 sky130_fd_sc_hd__mux2_1 _28749_ (.A0(_01209_),
    .A1(\cpuregs_rs1[0] ),
    .S(instr_timer),
    .X(_01210_));
 sky130_fd_sc_hd__mux2_1 _28750_ (.A0(_01209_),
    .A1(_01210_),
    .S(\cpu_state[2] ),
    .X(_02411_));
 sky130_fd_sc_hd__mux4_2 _28751_ (.A0(_01202_),
    .A1(_01203_),
    .A2(_01204_),
    .A3(_01205_),
    .S0(net440),
    .S1(net449),
    .X(_01206_));
 sky130_fd_sc_hd__mux4_2 _28752_ (.A0(_01181_),
    .A1(_01182_),
    .A2(_01183_),
    .A3(_01184_),
    .S0(net440),
    .S1(net449),
    .X(_01185_));
 sky130_fd_sc_hd__mux4_2 _28753_ (.A0(_01186_),
    .A1(_01187_),
    .A2(_01188_),
    .A3(_01189_),
    .S0(net443),
    .S1(_00358_),
    .X(_01190_));
 sky130_fd_sc_hd__mux4_2 _28754_ (.A0(_01191_),
    .A1(_01192_),
    .A2(_01193_),
    .A3(_01194_),
    .S0(net443),
    .S1(_00358_),
    .X(_01195_));
 sky130_fd_sc_hd__mux4_1 _28755_ (.A0(_01196_),
    .A1(_01197_),
    .A2(_01198_),
    .A3(_01199_),
    .S0(net443),
    .S1(_00358_),
    .X(_01200_));
 sky130_fd_sc_hd__mux4_1 _28756_ (.A0(_01185_),
    .A1(_01190_),
    .A2(_01195_),
    .A3(_01200_),
    .S0(net452),
    .S1(net454),
    .X(_01201_));
 sky130_fd_sc_hd__mux4_2 _28757_ (.A0(_01175_),
    .A1(_01176_),
    .A2(_01177_),
    .A3(_01178_),
    .S0(net440),
    .S1(net449),
    .X(_01179_));
 sky130_fd_sc_hd__mux4_2 _28758_ (.A0(_01154_),
    .A1(_01155_),
    .A2(_01156_),
    .A3(_01157_),
    .S0(net440),
    .S1(net449),
    .X(_01158_));
 sky130_fd_sc_hd__mux4_2 _28759_ (.A0(_01159_),
    .A1(_01160_),
    .A2(_01161_),
    .A3(_01162_),
    .S0(net443),
    .S1(_00358_),
    .X(_01163_));
 sky130_fd_sc_hd__mux4_2 _28760_ (.A0(_01164_),
    .A1(_01165_),
    .A2(_01166_),
    .A3(_01167_),
    .S0(net443),
    .S1(_00358_),
    .X(_01168_));
 sky130_fd_sc_hd__mux4_1 _28761_ (.A0(_01169_),
    .A1(_01170_),
    .A2(_01171_),
    .A3(_01172_),
    .S0(net443),
    .S1(_00358_),
    .X(_01173_));
 sky130_fd_sc_hd__mux4_1 _28762_ (.A0(_01158_),
    .A1(_01163_),
    .A2(_01168_),
    .A3(_01173_),
    .S0(net452),
    .S1(net454),
    .X(_01174_));
 sky130_fd_sc_hd__mux4_2 _28763_ (.A0(_01148_),
    .A1(_01149_),
    .A2(_01150_),
    .A3(_01151_),
    .S0(net440),
    .S1(net449),
    .X(_01152_));
 sky130_fd_sc_hd__mux4_2 _28764_ (.A0(_01127_),
    .A1(_01128_),
    .A2(_01129_),
    .A3(_01130_),
    .S0(net440),
    .S1(net449),
    .X(_01131_));
 sky130_fd_sc_hd__mux4_2 _28765_ (.A0(_01132_),
    .A1(_01133_),
    .A2(_01134_),
    .A3(_01135_),
    .S0(net443),
    .S1(_00358_),
    .X(_01136_));
 sky130_fd_sc_hd__mux4_2 _28766_ (.A0(_01137_),
    .A1(_01138_),
    .A2(_01139_),
    .A3(_01140_),
    .S0(net443),
    .S1(_00358_),
    .X(_01141_));
 sky130_fd_sc_hd__mux4_1 _28767_ (.A0(_01142_),
    .A1(_01143_),
    .A2(_01144_),
    .A3(_01145_),
    .S0(net443),
    .S1(_00358_),
    .X(_01146_));
 sky130_fd_sc_hd__mux4_1 _28768_ (.A0(_01131_),
    .A1(_01136_),
    .A2(_01141_),
    .A3(_01146_),
    .S0(net452),
    .S1(net454),
    .X(_01147_));
 sky130_fd_sc_hd__mux4_2 _28769_ (.A0(_01121_),
    .A1(_01122_),
    .A2(_01123_),
    .A3(_01124_),
    .S0(net440),
    .S1(net449),
    .X(_01125_));
 sky130_fd_sc_hd__mux4_2 _28770_ (.A0(_01100_),
    .A1(_01101_),
    .A2(_01102_),
    .A3(_01103_),
    .S0(net440),
    .S1(net449),
    .X(_01104_));
 sky130_fd_sc_hd__mux4_2 _28771_ (.A0(_01105_),
    .A1(_01106_),
    .A2(_01107_),
    .A3(_01108_),
    .S0(net443),
    .S1(_00358_),
    .X(_01109_));
 sky130_fd_sc_hd__mux4_2 _28772_ (.A0(_01110_),
    .A1(_01111_),
    .A2(_01112_),
    .A3(_01113_),
    .S0(net443),
    .S1(_00358_),
    .X(_01114_));
 sky130_fd_sc_hd__mux4_1 _28773_ (.A0(_01115_),
    .A1(_01116_),
    .A2(_01117_),
    .A3(_01118_),
    .S0(net443),
    .S1(_00358_),
    .X(_01119_));
 sky130_fd_sc_hd__mux4_1 _28774_ (.A0(_01104_),
    .A1(_01109_),
    .A2(_01114_),
    .A3(_01119_),
    .S0(net452),
    .S1(net454),
    .X(_01120_));
 sky130_fd_sc_hd__mux4_2 _28775_ (.A0(_01094_),
    .A1(_01095_),
    .A2(_01096_),
    .A3(_01097_),
    .S0(net440),
    .S1(net449),
    .X(_01098_));
 sky130_fd_sc_hd__mux4_2 _28776_ (.A0(_01073_),
    .A1(_01074_),
    .A2(_01075_),
    .A3(_01076_),
    .S0(net440),
    .S1(net449),
    .X(_01077_));
 sky130_fd_sc_hd__mux4_2 _28777_ (.A0(_01078_),
    .A1(_01079_),
    .A2(_01080_),
    .A3(_01081_),
    .S0(net441),
    .S1(net449),
    .X(_01082_));
 sky130_fd_sc_hd__mux4_2 _28778_ (.A0(_01083_),
    .A1(_01084_),
    .A2(_01085_),
    .A3(_01086_),
    .S0(net442),
    .S1(net450),
    .X(_01087_));
 sky130_fd_sc_hd__mux4_1 _28779_ (.A0(_01088_),
    .A1(_01089_),
    .A2(_01090_),
    .A3(_01091_),
    .S0(net441),
    .S1(net449),
    .X(_01092_));
 sky130_fd_sc_hd__mux4_2 _28780_ (.A0(_01077_),
    .A1(_01082_),
    .A2(_01087_),
    .A3(_01092_),
    .S0(net452),
    .S1(net454),
    .X(_01093_));
 sky130_fd_sc_hd__mux4_2 _28781_ (.A0(_01067_),
    .A1(_01068_),
    .A2(_01069_),
    .A3(_01070_),
    .S0(net441),
    .S1(net449),
    .X(_01071_));
 sky130_fd_sc_hd__mux4_2 _28782_ (.A0(_01046_),
    .A1(_01047_),
    .A2(_01048_),
    .A3(_01049_),
    .S0(net440),
    .S1(net449),
    .X(_01050_));
 sky130_fd_sc_hd__mux4_2 _28783_ (.A0(_01051_),
    .A1(_01052_),
    .A2(_01053_),
    .A3(_01054_),
    .S0(net441),
    .S1(net449),
    .X(_01055_));
 sky130_fd_sc_hd__mux4_2 _28784_ (.A0(_01056_),
    .A1(_01057_),
    .A2(_01058_),
    .A3(_01059_),
    .S0(net442),
    .S1(net450),
    .X(_01060_));
 sky130_fd_sc_hd__mux4_1 _28785_ (.A0(_01061_),
    .A1(_01062_),
    .A2(_01063_),
    .A3(_01064_),
    .S0(net441),
    .S1(net449),
    .X(_01065_));
 sky130_fd_sc_hd__mux4_1 _28786_ (.A0(_01050_),
    .A1(_01055_),
    .A2(_01060_),
    .A3(_01065_),
    .S0(net452),
    .S1(net454),
    .X(_01066_));
 sky130_fd_sc_hd__mux4_2 _28787_ (.A0(_01040_),
    .A1(_01041_),
    .A2(_01042_),
    .A3(_01043_),
    .S0(net440),
    .S1(net449),
    .X(_01044_));
 sky130_fd_sc_hd__mux4_2 _28788_ (.A0(_01019_),
    .A1(_01020_),
    .A2(_01021_),
    .A3(_01022_),
    .S0(net440),
    .S1(net449),
    .X(_01023_));
 sky130_fd_sc_hd__mux4_2 _28789_ (.A0(_01024_),
    .A1(_01025_),
    .A2(_01026_),
    .A3(_01027_),
    .S0(net441),
    .S1(net449),
    .X(_01028_));
 sky130_fd_sc_hd__mux4_2 _28790_ (.A0(_01029_),
    .A1(_01030_),
    .A2(_01031_),
    .A3(_01032_),
    .S0(net442),
    .S1(net450),
    .X(_01033_));
 sky130_fd_sc_hd__mux4_1 _28791_ (.A0(_01034_),
    .A1(_01035_),
    .A2(_01036_),
    .A3(_01037_),
    .S0(net441),
    .S1(net449),
    .X(_01038_));
 sky130_fd_sc_hd__mux4_2 _28792_ (.A0(_01023_),
    .A1(_01028_),
    .A2(_01033_),
    .A3(_01038_),
    .S0(net452),
    .S1(net454),
    .X(_01039_));
 sky130_fd_sc_hd__mux4_2 _28793_ (.A0(_01013_),
    .A1(_01014_),
    .A2(_01015_),
    .A3(_01016_),
    .S0(net441),
    .S1(net449),
    .X(_01017_));
 sky130_fd_sc_hd__mux4_2 _28794_ (.A0(_00992_),
    .A1(_00993_),
    .A2(_00994_),
    .A3(_00995_),
    .S0(net440),
    .S1(net449),
    .X(_00996_));
 sky130_fd_sc_hd__mux4_2 _28795_ (.A0(_00997_),
    .A1(_00998_),
    .A2(_00999_),
    .A3(_01000_),
    .S0(net441),
    .S1(net449),
    .X(_01001_));
 sky130_fd_sc_hd__mux4_2 _28796_ (.A0(_01002_),
    .A1(_01003_),
    .A2(_01004_),
    .A3(_01005_),
    .S0(net443),
    .S1(_00358_),
    .X(_01006_));
 sky130_fd_sc_hd__mux4_1 _28797_ (.A0(_01007_),
    .A1(_01008_),
    .A2(_01009_),
    .A3(_01010_),
    .S0(net441),
    .S1(net449),
    .X(_01011_));
 sky130_fd_sc_hd__mux4_1 _28798_ (.A0(_00996_),
    .A1(_01001_),
    .A2(_01006_),
    .A3(_01011_),
    .S0(net452),
    .S1(net454),
    .X(_01012_));
 sky130_fd_sc_hd__mux4_1 _28799_ (.A0(_00986_),
    .A1(_00987_),
    .A2(_00988_),
    .A3(_00989_),
    .S0(net442),
    .S1(net450),
    .X(_00990_));
 sky130_fd_sc_hd__mux4_2 _28800_ (.A0(_00965_),
    .A1(_00966_),
    .A2(_00967_),
    .A3(_00968_),
    .S0(net442),
    .S1(net450),
    .X(_00969_));
 sky130_fd_sc_hd__mux4_2 _28801_ (.A0(_00970_),
    .A1(_00971_),
    .A2(_00972_),
    .A3(_00973_),
    .S0(net439),
    .S1(net450),
    .X(_00974_));
 sky130_fd_sc_hd__mux4_2 _28802_ (.A0(_00975_),
    .A1(_00976_),
    .A2(_00977_),
    .A3(_00978_),
    .S0(net439),
    .S1(net450),
    .X(_00979_));
 sky130_fd_sc_hd__mux4_1 _28803_ (.A0(_00980_),
    .A1(_00981_),
    .A2(_00982_),
    .A3(_00983_),
    .S0(net442),
    .S1(net450),
    .X(_00984_));
 sky130_fd_sc_hd__mux4_2 _28804_ (.A0(_00969_),
    .A1(_00974_),
    .A2(_00979_),
    .A3(_00984_),
    .S0(net452),
    .S1(net454),
    .X(_00985_));
 sky130_fd_sc_hd__mux4_1 _28805_ (.A0(_00959_),
    .A1(_00960_),
    .A2(_00961_),
    .A3(_00962_),
    .S0(net442),
    .S1(net450),
    .X(_00963_));
 sky130_fd_sc_hd__mux4_2 _28806_ (.A0(_00938_),
    .A1(_00939_),
    .A2(_00940_),
    .A3(_00941_),
    .S0(net442),
    .S1(net450),
    .X(_00942_));
 sky130_fd_sc_hd__mux4_2 _28807_ (.A0(_00943_),
    .A1(_00944_),
    .A2(_00945_),
    .A3(_00946_),
    .S0(net439),
    .S1(net450),
    .X(_00947_));
 sky130_fd_sc_hd__mux4_2 _28808_ (.A0(_00948_),
    .A1(_00949_),
    .A2(_00950_),
    .A3(_00951_),
    .S0(net439),
    .S1(net450),
    .X(_00952_));
 sky130_fd_sc_hd__mux4_1 _28809_ (.A0(_00953_),
    .A1(_00954_),
    .A2(_00955_),
    .A3(_00956_),
    .S0(net442),
    .S1(net450),
    .X(_00957_));
 sky130_fd_sc_hd__mux4_2 _28810_ (.A0(_00942_),
    .A1(_00947_),
    .A2(_00952_),
    .A3(_00957_),
    .S0(net452),
    .S1(net454),
    .X(_00958_));
 sky130_fd_sc_hd__mux4_1 _28811_ (.A0(_00932_),
    .A1(_00933_),
    .A2(_00934_),
    .A3(_00935_),
    .S0(net442),
    .S1(net450),
    .X(_00936_));
 sky130_fd_sc_hd__mux4_2 _28812_ (.A0(_00911_),
    .A1(_00912_),
    .A2(_00913_),
    .A3(_00914_),
    .S0(net442),
    .S1(net450),
    .X(_00915_));
 sky130_fd_sc_hd__mux4_2 _28813_ (.A0(_00916_),
    .A1(_00917_),
    .A2(_00918_),
    .A3(_00919_),
    .S0(net439),
    .S1(net450),
    .X(_00920_));
 sky130_fd_sc_hd__mux4_2 _28814_ (.A0(_00921_),
    .A1(_00922_),
    .A2(_00923_),
    .A3(_00924_),
    .S0(net439),
    .S1(net448),
    .X(_00925_));
 sky130_fd_sc_hd__mux4_2 _28815_ (.A0(_00926_),
    .A1(_00927_),
    .A2(_00928_),
    .A3(_00929_),
    .S0(net442),
    .S1(net450),
    .X(_00930_));
 sky130_fd_sc_hd__mux4_2 _28816_ (.A0(_00915_),
    .A1(_00920_),
    .A2(_00925_),
    .A3(_00930_),
    .S0(net452),
    .S1(net454),
    .X(_00931_));
 sky130_fd_sc_hd__mux4_1 _28817_ (.A0(_00905_),
    .A1(_00906_),
    .A2(_00907_),
    .A3(_00908_),
    .S0(net442),
    .S1(net450),
    .X(_00909_));
 sky130_fd_sc_hd__mux4_2 _28818_ (.A0(_00884_),
    .A1(_00885_),
    .A2(_00886_),
    .A3(_00887_),
    .S0(net442),
    .S1(net450),
    .X(_00888_));
 sky130_fd_sc_hd__mux4_2 _28819_ (.A0(_00889_),
    .A1(_00890_),
    .A2(_00891_),
    .A3(_00892_),
    .S0(net439),
    .S1(net450),
    .X(_00893_));
 sky130_fd_sc_hd__mux4_2 _28820_ (.A0(_00894_),
    .A1(_00895_),
    .A2(_00896_),
    .A3(_00897_),
    .S0(net439),
    .S1(net448),
    .X(_00898_));
 sky130_fd_sc_hd__mux4_2 _28821_ (.A0(_00899_),
    .A1(_00900_),
    .A2(_00901_),
    .A3(_00902_),
    .S0(net442),
    .S1(net450),
    .X(_00903_));
 sky130_fd_sc_hd__mux4_2 _28822_ (.A0(_00888_),
    .A1(_00893_),
    .A2(_00898_),
    .A3(_00903_),
    .S0(net452),
    .S1(net454),
    .X(_00904_));
 sky130_fd_sc_hd__mux4_1 _28823_ (.A0(_00878_),
    .A1(_00879_),
    .A2(_00880_),
    .A3(_00881_),
    .S0(net439),
    .S1(net448),
    .X(_00882_));
 sky130_fd_sc_hd__mux4_2 _28824_ (.A0(_00857_),
    .A1(_00858_),
    .A2(_00859_),
    .A3(_00860_),
    .S0(net438),
    .S1(net448),
    .X(_00861_));
 sky130_fd_sc_hd__mux4_1 _28825_ (.A0(_00862_),
    .A1(_00863_),
    .A2(_00864_),
    .A3(_00865_),
    .S0(net438),
    .S1(net448),
    .X(_00866_));
 sky130_fd_sc_hd__mux4_2 _28826_ (.A0(_00867_),
    .A1(_00868_),
    .A2(_00869_),
    .A3(_00870_),
    .S0(net437),
    .S1(net447),
    .X(_00871_));
 sky130_fd_sc_hd__mux4_1 _28827_ (.A0(_00872_),
    .A1(_00873_),
    .A2(_00874_),
    .A3(_00875_),
    .S0(net438),
    .S1(net448),
    .X(_00876_));
 sky130_fd_sc_hd__mux4_2 _28828_ (.A0(_00861_),
    .A1(_00866_),
    .A2(_00871_),
    .A3(_00876_),
    .S0(_00360_),
    .S1(net453),
    .X(_00877_));
 sky130_fd_sc_hd__mux4_1 _28829_ (.A0(_00851_),
    .A1(_00852_),
    .A2(_00853_),
    .A3(_00854_),
    .S0(net438),
    .S1(net448),
    .X(_00855_));
 sky130_fd_sc_hd__mux4_2 _28830_ (.A0(_00830_),
    .A1(_00831_),
    .A2(_00832_),
    .A3(_00833_),
    .S0(net438),
    .S1(net448),
    .X(_00834_));
 sky130_fd_sc_hd__mux4_2 _28831_ (.A0(_00835_),
    .A1(_00836_),
    .A2(_00837_),
    .A3(_00838_),
    .S0(net438),
    .S1(net448),
    .X(_00839_));
 sky130_fd_sc_hd__mux4_2 _28832_ (.A0(_00840_),
    .A1(_00841_),
    .A2(_00842_),
    .A3(_00843_),
    .S0(net438),
    .S1(net448),
    .X(_00844_));
 sky130_fd_sc_hd__mux4_1 _28833_ (.A0(_00845_),
    .A1(_00846_),
    .A2(_00847_),
    .A3(_00848_),
    .S0(net438),
    .S1(net448),
    .X(_00849_));
 sky130_fd_sc_hd__mux4_2 _28834_ (.A0(_00834_),
    .A1(_00839_),
    .A2(_00844_),
    .A3(_00849_),
    .S0(_00360_),
    .S1(net453),
    .X(_00850_));
 sky130_fd_sc_hd__mux4_1 _28835_ (.A0(_00824_),
    .A1(_00825_),
    .A2(_00826_),
    .A3(_00827_),
    .S0(net439),
    .S1(net448),
    .X(_00828_));
 sky130_fd_sc_hd__mux4_2 _28836_ (.A0(_00803_),
    .A1(_00804_),
    .A2(_00805_),
    .A3(_00806_),
    .S0(net438),
    .S1(net448),
    .X(_00807_));
 sky130_fd_sc_hd__mux4_1 _28837_ (.A0(_00808_),
    .A1(_00809_),
    .A2(_00810_),
    .A3(_00811_),
    .S0(net438),
    .S1(net448),
    .X(_00812_));
 sky130_fd_sc_hd__mux4_2 _28838_ (.A0(_00813_),
    .A1(_00814_),
    .A2(_00815_),
    .A3(_00816_),
    .S0(net437),
    .S1(net447),
    .X(_00817_));
 sky130_fd_sc_hd__mux4_1 _28839_ (.A0(_00818_),
    .A1(_00819_),
    .A2(_00820_),
    .A3(_00821_),
    .S0(net438),
    .S1(net448),
    .X(_00822_));
 sky130_fd_sc_hd__mux4_2 _28840_ (.A0(_00807_),
    .A1(_00812_),
    .A2(_00817_),
    .A3(_00822_),
    .S0(_00360_),
    .S1(net453),
    .X(_00823_));
 sky130_fd_sc_hd__mux4_1 _28841_ (.A0(_00797_),
    .A1(_00798_),
    .A2(_00799_),
    .A3(_00800_),
    .S0(net439),
    .S1(net448),
    .X(_00801_));
 sky130_fd_sc_hd__mux4_1 _28842_ (.A0(_00776_),
    .A1(_00777_),
    .A2(_00778_),
    .A3(_00779_),
    .S0(net438),
    .S1(net448),
    .X(_00780_));
 sky130_fd_sc_hd__mux4_2 _28843_ (.A0(_00781_),
    .A1(_00782_),
    .A2(_00783_),
    .A3(_00784_),
    .S0(net438),
    .S1(net448),
    .X(_00785_));
 sky130_fd_sc_hd__mux4_2 _28844_ (.A0(_00786_),
    .A1(_00787_),
    .A2(_00788_),
    .A3(_00789_),
    .S0(net438),
    .S1(net448),
    .X(_00790_));
 sky130_fd_sc_hd__mux4_1 _28845_ (.A0(_00791_),
    .A1(_00792_),
    .A2(_00793_),
    .A3(_00794_),
    .S0(net438),
    .S1(net448),
    .X(_00795_));
 sky130_fd_sc_hd__mux4_2 _28846_ (.A0(_00780_),
    .A1(_00785_),
    .A2(_00790_),
    .A3(_00795_),
    .S0(_00360_),
    .S1(net453),
    .X(_00796_));
 sky130_fd_sc_hd__mux4_1 _28847_ (.A0(_00770_),
    .A1(_00771_),
    .A2(_00772_),
    .A3(_00773_),
    .S0(net435),
    .S1(net444),
    .X(_00774_));
 sky130_fd_sc_hd__mux4_2 _28848_ (.A0(_00749_),
    .A1(_00750_),
    .A2(_00751_),
    .A3(_00752_),
    .S0(net432),
    .S1(net444),
    .X(_00753_));
 sky130_fd_sc_hd__mux4_2 _28849_ (.A0(_00754_),
    .A1(_00755_),
    .A2(_00756_),
    .A3(_00757_),
    .S0(net436),
    .S1(net445),
    .X(_00758_));
 sky130_fd_sc_hd__mux4_2 _28850_ (.A0(_00759_),
    .A1(_00760_),
    .A2(_00761_),
    .A3(_00762_),
    .S0(net434),
    .S1(net445),
    .X(_00763_));
 sky130_fd_sc_hd__mux4_1 _28851_ (.A0(_00764_),
    .A1(_00765_),
    .A2(_00766_),
    .A3(_00767_),
    .S0(net435),
    .S1(net444),
    .X(_00768_));
 sky130_fd_sc_hd__mux4_2 _28852_ (.A0(_00753_),
    .A1(_00758_),
    .A2(_00763_),
    .A3(_00768_),
    .S0(net451),
    .S1(net453),
    .X(_00769_));
 sky130_fd_sc_hd__mux4_1 _28853_ (.A0(_00743_),
    .A1(_00744_),
    .A2(_00745_),
    .A3(_00746_),
    .S0(net435),
    .S1(net444),
    .X(_00747_));
 sky130_fd_sc_hd__mux4_2 _28854_ (.A0(_00722_),
    .A1(_00723_),
    .A2(_00724_),
    .A3(_00725_),
    .S0(net432),
    .S1(net444),
    .X(_00726_));
 sky130_fd_sc_hd__mux4_2 _28855_ (.A0(_00727_),
    .A1(_00728_),
    .A2(_00729_),
    .A3(_00730_),
    .S0(net436),
    .S1(net445),
    .X(_00731_));
 sky130_fd_sc_hd__mux4_2 _28856_ (.A0(_00732_),
    .A1(_00733_),
    .A2(_00734_),
    .A3(_00735_),
    .S0(net434),
    .S1(net445),
    .X(_00736_));
 sky130_fd_sc_hd__mux4_1 _28857_ (.A0(_00737_),
    .A1(_00738_),
    .A2(_00739_),
    .A3(_00740_),
    .S0(net435),
    .S1(net444),
    .X(_00741_));
 sky130_fd_sc_hd__mux4_2 _28858_ (.A0(_00726_),
    .A1(_00731_),
    .A2(_00736_),
    .A3(_00741_),
    .S0(net451),
    .S1(net453),
    .X(_00742_));
 sky130_fd_sc_hd__mux4_1 _28859_ (.A0(_00716_),
    .A1(_00717_),
    .A2(_00718_),
    .A3(_00719_),
    .S0(net432),
    .S1(net444),
    .X(_00720_));
 sky130_fd_sc_hd__mux4_2 _28860_ (.A0(_00695_),
    .A1(_00696_),
    .A2(_00697_),
    .A3(_00698_),
    .S0(net432),
    .S1(net444),
    .X(_00699_));
 sky130_fd_sc_hd__mux4_2 _28861_ (.A0(_00700_),
    .A1(_00701_),
    .A2(_00702_),
    .A3(_00703_),
    .S0(net436),
    .S1(net445),
    .X(_00704_));
 sky130_fd_sc_hd__mux4_2 _28862_ (.A0(_00705_),
    .A1(_00706_),
    .A2(_00707_),
    .A3(_00708_),
    .S0(net434),
    .S1(net445),
    .X(_00709_));
 sky130_fd_sc_hd__mux4_1 _28863_ (.A0(_00710_),
    .A1(_00711_),
    .A2(_00712_),
    .A3(_00713_),
    .S0(net436),
    .S1(net445),
    .X(_00714_));
 sky130_fd_sc_hd__mux4_2 _28864_ (.A0(_00699_),
    .A1(_00704_),
    .A2(_00709_),
    .A3(_00714_),
    .S0(net451),
    .S1(net453),
    .X(_00715_));
 sky130_fd_sc_hd__mux4_1 _28865_ (.A0(_00689_),
    .A1(_00690_),
    .A2(_00691_),
    .A3(_00692_),
    .S0(net435),
    .S1(net444),
    .X(_00693_));
 sky130_fd_sc_hd__mux4_2 _28866_ (.A0(_00668_),
    .A1(_00669_),
    .A2(_00670_),
    .A3(_00671_),
    .S0(net432),
    .S1(net444),
    .X(_00672_));
 sky130_fd_sc_hd__mux4_2 _28867_ (.A0(_00673_),
    .A1(_00674_),
    .A2(_00675_),
    .A3(_00676_),
    .S0(net436),
    .S1(net445),
    .X(_00677_));
 sky130_fd_sc_hd__mux4_2 _28868_ (.A0(_00678_),
    .A1(_00679_),
    .A2(_00680_),
    .A3(_00681_),
    .S0(net434),
    .S1(net445),
    .X(_00682_));
 sky130_fd_sc_hd__mux4_1 _28869_ (.A0(_00683_),
    .A1(_00684_),
    .A2(_00685_),
    .A3(_00686_),
    .S0(net432),
    .S1(net444),
    .X(_00687_));
 sky130_fd_sc_hd__mux4_2 _28870_ (.A0(_00672_),
    .A1(_00677_),
    .A2(_00682_),
    .A3(_00687_),
    .S0(net451),
    .S1(net453),
    .X(_00688_));
 sky130_fd_sc_hd__mux4_2 _28871_ (.A0(_00662_),
    .A1(_00663_),
    .A2(_00664_),
    .A3(_00665_),
    .S0(net432),
    .S1(net444),
    .X(_00666_));
 sky130_fd_sc_hd__mux4_2 _28872_ (.A0(_00641_),
    .A1(_00642_),
    .A2(_00643_),
    .A3(_00644_),
    .S0(net432),
    .S1(net444),
    .X(_00645_));
 sky130_fd_sc_hd__mux4_1 _28873_ (.A0(_00646_),
    .A1(_00647_),
    .A2(_00648_),
    .A3(_00649_),
    .S0(net434),
    .S1(net445),
    .X(_00650_));
 sky130_fd_sc_hd__mux4_2 _28874_ (.A0(_00651_),
    .A1(_00652_),
    .A2(_00653_),
    .A3(_00654_),
    .S0(net434),
    .S1(net445),
    .X(_00655_));
 sky130_fd_sc_hd__mux4_1 _28875_ (.A0(_00656_),
    .A1(_00657_),
    .A2(_00658_),
    .A3(_00659_),
    .S0(net434),
    .S1(net445),
    .X(_00660_));
 sky130_fd_sc_hd__mux4_2 _28876_ (.A0(_00645_),
    .A1(_00650_),
    .A2(_00655_),
    .A3(_00660_),
    .S0(net451),
    .S1(net453),
    .X(_00661_));
 sky130_fd_sc_hd__mux4_2 _28877_ (.A0(_00635_),
    .A1(_00636_),
    .A2(_00637_),
    .A3(_00638_),
    .S0(net432),
    .S1(net444),
    .X(_00639_));
 sky130_fd_sc_hd__mux4_2 _28878_ (.A0(_00614_),
    .A1(_00615_),
    .A2(_00616_),
    .A3(_00617_),
    .S0(net432),
    .S1(net444),
    .X(_00618_));
 sky130_fd_sc_hd__mux4_2 _28879_ (.A0(_00619_),
    .A1(_00620_),
    .A2(_00621_),
    .A3(_00622_),
    .S0(net434),
    .S1(net445),
    .X(_00623_));
 sky130_fd_sc_hd__mux4_2 _28880_ (.A0(_00624_),
    .A1(_00625_),
    .A2(_00626_),
    .A3(_00627_),
    .S0(net434),
    .S1(net445),
    .X(_00628_));
 sky130_fd_sc_hd__mux4_1 _28881_ (.A0(_00629_),
    .A1(_00630_),
    .A2(_00631_),
    .A3(_00632_),
    .S0(net432),
    .S1(net444),
    .X(_00633_));
 sky130_fd_sc_hd__mux4_2 _28882_ (.A0(_00618_),
    .A1(_00623_),
    .A2(_00628_),
    .A3(_00633_),
    .S0(net451),
    .S1(net453),
    .X(_00634_));
 sky130_fd_sc_hd__mux4_1 _28883_ (.A0(_00608_),
    .A1(_00609_),
    .A2(_00610_),
    .A3(_00611_),
    .S0(net432),
    .S1(net444),
    .X(_00612_));
 sky130_fd_sc_hd__mux4_1 _28884_ (.A0(_00587_),
    .A1(_00588_),
    .A2(_00589_),
    .A3(_00590_),
    .S0(net432),
    .S1(net444),
    .X(_00591_));
 sky130_fd_sc_hd__mux4_2 _28885_ (.A0(_00592_),
    .A1(_00593_),
    .A2(_00594_),
    .A3(_00595_),
    .S0(net434),
    .S1(net445),
    .X(_00596_));
 sky130_fd_sc_hd__mux4_2 _28886_ (.A0(_00597_),
    .A1(_00598_),
    .A2(_00599_),
    .A3(_00600_),
    .S0(net434),
    .S1(net445),
    .X(_00601_));
 sky130_fd_sc_hd__mux4_1 _28887_ (.A0(_00602_),
    .A1(_00603_),
    .A2(_00604_),
    .A3(_00605_),
    .S0(net432),
    .S1(net444),
    .X(_00606_));
 sky130_fd_sc_hd__mux4_2 _28888_ (.A0(_00591_),
    .A1(_00596_),
    .A2(_00601_),
    .A3(_00606_),
    .S0(net451),
    .S1(net453),
    .X(_00607_));
 sky130_fd_sc_hd__mux4_2 _28889_ (.A0(_00581_),
    .A1(_00582_),
    .A2(_00583_),
    .A3(_00584_),
    .S0(net432),
    .S1(net444),
    .X(_00585_));
 sky130_fd_sc_hd__mux4_2 _28890_ (.A0(_00560_),
    .A1(_00561_),
    .A2(_00562_),
    .A3(_00563_),
    .S0(net432),
    .S1(net444),
    .X(_00564_));
 sky130_fd_sc_hd__mux4_2 _28891_ (.A0(_00565_),
    .A1(_00566_),
    .A2(_00567_),
    .A3(_00568_),
    .S0(net434),
    .S1(net445),
    .X(_00569_));
 sky130_fd_sc_hd__mux4_2 _28892_ (.A0(_00570_),
    .A1(_00571_),
    .A2(_00572_),
    .A3(_00573_),
    .S0(net434),
    .S1(net445),
    .X(_00574_));
 sky130_fd_sc_hd__mux4_1 _28893_ (.A0(_00575_),
    .A1(_00576_),
    .A2(_00577_),
    .A3(_00578_),
    .S0(net434),
    .S1(net445),
    .X(_00579_));
 sky130_fd_sc_hd__mux4_2 _28894_ (.A0(_00564_),
    .A1(_00569_),
    .A2(_00574_),
    .A3(_00579_),
    .S0(net451),
    .S1(net453),
    .X(_00580_));
 sky130_fd_sc_hd__mux4_1 _28895_ (.A0(_00554_),
    .A1(_00555_),
    .A2(_00556_),
    .A3(_00557_),
    .S0(net433),
    .S1(net446),
    .X(_00558_));
 sky130_fd_sc_hd__mux4_2 _28896_ (.A0(_00533_),
    .A1(_00534_),
    .A2(_00535_),
    .A3(_00536_),
    .S0(net433),
    .S1(net446),
    .X(_00537_));
 sky130_fd_sc_hd__mux4_2 _28897_ (.A0(_00538_),
    .A1(_00539_),
    .A2(_00540_),
    .A3(_00541_),
    .S0(net435),
    .S1(net446),
    .X(_00542_));
 sky130_fd_sc_hd__mux4_2 _28898_ (.A0(_00543_),
    .A1(_00544_),
    .A2(_00545_),
    .A3(_00546_),
    .S0(net436),
    .S1(net447),
    .X(_00547_));
 sky130_fd_sc_hd__mux4_1 _28899_ (.A0(_00548_),
    .A1(_00549_),
    .A2(_00550_),
    .A3(_00551_),
    .S0(net435),
    .S1(net444),
    .X(_00552_));
 sky130_fd_sc_hd__mux4_2 _28900_ (.A0(_00537_),
    .A1(_00542_),
    .A2(_00547_),
    .A3(_00552_),
    .S0(net451),
    .S1(net453),
    .X(_00553_));
 sky130_fd_sc_hd__mux4_1 _28901_ (.A0(_00527_),
    .A1(_00528_),
    .A2(_00529_),
    .A3(_00530_),
    .S0(net433),
    .S1(net446),
    .X(_00531_));
 sky130_fd_sc_hd__mux4_2 _28902_ (.A0(_00506_),
    .A1(_00507_),
    .A2(_00508_),
    .A3(_00509_),
    .S0(net433),
    .S1(net446),
    .X(_00510_));
 sky130_fd_sc_hd__mux4_2 _28903_ (.A0(_00511_),
    .A1(_00512_),
    .A2(_00513_),
    .A3(_00514_),
    .S0(net436),
    .S1(net446),
    .X(_00515_));
 sky130_fd_sc_hd__mux4_2 _28904_ (.A0(_00516_),
    .A1(_00517_),
    .A2(_00518_),
    .A3(_00519_),
    .S0(net436),
    .S1(net446),
    .X(_00520_));
 sky130_fd_sc_hd__mux4_1 _28905_ (.A0(_00521_),
    .A1(_00522_),
    .A2(_00523_),
    .A3(_00524_),
    .S0(net435),
    .S1(net446),
    .X(_00525_));
 sky130_fd_sc_hd__mux4_2 _28906_ (.A0(_00510_),
    .A1(_00515_),
    .A2(_00520_),
    .A3(_00525_),
    .S0(net451),
    .S1(net453),
    .X(_00526_));
 sky130_fd_sc_hd__mux4_1 _28907_ (.A0(_00500_),
    .A1(_00501_),
    .A2(_00502_),
    .A3(_00503_),
    .S0(net433),
    .S1(net446),
    .X(_00504_));
 sky130_fd_sc_hd__mux4_2 _28908_ (.A0(_00479_),
    .A1(_00480_),
    .A2(_00481_),
    .A3(_00482_),
    .S0(net433),
    .S1(net446),
    .X(_00483_));
 sky130_fd_sc_hd__mux4_2 _28909_ (.A0(_00484_),
    .A1(_00485_),
    .A2(_00486_),
    .A3(_00487_),
    .S0(net435),
    .S1(net446),
    .X(_00488_));
 sky130_fd_sc_hd__mux4_2 _28910_ (.A0(_00489_),
    .A1(_00490_),
    .A2(_00491_),
    .A3(_00492_),
    .S0(net436),
    .S1(net447),
    .X(_00493_));
 sky130_fd_sc_hd__mux4_1 _28911_ (.A0(_00494_),
    .A1(_00495_),
    .A2(_00496_),
    .A3(_00497_),
    .S0(net433),
    .S1(net446),
    .X(_00498_));
 sky130_fd_sc_hd__mux4_2 _28912_ (.A0(_00483_),
    .A1(_00488_),
    .A2(_00493_),
    .A3(_00498_),
    .S0(net451),
    .S1(net453),
    .X(_00499_));
 sky130_fd_sc_hd__mux4_1 _28913_ (.A0(_00473_),
    .A1(_00474_),
    .A2(_00475_),
    .A3(_00476_),
    .S0(net433),
    .S1(net446),
    .X(_00477_));
 sky130_fd_sc_hd__mux4_2 _28914_ (.A0(_00452_),
    .A1(_00453_),
    .A2(_00454_),
    .A3(_00455_),
    .S0(net433),
    .S1(net446),
    .X(_00456_));
 sky130_fd_sc_hd__mux4_2 _28915_ (.A0(_00457_),
    .A1(_00458_),
    .A2(_00459_),
    .A3(_00460_),
    .S0(net435),
    .S1(net446),
    .X(_00461_));
 sky130_fd_sc_hd__mux4_2 _28916_ (.A0(_00462_),
    .A1(_00463_),
    .A2(_00464_),
    .A3(_00465_),
    .S0(net436),
    .S1(net447),
    .X(_00466_));
 sky130_fd_sc_hd__mux4_1 _28917_ (.A0(_00467_),
    .A1(_00468_),
    .A2(_00469_),
    .A3(_00470_),
    .S0(net435),
    .S1(net446),
    .X(_00471_));
 sky130_fd_sc_hd__mux4_2 _28918_ (.A0(_00456_),
    .A1(_00461_),
    .A2(_00466_),
    .A3(_00471_),
    .S0(net451),
    .S1(net453),
    .X(_00472_));
 sky130_fd_sc_hd__mux4_1 _28919_ (.A0(_00446_),
    .A1(_00447_),
    .A2(_00448_),
    .A3(_00449_),
    .S0(net433),
    .S1(net446),
    .X(_00450_));
 sky130_fd_sc_hd__mux4_2 _28920_ (.A0(_00425_),
    .A1(_00426_),
    .A2(_00427_),
    .A3(_00428_),
    .S0(net437),
    .S1(net447),
    .X(_00429_));
 sky130_fd_sc_hd__mux4_2 _28921_ (.A0(_00430_),
    .A1(_00431_),
    .A2(_00432_),
    .A3(_00433_),
    .S0(net437),
    .S1(net447),
    .X(_00434_));
 sky130_fd_sc_hd__mux4_2 _28922_ (.A0(_00435_),
    .A1(_00436_),
    .A2(_00437_),
    .A3(_00438_),
    .S0(net436),
    .S1(net447),
    .X(_00439_));
 sky130_fd_sc_hd__mux4_1 _28923_ (.A0(_00440_),
    .A1(_00441_),
    .A2(_00442_),
    .A3(_00443_),
    .S0(net437),
    .S1(net447),
    .X(_00444_));
 sky130_fd_sc_hd__mux4_2 _28924_ (.A0(_00429_),
    .A1(_00434_),
    .A2(_00439_),
    .A3(_00444_),
    .S0(net451),
    .S1(net453),
    .X(_00445_));
 sky130_fd_sc_hd__mux4_1 _28925_ (.A0(_00419_),
    .A1(_00420_),
    .A2(_00421_),
    .A3(_00422_),
    .S0(net433),
    .S1(net446),
    .X(_00423_));
 sky130_fd_sc_hd__mux4_2 _28926_ (.A0(_00398_),
    .A1(_00399_),
    .A2(_00400_),
    .A3(_00401_),
    .S0(net437),
    .S1(net447),
    .X(_00402_));
 sky130_fd_sc_hd__mux4_2 _28927_ (.A0(_00403_),
    .A1(_00404_),
    .A2(_00405_),
    .A3(_00406_),
    .S0(net437),
    .S1(net447),
    .X(_00407_));
 sky130_fd_sc_hd__mux4_2 _28928_ (.A0(_00408_),
    .A1(_00409_),
    .A2(_00410_),
    .A3(_00411_),
    .S0(net436),
    .S1(net447),
    .X(_00412_));
 sky130_fd_sc_hd__mux4_1 _28929_ (.A0(_00413_),
    .A1(_00414_),
    .A2(_00415_),
    .A3(_00416_),
    .S0(net437),
    .S1(net447),
    .X(_00417_));
 sky130_fd_sc_hd__mux4_2 _28930_ (.A0(_00402_),
    .A1(_00407_),
    .A2(_00412_),
    .A3(_00417_),
    .S0(_00360_),
    .S1(net453),
    .X(_00418_));
 sky130_fd_sc_hd__mux4_1 _28931_ (.A0(_00392_),
    .A1(_00393_),
    .A2(_00394_),
    .A3(_00395_),
    .S0(net433),
    .S1(net446),
    .X(_00396_));
 sky130_fd_sc_hd__mux4_2 _28932_ (.A0(_00371_),
    .A1(_00372_),
    .A2(_00373_),
    .A3(_00374_),
    .S0(net437),
    .S1(net447),
    .X(_00375_));
 sky130_fd_sc_hd__mux4_2 _28933_ (.A0(_00376_),
    .A1(_00377_),
    .A2(_00378_),
    .A3(_00379_),
    .S0(net437),
    .S1(net447),
    .X(_00380_));
 sky130_fd_sc_hd__mux4_2 _28934_ (.A0(_00381_),
    .A1(_00382_),
    .A2(_00383_),
    .A3(_00384_),
    .S0(net436),
    .S1(net447),
    .X(_00385_));
 sky130_fd_sc_hd__mux4_1 _28935_ (.A0(_00386_),
    .A1(_00387_),
    .A2(_00388_),
    .A3(_00389_),
    .S0(net437),
    .S1(net447),
    .X(_00390_));
 sky130_fd_sc_hd__mux4_2 _28936_ (.A0(_00375_),
    .A1(_00380_),
    .A2(_00385_),
    .A3(_00390_),
    .S0(net451),
    .S1(net453),
    .X(_00391_));
 sky130_fd_sc_hd__mux4_1 _28937_ (.A0(\cpuregs[16][0] ),
    .A1(\cpuregs[17][0] ),
    .A2(\cpuregs[18][0] ),
    .A3(\cpuregs[19][0] ),
    .S0(net433),
    .S1(net446),
    .X(_00369_));
 sky130_fd_sc_hd__mux4_2 _28938_ (.A0(\cpuregs[0][0] ),
    .A1(\cpuregs[1][0] ),
    .A2(\cpuregs[2][0] ),
    .A3(\cpuregs[3][0] ),
    .S0(net437),
    .S1(net447),
    .X(_00359_));
 sky130_fd_sc_hd__mux4_2 _28939_ (.A0(\cpuregs[4][0] ),
    .A1(\cpuregs[5][0] ),
    .A2(\cpuregs[6][0] ),
    .A3(\cpuregs[7][0] ),
    .S0(net437),
    .S1(net447),
    .X(_00361_));
 sky130_fd_sc_hd__mux4_2 _28940_ (.A0(\cpuregs[8][0] ),
    .A1(\cpuregs[9][0] ),
    .A2(\cpuregs[10][0] ),
    .A3(\cpuregs[11][0] ),
    .S0(net437),
    .S1(net447),
    .X(_00363_));
 sky130_fd_sc_hd__mux4_1 _28941_ (.A0(\cpuregs[12][0] ),
    .A1(\cpuregs[13][0] ),
    .A2(\cpuregs[14][0] ),
    .A3(\cpuregs[15][0] ),
    .S0(net437),
    .S1(net447),
    .X(_00364_));
 sky130_fd_sc_hd__mux4_2 _28942_ (.A0(_00359_),
    .A1(_00361_),
    .A2(_00363_),
    .A3(_00364_),
    .S0(_00360_),
    .S1(net453),
    .X(_00365_));
 sky130_fd_sc_hd__mux4_1 _28943_ (.A0(_02581_),
    .A1(_01681_),
    .A2(_01679_),
    .A3(_02581_),
    .S0(net412),
    .S1(net431),
    .X(_01682_));
 sky130_fd_sc_hd__mux4_1 _28944_ (.A0(_02580_),
    .A1(_01677_),
    .A2(_01675_),
    .A3(_02580_),
    .S0(net412),
    .S1(net431),
    .X(_01678_));
 sky130_fd_sc_hd__mux4_1 _28945_ (.A0(_02579_),
    .A1(_01673_),
    .A2(_01671_),
    .A3(_02579_),
    .S0(net412),
    .S1(net431),
    .X(_01674_));
 sky130_fd_sc_hd__mux4_1 _28946_ (.A0(_02578_),
    .A1(_01669_),
    .A2(_01667_),
    .A3(_02578_),
    .S0(net412),
    .S1(net431),
    .X(_01670_));
 sky130_fd_sc_hd__mux4_1 _28947_ (.A0(_02577_),
    .A1(_01665_),
    .A2(_01663_),
    .A3(_02577_),
    .S0(net412),
    .S1(net431),
    .X(_01666_));
 sky130_fd_sc_hd__mux4_1 _28948_ (.A0(_02576_),
    .A1(_01661_),
    .A2(_01659_),
    .A3(_02576_),
    .S0(net412),
    .S1(net431),
    .X(_01662_));
 sky130_fd_sc_hd__mux4_1 _28949_ (.A0(_02575_),
    .A1(_01657_),
    .A2(_01655_),
    .A3(_02575_),
    .S0(net412),
    .S1(net431),
    .X(_01658_));
 sky130_fd_sc_hd__mux4_1 _28950_ (.A0(_02574_),
    .A1(_01653_),
    .A2(_01651_),
    .A3(_02574_),
    .S0(net412),
    .S1(net431),
    .X(_01654_));
 sky130_fd_sc_hd__mux4_1 _28951_ (.A0(_02573_),
    .A1(_01649_),
    .A2(_01647_),
    .A3(_02573_),
    .S0(net412),
    .S1(net431),
    .X(_01650_));
 sky130_fd_sc_hd__mux4_1 _28952_ (.A0(_02572_),
    .A1(_01645_),
    .A2(_01643_),
    .A3(_02572_),
    .S0(net412),
    .S1(net431),
    .X(_01646_));
 sky130_fd_sc_hd__mux4_1 _28953_ (.A0(_02570_),
    .A1(_01641_),
    .A2(_01639_),
    .A3(_02570_),
    .S0(net412),
    .S1(net431),
    .X(_01642_));
 sky130_fd_sc_hd__mux4_1 _28954_ (.A0(_02569_),
    .A1(_01637_),
    .A2(_01635_),
    .A3(_02569_),
    .S0(net412),
    .S1(net431),
    .X(_01638_));
 sky130_fd_sc_hd__mux4_1 _28955_ (.A0(_02568_),
    .A1(_01633_),
    .A2(_01631_),
    .A3(_02568_),
    .S0(net412),
    .S1(net431),
    .X(_01634_));
 sky130_fd_sc_hd__mux4_1 _28956_ (.A0(_02567_),
    .A1(_01629_),
    .A2(_01627_),
    .A3(_02567_),
    .S0(net412),
    .S1(net431),
    .X(_01630_));
 sky130_fd_sc_hd__mux4_1 _28957_ (.A0(_02566_),
    .A1(_01625_),
    .A2(_01623_),
    .A3(_02566_),
    .S0(net412),
    .S1(net431),
    .X(_01626_));
 sky130_fd_sc_hd__mux4_1 _28958_ (.A0(_02565_),
    .A1(_01621_),
    .A2(_01619_),
    .A3(_02565_),
    .S0(net412),
    .S1(net431),
    .X(_01622_));
 sky130_fd_sc_hd__mux4_1 _28959_ (.A0(_02564_),
    .A1(_01617_),
    .A2(_01615_),
    .A3(_02564_),
    .S0(net412),
    .S1(net431),
    .X(_01618_));
 sky130_fd_sc_hd__mux4_1 _28960_ (.A0(_02563_),
    .A1(_01613_),
    .A2(_01611_),
    .A3(_02563_),
    .S0(net412),
    .S1(net431),
    .X(_01614_));
 sky130_fd_sc_hd__mux4_1 _28961_ (.A0(_02562_),
    .A1(_01609_),
    .A2(_01607_),
    .A3(_02562_),
    .S0(net412),
    .S1(net431),
    .X(_01610_));
 sky130_fd_sc_hd__mux4_1 _28962_ (.A0(_02561_),
    .A1(_01605_),
    .A2(_01603_),
    .A3(_02561_),
    .S0(net412),
    .S1(net431),
    .X(_01606_));
 sky130_fd_sc_hd__mux4_1 _28963_ (.A0(_02589_),
    .A1(_01601_),
    .A2(_01599_),
    .A3(_02589_),
    .S0(_14285_),
    .S1(net431),
    .X(_01602_));
 sky130_fd_sc_hd__mux4_1 _28964_ (.A0(_02588_),
    .A1(_01597_),
    .A2(_01595_),
    .A3(_02588_),
    .S0(_14285_),
    .S1(net431),
    .X(_01598_));
 sky130_fd_sc_hd__mux4_1 _28965_ (.A0(_02587_),
    .A1(_01593_),
    .A2(_01591_),
    .A3(_02587_),
    .S0(_14285_),
    .S1(net431),
    .X(_01594_));
 sky130_fd_sc_hd__mux4_1 _28966_ (.A0(_02586_),
    .A1(_01589_),
    .A2(_01587_),
    .A3(_02586_),
    .S0(_14285_),
    .S1(net431),
    .X(_01590_));
 sky130_fd_sc_hd__mux4_1 _28967_ (.A0(_02585_),
    .A1(_01585_),
    .A2(_01583_),
    .A3(_02585_),
    .S0(_14285_),
    .S1(net431),
    .X(_01586_));
 sky130_fd_sc_hd__mux4_1 _28968_ (.A0(_02584_),
    .A1(_01581_),
    .A2(_01579_),
    .A3(_02584_),
    .S0(_14285_),
    .S1(net431),
    .X(_01582_));
 sky130_fd_sc_hd__mux4_1 _28969_ (.A0(_02583_),
    .A1(_01577_),
    .A2(_01575_),
    .A3(_02583_),
    .S0(_14285_),
    .S1(net431),
    .X(_01578_));
 sky130_fd_sc_hd__mux4_1 _28970_ (.A0(_02582_),
    .A1(_01573_),
    .A2(_01571_),
    .A3(_02582_),
    .S0(_14285_),
    .S1(net431),
    .X(_01574_));
 sky130_fd_sc_hd__mux4_1 _28971_ (.A0(_02571_),
    .A1(_01569_),
    .A2(_01567_),
    .A3(_02571_),
    .S0(_14285_),
    .S1(net431),
    .X(_01570_));
 sky130_fd_sc_hd__dfxtp_1 _28972_ (.D(_02687_),
    .Q(\alu_shl[0] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _28973_ (.D(_02688_),
    .Q(\alu_shl[1] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _28974_ (.D(_02689_),
    .Q(\alu_shl[2] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _28975_ (.D(_02690_),
    .Q(\alu_shl[3] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _28976_ (.D(_02691_),
    .Q(\alu_shl[4] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _28977_ (.D(_02692_),
    .Q(\alu_shl[5] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _28978_ (.D(_02693_),
    .Q(\alu_shl[6] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _28979_ (.D(_02694_),
    .Q(\alu_shl[7] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _28980_ (.D(_02695_),
    .Q(\alu_shl[8] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _28981_ (.D(_02696_),
    .Q(\alu_shl[9] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _28982_ (.D(_02697_),
    .Q(\alu_shl[10] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _28983_ (.D(_02698_),
    .Q(\alu_shl[11] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _28984_ (.D(_02699_),
    .Q(\alu_shl[12] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _28985_ (.D(_02700_),
    .Q(\alu_shl[13] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _28986_ (.D(_02701_),
    .Q(\alu_shl[14] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _28987_ (.D(_02702_),
    .Q(\alu_shl[15] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _28988_ (.D(_02703_),
    .Q(alu_wait),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _28989_ (.D(_02704_),
    .Q(\latched_rd[3] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _28990_ (.D(_02705_),
    .Q(\latched_rd[2] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _28991_ (.D(_02706_),
    .Q(\latched_rd[1] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _28992_ (.D(_02707_),
    .Q(\latched_rd[0] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _28993_ (.D(_02708_),
    .Q(\decoded_imm[31] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _28994_ (.D(_02709_),
    .Q(\decoded_imm[30] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _28995_ (.D(_02710_),
    .Q(\decoded_imm[29] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _28996_ (.D(_02711_),
    .Q(\decoded_imm[28] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _28997_ (.D(_02712_),
    .Q(\decoded_imm[27] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _28998_ (.D(_02713_),
    .Q(\decoded_imm[26] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _28999_ (.D(_02714_),
    .Q(\decoded_imm[25] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29000_ (.D(_02715_),
    .Q(\decoded_imm[24] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _29001_ (.D(_02716_),
    .Q(\decoded_imm[23] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _29002_ (.D(_02717_),
    .Q(\decoded_imm[22] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _29003_ (.D(_02718_),
    .Q(\decoded_imm[21] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _29004_ (.D(_02719_),
    .Q(\decoded_imm[20] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _29005_ (.D(_02720_),
    .Q(\decoded_imm[19] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _29006_ (.D(_02721_),
    .Q(\decoded_imm[18] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29007_ (.D(_02722_),
    .Q(\decoded_imm[17] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _29008_ (.D(_02723_),
    .Q(\decoded_imm[16] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _29009_ (.D(_02724_),
    .Q(\decoded_imm[15] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29010_ (.D(_02725_),
    .Q(\decoded_imm[14] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29011_ (.D(_02726_),
    .Q(\decoded_imm[13] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29012_ (.D(_02727_),
    .Q(\decoded_imm[12] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29013_ (.D(_02728_),
    .Q(\decoded_imm[11] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29014_ (.D(_02729_),
    .Q(\decoded_imm[10] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29015_ (.D(_02730_),
    .Q(\decoded_imm[9] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29016_ (.D(_02731_),
    .Q(\decoded_imm[8] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29017_ (.D(_02732_),
    .Q(\decoded_imm[7] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29018_ (.D(_02733_),
    .Q(\decoded_imm[6] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29019_ (.D(_02734_),
    .Q(\decoded_imm[5] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29020_ (.D(_02735_),
    .Q(\decoded_imm[4] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29021_ (.D(_02736_),
    .Q(\decoded_imm[3] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29022_ (.D(_02737_),
    .Q(\decoded_imm[2] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _29023_ (.D(_02738_),
    .Q(\decoded_imm[1] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29024_ (.D(_02739_),
    .Q(\irq_pending[31] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29025_ (.D(_02740_),
    .Q(\irq_pending[30] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29026_ (.D(_02741_),
    .Q(\irq_pending[29] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29027_ (.D(_02742_),
    .Q(\irq_pending[28] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29028_ (.D(_02743_),
    .Q(\irq_pending[27] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29029_ (.D(_02744_),
    .Q(\irq_pending[26] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29030_ (.D(_02745_),
    .Q(\irq_pending[25] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29031_ (.D(_02746_),
    .Q(\irq_pending[24] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29032_ (.D(_02747_),
    .Q(\irq_pending[23] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _29033_ (.D(_02748_),
    .Q(\irq_pending[22] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _29034_ (.D(_02749_),
    .Q(\irq_pending[21] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _29035_ (.D(_02750_),
    .Q(\irq_pending[20] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _29036_ (.D(_02751_),
    .Q(\irq_pending[19] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _29037_ (.D(_02752_),
    .Q(\irq_pending[18] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _29038_ (.D(_02753_),
    .Q(\irq_pending[17] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _29039_ (.D(_02754_),
    .Q(\irq_pending[16] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _29040_ (.D(_02755_),
    .Q(\irq_pending[15] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _29041_ (.D(_02756_),
    .Q(\irq_pending[14] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _29042_ (.D(_02757_),
    .Q(\irq_pending[13] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _29043_ (.D(_02758_),
    .Q(\irq_pending[12] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _29044_ (.D(_02759_),
    .Q(\irq_pending[11] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _29045_ (.D(_02760_),
    .Q(\irq_pending[10] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _29046_ (.D(_02761_),
    .Q(\irq_pending[9] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _29047_ (.D(_02762_),
    .Q(\irq_pending[8] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _29048_ (.D(_02763_),
    .Q(\irq_pending[7] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _29049_ (.D(_02764_),
    .Q(\irq_pending[6] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _29050_ (.D(_02765_),
    .Q(\irq_pending[5] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _29051_ (.D(_02766_),
    .Q(\irq_pending[4] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _29052_ (.D(_02767_),
    .Q(\irq_pending[3] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _29053_ (.D(_02768_),
    .Q(\irq_pending[1] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _29054_ (.D(_02769_),
    .Q(\irq_pending[0] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29055_ (.D(_02770_),
    .Q(\reg_next_pc[0] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29056_ (.D(_00045_),
    .Q(\mem_wordsize[0] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _29057_ (.D(_00046_),
    .Q(\mem_wordsize[1] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _29058_ (.D(_00047_),
    .Q(\mem_wordsize[2] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29059_ (.D(_14287_),
    .Q(\reg_out[0] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29060_ (.D(_14298_),
    .Q(\reg_out[1] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29061_ (.D(_14309_),
    .Q(\reg_out[2] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29062_ (.D(_14312_),
    .Q(\reg_out[3] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29063_ (.D(_14313_),
    .Q(\reg_out[4] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29064_ (.D(_14314_),
    .Q(\reg_out[5] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29065_ (.D(_14315_),
    .Q(\reg_out[6] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29066_ (.D(_14316_),
    .Q(\reg_out[7] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29067_ (.D(_14317_),
    .Q(\reg_out[8] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29068_ (.D(_14318_),
    .Q(\reg_out[9] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29069_ (.D(_14288_),
    .Q(\reg_out[10] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29070_ (.D(_14289_),
    .Q(\reg_out[11] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29071_ (.D(_14290_),
    .Q(\reg_out[12] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29072_ (.D(_14291_),
    .Q(\reg_out[13] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29073_ (.D(_14292_),
    .Q(\reg_out[14] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29074_ (.D(_14293_),
    .Q(\reg_out[15] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29075_ (.D(_14294_),
    .Q(\reg_out[16] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29076_ (.D(_14295_),
    .Q(\reg_out[17] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29077_ (.D(_14296_),
    .Q(\reg_out[18] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29078_ (.D(_14297_),
    .Q(\reg_out[19] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29079_ (.D(_14299_),
    .Q(\reg_out[20] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29080_ (.D(_14300_),
    .Q(\reg_out[21] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29081_ (.D(_14301_),
    .Q(\reg_out[22] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29082_ (.D(_14302_),
    .Q(\reg_out[23] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29083_ (.D(_14303_),
    .Q(\reg_out[24] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29084_ (.D(_14304_),
    .Q(\reg_out[25] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29085_ (.D(_14305_),
    .Q(\reg_out[26] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29086_ (.D(_14306_),
    .Q(\reg_out[27] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29087_ (.D(_14307_),
    .Q(\reg_out[28] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29088_ (.D(_14308_),
    .Q(\reg_out[29] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29089_ (.D(_14310_),
    .Q(\reg_out[30] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29090_ (.D(_14311_),
    .Q(\reg_out[31] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _29091_ (.D(_00004_),
    .Q(\irq_pending[2] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _29092_ (.D(_00003_),
    .Q(decoder_trigger),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29093_ (.D(\alu_out[0] ),
    .Q(\alu_out_q[0] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29094_ (.D(\alu_out[1] ),
    .Q(\alu_out_q[1] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29095_ (.D(\alu_out[2] ),
    .Q(\alu_out_q[2] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29096_ (.D(\alu_out[3] ),
    .Q(\alu_out_q[3] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29097_ (.D(\alu_out[4] ),
    .Q(\alu_out_q[4] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29098_ (.D(\alu_out[5] ),
    .Q(\alu_out_q[5] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29099_ (.D(\alu_out[6] ),
    .Q(\alu_out_q[6] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29100_ (.D(\alu_out[7] ),
    .Q(\alu_out_q[7] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29101_ (.D(\alu_out[8] ),
    .Q(\alu_out_q[8] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29102_ (.D(\alu_out[9] ),
    .Q(\alu_out_q[9] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29103_ (.D(\alu_out[10] ),
    .Q(\alu_out_q[10] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29104_ (.D(\alu_out[11] ),
    .Q(\alu_out_q[11] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29105_ (.D(\alu_out[12] ),
    .Q(\alu_out_q[12] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29106_ (.D(\alu_out[13] ),
    .Q(\alu_out_q[13] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29107_ (.D(\alu_out[14] ),
    .Q(\alu_out_q[14] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29108_ (.D(\alu_out[15] ),
    .Q(\alu_out_q[15] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29109_ (.D(\alu_out[16] ),
    .Q(\alu_out_q[16] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29110_ (.D(\alu_out[17] ),
    .Q(\alu_out_q[17] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29111_ (.D(\alu_out[18] ),
    .Q(\alu_out_q[18] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29112_ (.D(\alu_out[19] ),
    .Q(\alu_out_q[19] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29113_ (.D(\alu_out[20] ),
    .Q(\alu_out_q[20] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29114_ (.D(\alu_out[21] ),
    .Q(\alu_out_q[21] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29115_ (.D(\alu_out[22] ),
    .Q(\alu_out_q[22] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29116_ (.D(\alu_out[23] ),
    .Q(\alu_out_q[23] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29117_ (.D(\alu_out[24] ),
    .Q(\alu_out_q[24] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29118_ (.D(\alu_out[25] ),
    .Q(\alu_out_q[25] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29119_ (.D(\alu_out[26] ),
    .Q(\alu_out_q[26] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29120_ (.D(\alu_out[27] ),
    .Q(\alu_out_q[27] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29121_ (.D(\alu_out[28] ),
    .Q(\alu_out_q[28] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29122_ (.D(\alu_out[29] ),
    .Q(\alu_out_q[29] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _29123_ (.D(\alu_out[30] ),
    .Q(\alu_out_q[30] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29124_ (.D(\alu_out[31] ),
    .Q(\alu_out_q[31] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _29125_ (.D(_00005_),
    .Q(is_lui_auipc_jal),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29126_ (.D(_00006_),
    .Q(is_slti_blt_slt),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29127_ (.D(_00007_),
    .Q(is_sltiu_bltu_sltu),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29128_ (.D(_02591_),
    .Q(\alu_add_sub[0] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29129_ (.D(_02602_),
    .Q(\alu_add_sub[1] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29130_ (.D(_02613_),
    .Q(\alu_add_sub[2] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29131_ (.D(_02616_),
    .Q(\alu_add_sub[3] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29132_ (.D(_02617_),
    .Q(\alu_add_sub[4] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29133_ (.D(_02618_),
    .Q(\alu_add_sub[5] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29134_ (.D(_02619_),
    .Q(\alu_add_sub[6] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29135_ (.D(_02620_),
    .Q(\alu_add_sub[7] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29136_ (.D(_02621_),
    .Q(\alu_add_sub[8] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29137_ (.D(_02622_),
    .Q(\alu_add_sub[9] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29138_ (.D(_02592_),
    .Q(\alu_add_sub[10] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29139_ (.D(_02593_),
    .Q(\alu_add_sub[11] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29140_ (.D(_02594_),
    .Q(\alu_add_sub[12] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29141_ (.D(_02595_),
    .Q(\alu_add_sub[13] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29142_ (.D(_02596_),
    .Q(\alu_add_sub[14] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29143_ (.D(_02597_),
    .Q(\alu_add_sub[15] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29144_ (.D(_02598_),
    .Q(\alu_add_sub[16] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29145_ (.D(_02599_),
    .Q(\alu_add_sub[17] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29146_ (.D(_02600_),
    .Q(\alu_add_sub[18] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29147_ (.D(_02601_),
    .Q(\alu_add_sub[19] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29148_ (.D(_02603_),
    .Q(\alu_add_sub[20] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29149_ (.D(_02604_),
    .Q(\alu_add_sub[21] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29150_ (.D(_02605_),
    .Q(\alu_add_sub[22] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29151_ (.D(_02606_),
    .Q(\alu_add_sub[23] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29152_ (.D(_02607_),
    .Q(\alu_add_sub[24] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29153_ (.D(_02608_),
    .Q(\alu_add_sub[25] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29154_ (.D(_02609_),
    .Q(\alu_add_sub[26] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29155_ (.D(_02610_),
    .Q(\alu_add_sub[27] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29156_ (.D(_02611_),
    .Q(\alu_add_sub[28] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29157_ (.D(_02612_),
    .Q(\alu_add_sub[29] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29158_ (.D(_02614_),
    .Q(\alu_add_sub[30] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29159_ (.D(_02615_),
    .Q(\alu_add_sub[31] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29160_ (.D(_14322_),
    .Q(\alu_shl[16] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29161_ (.D(_14323_),
    .Q(\alu_shl[17] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29162_ (.D(_14324_),
    .Q(\alu_shl[18] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29163_ (.D(_14325_),
    .Q(\alu_shl[19] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29164_ (.D(_14326_),
    .Q(\alu_shl[20] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29165_ (.D(_14327_),
    .Q(\alu_shl[21] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29166_ (.D(_14328_),
    .Q(\alu_shl[22] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29167_ (.D(_14329_),
    .Q(\alu_shl[23] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29168_ (.D(_14330_),
    .Q(\alu_shl[24] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29169_ (.D(_14331_),
    .Q(\alu_shl[25] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29170_ (.D(_14332_),
    .Q(\alu_shl[26] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29171_ (.D(_14333_),
    .Q(\alu_shl[27] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29172_ (.D(_14334_),
    .Q(\alu_shl[28] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29173_ (.D(_14335_),
    .Q(\alu_shl[29] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29174_ (.D(_14336_),
    .Q(\alu_shl[30] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29175_ (.D(_14337_),
    .Q(\alu_shl[31] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29176_ (.D(_14338_),
    .Q(\alu_shr[0] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29177_ (.D(_14349_),
    .Q(\alu_shr[1] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29178_ (.D(_14360_),
    .Q(\alu_shr[2] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29179_ (.D(_14363_),
    .Q(\alu_shr[3] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29180_ (.D(_14364_),
    .Q(\alu_shr[4] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29181_ (.D(_14365_),
    .Q(\alu_shr[5] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29182_ (.D(_14366_),
    .Q(\alu_shr[6] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29183_ (.D(_14367_),
    .Q(\alu_shr[7] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29184_ (.D(_14368_),
    .Q(\alu_shr[8] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29185_ (.D(_14369_),
    .Q(\alu_shr[9] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29186_ (.D(_14339_),
    .Q(\alu_shr[10] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29187_ (.D(_14340_),
    .Q(\alu_shr[11] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29188_ (.D(_14341_),
    .Q(\alu_shr[12] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29189_ (.D(_14342_),
    .Q(\alu_shr[13] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29190_ (.D(_14343_),
    .Q(\alu_shr[14] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29191_ (.D(_14344_),
    .Q(\alu_shr[15] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29192_ (.D(_14345_),
    .Q(\alu_shr[16] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29193_ (.D(_14346_),
    .Q(\alu_shr[17] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29194_ (.D(_14347_),
    .Q(\alu_shr[18] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29195_ (.D(_14348_),
    .Q(\alu_shr[19] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29196_ (.D(_14350_),
    .Q(\alu_shr[20] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29197_ (.D(_14351_),
    .Q(\alu_shr[21] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29198_ (.D(_14352_),
    .Q(\alu_shr[22] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29199_ (.D(_14353_),
    .Q(\alu_shr[23] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29200_ (.D(_14354_),
    .Q(\alu_shr[24] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29201_ (.D(_14355_),
    .Q(\alu_shr[25] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29202_ (.D(_14356_),
    .Q(\alu_shr[26] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29203_ (.D(_14357_),
    .Q(\alu_shr[27] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29204_ (.D(_14358_),
    .Q(\alu_shr[28] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29205_ (.D(_14359_),
    .Q(\alu_shr[29] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29206_ (.D(_14361_),
    .Q(\alu_shr[30] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29207_ (.D(_14362_),
    .Q(\alu_shr[31] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _29208_ (.D(_00000_),
    .Q(alu_eq),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _29209_ (.D(_00002_),
    .Q(alu_ltu),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _29210_ (.D(_00001_),
    .Q(alu_lts),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29211_ (.D(_02623_),
    .Q(\pcpi_mul.rd[0] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29212_ (.D(_02624_),
    .Q(\pcpi_mul.rd[1] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29213_ (.D(_02625_),
    .Q(\pcpi_mul.rd[2] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29214_ (.D(_02626_),
    .Q(\pcpi_mul.rd[3] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29215_ (.D(_02627_),
    .Q(\pcpi_mul.rd[4] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29216_ (.D(_02628_),
    .Q(\pcpi_mul.rd[5] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29217_ (.D(_02683_),
    .Q(\pcpi_mul.rd[6] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29218_ (.D(_02684_),
    .Q(\pcpi_mul.rd[7] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29219_ (.D(_02685_),
    .Q(\pcpi_mul.rd[8] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29220_ (.D(_02686_),
    .Q(\pcpi_mul.rd[9] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29221_ (.D(_02629_),
    .Q(\pcpi_mul.rd[10] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _29222_ (.D(_02630_),
    .Q(\pcpi_mul.rd[11] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _29223_ (.D(_02631_),
    .Q(\pcpi_mul.rd[12] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _29224_ (.D(_02632_),
    .Q(\pcpi_mul.rd[13] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _29225_ (.D(_02633_),
    .Q(\pcpi_mul.rd[14] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _29226_ (.D(_02634_),
    .Q(\pcpi_mul.rd[15] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29227_ (.D(_02635_),
    .Q(\pcpi_mul.rd[16] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _29228_ (.D(_02636_),
    .Q(\pcpi_mul.rd[17] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29229_ (.D(_02637_),
    .Q(\pcpi_mul.rd[18] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29230_ (.D(_02638_),
    .Q(\pcpi_mul.rd[19] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29231_ (.D(_02639_),
    .Q(\pcpi_mul.rd[20] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29232_ (.D(_02640_),
    .Q(\pcpi_mul.rd[21] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29233_ (.D(_02641_),
    .Q(\pcpi_mul.rd[22] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29234_ (.D(_02642_),
    .Q(\pcpi_mul.rd[23] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29235_ (.D(_02643_),
    .Q(\pcpi_mul.rd[24] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29236_ (.D(_02644_),
    .Q(\pcpi_mul.rd[25] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29237_ (.D(_02645_),
    .Q(\pcpi_mul.rd[26] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29238_ (.D(_02646_),
    .Q(\pcpi_mul.rd[27] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29239_ (.D(_02647_),
    .Q(\pcpi_mul.rd[28] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29240_ (.D(_02648_),
    .Q(\pcpi_mul.rd[29] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29241_ (.D(_02649_),
    .Q(\pcpi_mul.rd[30] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29242_ (.D(_02650_),
    .Q(\pcpi_mul.rd[31] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29243_ (.D(_02651_),
    .Q(\pcpi_mul.rd[32] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29244_ (.D(_02652_),
    .Q(\pcpi_mul.rd[33] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29245_ (.D(_02653_),
    .Q(\pcpi_mul.rd[34] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29246_ (.D(_02654_),
    .Q(\pcpi_mul.rd[35] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29247_ (.D(_02655_),
    .Q(\pcpi_mul.rd[36] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29248_ (.D(_02656_),
    .Q(\pcpi_mul.rd[37] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29249_ (.D(_02657_),
    .Q(\pcpi_mul.rd[38] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _29250_ (.D(_02658_),
    .Q(\pcpi_mul.rd[39] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29251_ (.D(_02659_),
    .Q(\pcpi_mul.rd[40] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _29252_ (.D(_02660_),
    .Q(\pcpi_mul.rd[41] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _29253_ (.D(_02661_),
    .Q(\pcpi_mul.rd[42] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _29254_ (.D(_02662_),
    .Q(\pcpi_mul.rd[43] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _29255_ (.D(_02663_),
    .Q(\pcpi_mul.rd[44] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _29256_ (.D(_02664_),
    .Q(\pcpi_mul.rd[45] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _29257_ (.D(_02665_),
    .Q(\pcpi_mul.rd[46] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _29258_ (.D(_02666_),
    .Q(\pcpi_mul.rd[47] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _29259_ (.D(_02667_),
    .Q(\pcpi_mul.rd[48] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _29260_ (.D(_02668_),
    .Q(\pcpi_mul.rd[49] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _29261_ (.D(_02669_),
    .Q(\pcpi_mul.rd[50] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _29262_ (.D(_02670_),
    .Q(\pcpi_mul.rd[51] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _29263_ (.D(_02671_),
    .Q(\pcpi_mul.rd[52] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _29264_ (.D(_02672_),
    .Q(\pcpi_mul.rd[53] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _29265_ (.D(_02673_),
    .Q(\pcpi_mul.rd[54] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _29266_ (.D(_02674_),
    .Q(\pcpi_mul.rd[55] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _29267_ (.D(_02675_),
    .Q(\pcpi_mul.rd[56] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _29268_ (.D(_02676_),
    .Q(\pcpi_mul.rd[57] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _29269_ (.D(_02677_),
    .Q(\pcpi_mul.rd[58] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _29270_ (.D(_02678_),
    .Q(\pcpi_mul.rd[59] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29271_ (.D(_02679_),
    .Q(\pcpi_mul.rd[60] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29272_ (.D(_02680_),
    .Q(\pcpi_mul.rd[61] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29273_ (.D(_02681_),
    .Q(\pcpi_mul.rd[62] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29274_ (.D(_02682_),
    .Q(\pcpi_mul.rd[63] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _29275_ (.D(\pcpi_mul.instr_any_mulh ),
    .Q(\pcpi_mul.shift_out ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29276_ (.D(_00038_),
    .Q(\cpu_state[0] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29277_ (.D(_00039_),
    .Q(\cpu_state[1] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _29278_ (.D(_00040_),
    .Q(\cpu_state[2] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _29279_ (.D(_00041_),
    .Q(\cpu_state[3] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29280_ (.D(_00042_),
    .Q(\cpu_state[4] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29281_ (.D(_00043_),
    .Q(\cpu_state[5] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29282_ (.D(_00044_),
    .Q(\cpu_state[6] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29283_ (.D(_02771_),
    .Q(\cpuregs[8][0] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29284_ (.D(_02772_),
    .Q(\cpuregs[8][1] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29285_ (.D(_02773_),
    .Q(\cpuregs[8][2] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29286_ (.D(_02774_),
    .Q(\cpuregs[8][3] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29287_ (.D(_02775_),
    .Q(\cpuregs[8][4] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29288_ (.D(_02776_),
    .Q(\cpuregs[8][5] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29289_ (.D(_02777_),
    .Q(\cpuregs[8][6] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29290_ (.D(_02778_),
    .Q(\cpuregs[8][7] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29291_ (.D(_02779_),
    .Q(\cpuregs[8][8] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29292_ (.D(_02780_),
    .Q(\cpuregs[8][9] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29293_ (.D(_02781_),
    .Q(\cpuregs[8][10] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29294_ (.D(_02782_),
    .Q(\cpuregs[8][11] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29295_ (.D(_02783_),
    .Q(\cpuregs[8][12] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29296_ (.D(_02784_),
    .Q(\cpuregs[8][13] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29297_ (.D(_02785_),
    .Q(\cpuregs[8][14] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29298_ (.D(_02786_),
    .Q(\cpuregs[8][15] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29299_ (.D(_02787_),
    .Q(\cpuregs[8][16] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29300_ (.D(_02788_),
    .Q(\cpuregs[8][17] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29301_ (.D(_02789_),
    .Q(\cpuregs[8][18] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29302_ (.D(_02790_),
    .Q(\cpuregs[8][19] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29303_ (.D(_02791_),
    .Q(\cpuregs[8][20] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29304_ (.D(_02792_),
    .Q(\cpuregs[8][21] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29305_ (.D(_02793_),
    .Q(\cpuregs[8][22] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29306_ (.D(_02794_),
    .Q(\cpuregs[8][23] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29307_ (.D(_02795_),
    .Q(\cpuregs[8][24] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29308_ (.D(_02796_),
    .Q(\cpuregs[8][25] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29309_ (.D(_02797_),
    .Q(\cpuregs[8][26] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29310_ (.D(_02798_),
    .Q(\cpuregs[8][27] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29311_ (.D(_02799_),
    .Q(\cpuregs[8][28] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29312_ (.D(_02800_),
    .Q(\cpuregs[8][29] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29313_ (.D(_02801_),
    .Q(\cpuregs[8][30] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29314_ (.D(_02802_),
    .Q(\cpuregs[8][31] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29315_ (.D(_02803_),
    .Q(\cpuregs[14][0] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29316_ (.D(_02804_),
    .Q(\cpuregs[14][1] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29317_ (.D(_02805_),
    .Q(\cpuregs[14][2] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29318_ (.D(_02806_),
    .Q(\cpuregs[14][3] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29319_ (.D(_02807_),
    .Q(\cpuregs[14][4] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29320_ (.D(_02808_),
    .Q(\cpuregs[14][5] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29321_ (.D(_02809_),
    .Q(\cpuregs[14][6] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29322_ (.D(_02810_),
    .Q(\cpuregs[14][7] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29323_ (.D(_02811_),
    .Q(\cpuregs[14][8] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29324_ (.D(_02812_),
    .Q(\cpuregs[14][9] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29325_ (.D(_02813_),
    .Q(\cpuregs[14][10] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29326_ (.D(_02814_),
    .Q(\cpuregs[14][11] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29327_ (.D(_02815_),
    .Q(\cpuregs[14][12] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29328_ (.D(_02816_),
    .Q(\cpuregs[14][13] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29329_ (.D(_02817_),
    .Q(\cpuregs[14][14] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29330_ (.D(_02818_),
    .Q(\cpuregs[14][15] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29331_ (.D(_02819_),
    .Q(\cpuregs[14][16] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29332_ (.D(_02820_),
    .Q(\cpuregs[14][17] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29333_ (.D(_02821_),
    .Q(\cpuregs[14][18] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29334_ (.D(_02822_),
    .Q(\cpuregs[14][19] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29335_ (.D(_02823_),
    .Q(\cpuregs[14][20] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29336_ (.D(_02824_),
    .Q(\cpuregs[14][21] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29337_ (.D(_02825_),
    .Q(\cpuregs[14][22] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29338_ (.D(_02826_),
    .Q(\cpuregs[14][23] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29339_ (.D(_02827_),
    .Q(\cpuregs[14][24] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29340_ (.D(_02828_),
    .Q(\cpuregs[14][25] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29341_ (.D(_02829_),
    .Q(\cpuregs[14][26] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29342_ (.D(_02830_),
    .Q(\cpuregs[14][27] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29343_ (.D(_02831_),
    .Q(\cpuregs[14][28] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29344_ (.D(_02832_),
    .Q(\cpuregs[14][29] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29345_ (.D(_02833_),
    .Q(\cpuregs[14][30] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29346_ (.D(_02834_),
    .Q(\cpuregs[14][31] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29347_ (.D(_02835_),
    .Q(\cpuregs[0][0] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29348_ (.D(_02836_),
    .Q(\cpuregs[0][1] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29349_ (.D(_02837_),
    .Q(\cpuregs[0][2] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29350_ (.D(_02838_),
    .Q(\cpuregs[0][3] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29351_ (.D(_02839_),
    .Q(\cpuregs[0][4] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29352_ (.D(_02840_),
    .Q(\cpuregs[0][5] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29353_ (.D(_02841_),
    .Q(\cpuregs[0][6] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29354_ (.D(_02842_),
    .Q(\cpuregs[0][7] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29355_ (.D(_02843_),
    .Q(\cpuregs[0][8] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29356_ (.D(_02844_),
    .Q(\cpuregs[0][9] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29357_ (.D(_02845_),
    .Q(\cpuregs[0][10] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29358_ (.D(_02846_),
    .Q(\cpuregs[0][11] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29359_ (.D(_02847_),
    .Q(\cpuregs[0][12] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29360_ (.D(_02848_),
    .Q(\cpuregs[0][13] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29361_ (.D(_02849_),
    .Q(\cpuregs[0][14] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29362_ (.D(_02850_),
    .Q(\cpuregs[0][15] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29363_ (.D(_02851_),
    .Q(\cpuregs[0][16] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29364_ (.D(_02852_),
    .Q(\cpuregs[0][17] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29365_ (.D(_02853_),
    .Q(\cpuregs[0][18] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29366_ (.D(_02854_),
    .Q(\cpuregs[0][19] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29367_ (.D(_02855_),
    .Q(\cpuregs[0][20] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29368_ (.D(_02856_),
    .Q(\cpuregs[0][21] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29369_ (.D(_02857_),
    .Q(\cpuregs[0][22] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29370_ (.D(_02858_),
    .Q(\cpuregs[0][23] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29371_ (.D(_02859_),
    .Q(\cpuregs[0][24] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29372_ (.D(_02860_),
    .Q(\cpuregs[0][25] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29373_ (.D(_02861_),
    .Q(\cpuregs[0][26] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29374_ (.D(_02862_),
    .Q(\cpuregs[0][27] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29375_ (.D(_02863_),
    .Q(\cpuregs[0][28] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29376_ (.D(_02864_),
    .Q(\cpuregs[0][29] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29377_ (.D(_02865_),
    .Q(\cpuregs[0][30] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29378_ (.D(_02866_),
    .Q(\cpuregs[0][31] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29379_ (.D(_02867_),
    .Q(\cpuregs[10][0] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29380_ (.D(_02868_),
    .Q(\cpuregs[10][1] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29381_ (.D(_02869_),
    .Q(\cpuregs[10][2] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29382_ (.D(_02870_),
    .Q(\cpuregs[10][3] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29383_ (.D(_02871_),
    .Q(\cpuregs[10][4] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29384_ (.D(_02872_),
    .Q(\cpuregs[10][5] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29385_ (.D(_02873_),
    .Q(\cpuregs[10][6] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29386_ (.D(_02874_),
    .Q(\cpuregs[10][7] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29387_ (.D(_02875_),
    .Q(\cpuregs[10][8] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29388_ (.D(_02876_),
    .Q(\cpuregs[10][9] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29389_ (.D(_02877_),
    .Q(\cpuregs[10][10] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29390_ (.D(_02878_),
    .Q(\cpuregs[10][11] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29391_ (.D(_02879_),
    .Q(\cpuregs[10][12] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29392_ (.D(_02880_),
    .Q(\cpuregs[10][13] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29393_ (.D(_02881_),
    .Q(\cpuregs[10][14] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29394_ (.D(_02882_),
    .Q(\cpuregs[10][15] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29395_ (.D(_02883_),
    .Q(\cpuregs[10][16] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29396_ (.D(_02884_),
    .Q(\cpuregs[10][17] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29397_ (.D(_02885_),
    .Q(\cpuregs[10][18] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29398_ (.D(_02886_),
    .Q(\cpuregs[10][19] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29399_ (.D(_02887_),
    .Q(\cpuregs[10][20] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29400_ (.D(_02888_),
    .Q(\cpuregs[10][21] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29401_ (.D(_02889_),
    .Q(\cpuregs[10][22] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29402_ (.D(_02890_),
    .Q(\cpuregs[10][23] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29403_ (.D(_02891_),
    .Q(\cpuregs[10][24] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29404_ (.D(_02892_),
    .Q(\cpuregs[10][25] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29405_ (.D(_02893_),
    .Q(\cpuregs[10][26] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29406_ (.D(_02894_),
    .Q(\cpuregs[10][27] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29407_ (.D(_02895_),
    .Q(\cpuregs[10][28] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29408_ (.D(_02896_),
    .Q(\cpuregs[10][29] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29409_ (.D(_02897_),
    .Q(\cpuregs[10][30] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29410_ (.D(_02898_),
    .Q(\cpuregs[10][31] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29411_ (.D(_02899_),
    .Q(\cpuregs[18][0] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29412_ (.D(_02900_),
    .Q(\cpuregs[18][1] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29413_ (.D(_02901_),
    .Q(\cpuregs[18][2] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29414_ (.D(_02902_),
    .Q(\cpuregs[18][3] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29415_ (.D(_02903_),
    .Q(\cpuregs[18][4] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29416_ (.D(_02904_),
    .Q(\cpuregs[18][5] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29417_ (.D(_02905_),
    .Q(\cpuregs[18][6] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29418_ (.D(_02906_),
    .Q(\cpuregs[18][7] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29419_ (.D(_02907_),
    .Q(\cpuregs[18][8] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29420_ (.D(_02908_),
    .Q(\cpuregs[18][9] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29421_ (.D(_02909_),
    .Q(\cpuregs[18][10] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29422_ (.D(_02910_),
    .Q(\cpuregs[18][11] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29423_ (.D(_02911_),
    .Q(\cpuregs[18][12] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29424_ (.D(_02912_),
    .Q(\cpuregs[18][13] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29425_ (.D(_02913_),
    .Q(\cpuregs[18][14] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29426_ (.D(_02914_),
    .Q(\cpuregs[18][15] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29427_ (.D(_02915_),
    .Q(\cpuregs[18][16] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29428_ (.D(_02916_),
    .Q(\cpuregs[18][17] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29429_ (.D(_02917_),
    .Q(\cpuregs[18][18] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29430_ (.D(_02918_),
    .Q(\cpuregs[18][19] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29431_ (.D(_02919_),
    .Q(\cpuregs[18][20] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29432_ (.D(_02920_),
    .Q(\cpuregs[18][21] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29433_ (.D(_02921_),
    .Q(\cpuregs[18][22] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29434_ (.D(_02922_),
    .Q(\cpuregs[18][23] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29435_ (.D(_02923_),
    .Q(\cpuregs[18][24] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29436_ (.D(_02924_),
    .Q(\cpuregs[18][25] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29437_ (.D(_02925_),
    .Q(\cpuregs[18][26] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29438_ (.D(_02926_),
    .Q(\cpuregs[18][27] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29439_ (.D(_02927_),
    .Q(\cpuregs[18][28] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29440_ (.D(_02928_),
    .Q(\cpuregs[18][29] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29441_ (.D(_02929_),
    .Q(\cpuregs[18][30] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29442_ (.D(_02930_),
    .Q(\cpuregs[18][31] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29443_ (.D(_02931_),
    .Q(\mem_rdata_q[0] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29444_ (.D(_02932_),
    .Q(\mem_rdata_q[1] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29445_ (.D(_02933_),
    .Q(\mem_rdata_q[2] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29446_ (.D(_02934_),
    .Q(\mem_rdata_q[3] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29447_ (.D(_02935_),
    .Q(\mem_rdata_q[4] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29448_ (.D(_02936_),
    .Q(\mem_rdata_q[5] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29449_ (.D(_02937_),
    .Q(\mem_rdata_q[6] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _29450_ (.D(_02938_),
    .Q(\mem_rdata_q[7] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _29451_ (.D(_02939_),
    .Q(\mem_rdata_q[8] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _29452_ (.D(_02940_),
    .Q(\mem_rdata_q[9] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _29453_ (.D(_02941_),
    .Q(\mem_rdata_q[10] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _29454_ (.D(_02942_),
    .Q(\mem_rdata_q[11] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29455_ (.D(_02943_),
    .Q(\mem_rdata_q[12] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29456_ (.D(_02944_),
    .Q(\mem_rdata_q[13] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29457_ (.D(_02945_),
    .Q(\mem_rdata_q[14] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _29458_ (.D(_02946_),
    .Q(\mem_rdata_q[15] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _29459_ (.D(_02947_),
    .Q(\mem_rdata_q[16] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _29460_ (.D(_02948_),
    .Q(\mem_rdata_q[17] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _29461_ (.D(_02949_),
    .Q(\mem_rdata_q[18] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _29462_ (.D(_02950_),
    .Q(\mem_rdata_q[19] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _29463_ (.D(_02951_),
    .Q(\mem_rdata_q[20] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29464_ (.D(_02952_),
    .Q(\mem_rdata_q[21] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _29465_ (.D(_02953_),
    .Q(\mem_rdata_q[22] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _29466_ (.D(_02954_),
    .Q(\mem_rdata_q[23] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29467_ (.D(_02955_),
    .Q(\mem_rdata_q[24] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29468_ (.D(_02956_),
    .Q(\mem_rdata_q[25] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29469_ (.D(_02957_),
    .Q(\mem_rdata_q[26] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29470_ (.D(_02958_),
    .Q(\mem_rdata_q[27] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29471_ (.D(_02959_),
    .Q(\mem_rdata_q[28] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29472_ (.D(_02960_),
    .Q(\mem_rdata_q[29] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29473_ (.D(_02961_),
    .Q(\mem_rdata_q[30] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29474_ (.D(_02962_),
    .Q(\mem_rdata_q[31] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29475_ (.D(_02963_),
    .Q(\cpuregs[2][0] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29476_ (.D(_02964_),
    .Q(\cpuregs[2][1] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29477_ (.D(_02965_),
    .Q(\cpuregs[2][2] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29478_ (.D(_02966_),
    .Q(\cpuregs[2][3] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29479_ (.D(_02967_),
    .Q(\cpuregs[2][4] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29480_ (.D(_02968_),
    .Q(\cpuregs[2][5] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29481_ (.D(_02969_),
    .Q(\cpuregs[2][6] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29482_ (.D(_02970_),
    .Q(\cpuregs[2][7] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29483_ (.D(_02971_),
    .Q(\cpuregs[2][8] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29484_ (.D(_02972_),
    .Q(\cpuregs[2][9] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29485_ (.D(_02973_),
    .Q(\cpuregs[2][10] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29486_ (.D(_02974_),
    .Q(\cpuregs[2][11] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29487_ (.D(_02975_),
    .Q(\cpuregs[2][12] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29488_ (.D(_02976_),
    .Q(\cpuregs[2][13] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29489_ (.D(_02977_),
    .Q(\cpuregs[2][14] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29490_ (.D(_02978_),
    .Q(\cpuregs[2][15] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29491_ (.D(_02979_),
    .Q(\cpuregs[2][16] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29492_ (.D(_02980_),
    .Q(\cpuregs[2][17] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29493_ (.D(_02981_),
    .Q(\cpuregs[2][18] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29494_ (.D(_02982_),
    .Q(\cpuregs[2][19] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29495_ (.D(_02983_),
    .Q(\cpuregs[2][20] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29496_ (.D(_02984_),
    .Q(\cpuregs[2][21] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29497_ (.D(_02985_),
    .Q(\cpuregs[2][22] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29498_ (.D(_02986_),
    .Q(\cpuregs[2][23] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29499_ (.D(_02987_),
    .Q(\cpuregs[2][24] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29500_ (.D(_02988_),
    .Q(\cpuregs[2][25] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29501_ (.D(_02989_),
    .Q(\cpuregs[2][26] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29502_ (.D(_02990_),
    .Q(\cpuregs[2][27] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29503_ (.D(_02991_),
    .Q(\cpuregs[2][28] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29504_ (.D(_02992_),
    .Q(\cpuregs[2][29] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29505_ (.D(_02993_),
    .Q(\cpuregs[2][30] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29506_ (.D(_02994_),
    .Q(\cpuregs[2][31] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29507_ (.D(_02995_),
    .Q(\cpuregs[5][0] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29508_ (.D(_02996_),
    .Q(\cpuregs[5][1] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29509_ (.D(_02997_),
    .Q(\cpuregs[5][2] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29510_ (.D(_02998_),
    .Q(\cpuregs[5][3] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29511_ (.D(_02999_),
    .Q(\cpuregs[5][4] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29512_ (.D(_03000_),
    .Q(\cpuregs[5][5] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29513_ (.D(_03001_),
    .Q(\cpuregs[5][6] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29514_ (.D(_03002_),
    .Q(\cpuregs[5][7] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29515_ (.D(_03003_),
    .Q(\cpuregs[5][8] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29516_ (.D(_03004_),
    .Q(\cpuregs[5][9] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29517_ (.D(_03005_),
    .Q(\cpuregs[5][10] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29518_ (.D(_03006_),
    .Q(\cpuregs[5][11] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29519_ (.D(_03007_),
    .Q(\cpuregs[5][12] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29520_ (.D(_03008_),
    .Q(\cpuregs[5][13] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29521_ (.D(_03009_),
    .Q(\cpuregs[5][14] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29522_ (.D(_03010_),
    .Q(\cpuregs[5][15] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29523_ (.D(_03011_),
    .Q(\cpuregs[5][16] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29524_ (.D(_03012_),
    .Q(\cpuregs[5][17] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29525_ (.D(_03013_),
    .Q(\cpuregs[5][18] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29526_ (.D(_03014_),
    .Q(\cpuregs[5][19] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29527_ (.D(_03015_),
    .Q(\cpuregs[5][20] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29528_ (.D(_03016_),
    .Q(\cpuregs[5][21] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29529_ (.D(_03017_),
    .Q(\cpuregs[5][22] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29530_ (.D(_03018_),
    .Q(\cpuregs[5][23] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29531_ (.D(_03019_),
    .Q(\cpuregs[5][24] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29532_ (.D(_03020_),
    .Q(\cpuregs[5][25] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29533_ (.D(_03021_),
    .Q(\cpuregs[5][26] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29534_ (.D(_03022_),
    .Q(\cpuregs[5][27] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29535_ (.D(_03023_),
    .Q(\cpuregs[5][28] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29536_ (.D(_03024_),
    .Q(\cpuregs[5][29] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29537_ (.D(_03025_),
    .Q(\cpuregs[5][30] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29538_ (.D(_03026_),
    .Q(\cpuregs[5][31] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29539_ (.D(_03027_),
    .Q(\pcpi_mul.rs1[0] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29540_ (.D(_03028_),
    .Q(\pcpi_mul.rs1[1] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29541_ (.D(_03029_),
    .Q(\pcpi_mul.rs1[2] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29542_ (.D(_03030_),
    .Q(\pcpi_mul.rs1[3] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29543_ (.D(_03031_),
    .Q(\pcpi_mul.rs1[4] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29544_ (.D(_03032_),
    .Q(\pcpi_mul.rs1[5] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29545_ (.D(_03033_),
    .Q(\pcpi_mul.rs1[6] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29546_ (.D(_03034_),
    .Q(\pcpi_mul.rs1[7] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29547_ (.D(_03035_),
    .Q(\pcpi_mul.rs1[8] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29548_ (.D(_03036_),
    .Q(\pcpi_mul.rs1[9] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29549_ (.D(_03037_),
    .Q(\pcpi_mul.rs1[10] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _29550_ (.D(_03038_),
    .Q(\pcpi_mul.rs1[11] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29551_ (.D(_03039_),
    .Q(\pcpi_mul.rs1[12] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29552_ (.D(_03040_),
    .Q(\pcpi_mul.rs1[13] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29553_ (.D(_03041_),
    .Q(\pcpi_mul.rs1[14] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29554_ (.D(_03042_),
    .Q(\pcpi_mul.rs1[15] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29555_ (.D(_03043_),
    .Q(\pcpi_mul.rs1[16] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29556_ (.D(_03044_),
    .Q(\pcpi_mul.rs1[17] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29557_ (.D(_03045_),
    .Q(\pcpi_mul.rs1[18] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29558_ (.D(_03046_),
    .Q(\pcpi_mul.rs1[19] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29559_ (.D(_03047_),
    .Q(\pcpi_mul.rs1[20] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29560_ (.D(_03048_),
    .Q(\pcpi_mul.rs1[21] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29561_ (.D(_03049_),
    .Q(\pcpi_mul.rs1[22] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29562_ (.D(_03050_),
    .Q(\pcpi_mul.rs1[23] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29563_ (.D(_03051_),
    .Q(\pcpi_mul.rs1[24] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29564_ (.D(_03052_),
    .Q(\pcpi_mul.rs1[25] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29565_ (.D(_03053_),
    .Q(\pcpi_mul.rs1[26] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29566_ (.D(_03054_),
    .Q(\pcpi_mul.rs1[27] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29567_ (.D(_03055_),
    .Q(\pcpi_mul.rs1[28] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _29568_ (.D(_03056_),
    .Q(\pcpi_mul.rs1[29] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _29569_ (.D(_03057_),
    .Q(\pcpi_mul.rs1[30] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29570_ (.D(_03058_),
    .Q(\pcpi_mul.rs1[31] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _29571_ (.D(_03059_),
    .Q(net156),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _29572_ (.D(_03060_),
    .Q(net159),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _29573_ (.D(_03061_),
    .Q(net160),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _29574_ (.D(_03062_),
    .Q(net161),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _29575_ (.D(_03063_),
    .Q(net162),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _29576_ (.D(_03064_),
    .Q(net163),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29577_ (.D(_03065_),
    .Q(net164),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _29578_ (.D(_03066_),
    .Q(net165),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _29579_ (.D(_03067_),
    .Q(net135),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _29580_ (.D(_03068_),
    .Q(net136),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _29581_ (.D(_03069_),
    .Q(net137),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _29582_ (.D(_03070_),
    .Q(net138),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _29583_ (.D(_03071_),
    .Q(net139),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29584_ (.D(_03072_),
    .Q(net140),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _29585_ (.D(_03073_),
    .Q(net141),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _29586_ (.D(_03074_),
    .Q(net142),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _29587_ (.D(_03075_),
    .Q(net143),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _29588_ (.D(_03076_),
    .Q(net144),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _29589_ (.D(_03077_),
    .Q(net146),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _29590_ (.D(_03078_),
    .Q(net147),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _29591_ (.D(_03079_),
    .Q(net148),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _29592_ (.D(_03080_),
    .Q(net149),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _29593_ (.D(_03081_),
    .Q(net150),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _29594_ (.D(_03082_),
    .Q(net151),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _29595_ (.D(_03083_),
    .Q(net152),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _29596_ (.D(_03084_),
    .Q(net153),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _29597_ (.D(_03085_),
    .Q(net154),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _29598_ (.D(_03086_),
    .Q(net155),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29599_ (.D(_03087_),
    .Q(net157),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _29600_ (.D(_03088_),
    .Q(net158),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _29601_ (.D(_03089_),
    .Q(net306),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _29602_ (.D(_03090_),
    .Q(net317),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _29603_ (.D(_03091_),
    .Q(net328),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _29604_ (.D(_03092_),
    .Q(net331),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _29605_ (.D(_03093_),
    .Q(net332),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _29606_ (.D(_03094_),
    .Q(net333),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _29607_ (.D(_03095_),
    .Q(net334),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _29608_ (.D(_03096_),
    .Q(net335),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _29609_ (.D(_03097_),
    .Q(net336),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _29610_ (.D(_03098_),
    .Q(net337),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _29611_ (.D(_03099_),
    .Q(net307),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _29612_ (.D(_03100_),
    .Q(net308),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _29613_ (.D(_03101_),
    .Q(net309),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _29614_ (.D(_03102_),
    .Q(net310),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _29615_ (.D(_03103_),
    .Q(net311),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _29616_ (.D(_03104_),
    .Q(net312),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _29617_ (.D(_03105_),
    .Q(net313),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _29618_ (.D(_03106_),
    .Q(net314),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _29619_ (.D(_03107_),
    .Q(net315),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _29620_ (.D(_03108_),
    .Q(net316),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _29621_ (.D(_03109_),
    .Q(net318),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _29622_ (.D(_03110_),
    .Q(net319),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _29623_ (.D(_03111_),
    .Q(net320),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _29624_ (.D(_03112_),
    .Q(net321),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _29625_ (.D(_03113_),
    .Q(net322),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _29626_ (.D(_03114_),
    .Q(net323),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _29627_ (.D(_03115_),
    .Q(net324),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _29628_ (.D(_03116_),
    .Q(net325),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _29629_ (.D(_03117_),
    .Q(net326),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _29630_ (.D(_03118_),
    .Q(net327),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _29631_ (.D(_03119_),
    .Q(net329),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _29632_ (.D(_03120_),
    .Q(net330),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _29633_ (.D(_03121_),
    .Q(net274),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _29634_ (.D(_03122_),
    .Q(net285),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _29635_ (.D(_03123_),
    .Q(net296),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _29636_ (.D(_03124_),
    .Q(net299),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _29637_ (.D(_03125_),
    .Q(net300),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _29638_ (.D(_03126_),
    .Q(net301),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _29639_ (.D(_03127_),
    .Q(net302),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _29640_ (.D(_03128_),
    .Q(net303),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _29641_ (.D(_03129_),
    .Q(net304),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _29642_ (.D(_03130_),
    .Q(net305),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _29643_ (.D(_03131_),
    .Q(net275),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _29644_ (.D(_03132_),
    .Q(net276),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _29645_ (.D(_03133_),
    .Q(net277),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _29646_ (.D(_03134_),
    .Q(net278),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _29647_ (.D(_03135_),
    .Q(net279),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _29648_ (.D(_03136_),
    .Q(net280),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _29649_ (.D(_03137_),
    .Q(net281),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _29650_ (.D(_03138_),
    .Q(net282),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _29651_ (.D(_03139_),
    .Q(net283),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _29652_ (.D(_03140_),
    .Q(net284),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _29653_ (.D(_03141_),
    .Q(net286),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _29654_ (.D(_03142_),
    .Q(net287),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _29655_ (.D(_03143_),
    .Q(net288),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _29656_ (.D(_03144_),
    .Q(net289),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _29657_ (.D(_03145_),
    .Q(net290),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _29658_ (.D(_03146_),
    .Q(net291),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _29659_ (.D(_03147_),
    .Q(net292),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _29660_ (.D(_03148_),
    .Q(net293),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _29661_ (.D(_03149_),
    .Q(net294),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _29662_ (.D(_03150_),
    .Q(net295),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _29663_ (.D(_03151_),
    .Q(net297),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _29664_ (.D(_03152_),
    .Q(net298),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29665_ (.D(_03153_),
    .Q(instr_lui),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29666_ (.D(_03154_),
    .Q(instr_auipc),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _29667_ (.D(_03155_),
    .Q(instr_jal),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29668_ (.D(_03156_),
    .Q(instr_jalr),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29669_ (.D(_03157_),
    .Q(instr_lb),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29670_ (.D(_03158_),
    .Q(instr_lh),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29671_ (.D(_03159_),
    .Q(instr_lw),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29672_ (.D(_03160_),
    .Q(instr_lbu),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29673_ (.D(_03161_),
    .Q(instr_lhu),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29674_ (.D(_03162_),
    .Q(instr_sb),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29675_ (.D(_03163_),
    .Q(instr_sh),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29676_ (.D(_03164_),
    .Q(instr_sw),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29677_ (.D(_03165_),
    .Q(instr_slli),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29678_ (.D(_03166_),
    .Q(instr_srli),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _29679_ (.D(_03167_),
    .Q(instr_srai),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29680_ (.D(_03168_),
    .Q(instr_rdcycle),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29681_ (.D(_03169_),
    .Q(instr_rdcycleh),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29682_ (.D(_03170_),
    .Q(instr_rdinstr),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29683_ (.D(_03171_),
    .Q(instr_rdinstrh),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _29684_ (.D(_03172_),
    .Q(instr_ecall_ebreak),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29685_ (.D(_03173_),
    .Q(instr_getq),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29686_ (.D(_03174_),
    .Q(instr_setq),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29687_ (.D(_03175_),
    .Q(instr_retirq),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _29688_ (.D(_03176_),
    .Q(instr_maskirq),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _29689_ (.D(_03177_),
    .Q(instr_waitirq),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _29690_ (.D(_03178_),
    .Q(instr_timer),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29691_ (.D(_03179_),
    .Q(\decoded_rd[0] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _29692_ (.D(_03180_),
    .Q(\decoded_rd[1] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _29693_ (.D(_03181_),
    .Q(\decoded_rd[2] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _29694_ (.D(_03182_),
    .Q(\decoded_rd[3] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29695_ (.D(_03183_),
    .Q(\decoded_rd[4] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29696_ (.D(_03184_),
    .Q(\decoded_imm[0] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _29697_ (.D(_03185_),
    .Q(\decoded_imm_uj[1] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _29698_ (.D(_03186_),
    .Q(\decoded_imm_uj[2] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _29699_ (.D(_03187_),
    .Q(\decoded_imm_uj[3] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _29700_ (.D(_03188_),
    .Q(\decoded_imm_uj[4] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29701_ (.D(_03189_),
    .Q(\decoded_imm_uj[5] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29702_ (.D(_03190_),
    .Q(\decoded_imm_uj[6] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29703_ (.D(_03191_),
    .Q(\decoded_imm_uj[7] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29704_ (.D(_03192_),
    .Q(\decoded_imm_uj[8] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29705_ (.D(_03193_),
    .Q(\decoded_imm_uj[9] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29706_ (.D(_03194_),
    .Q(\decoded_imm_uj[10] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _29707_ (.D(_03195_),
    .Q(\decoded_imm_uj[11] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29708_ (.D(_03196_),
    .Q(\decoded_imm_uj[12] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29709_ (.D(_03197_),
    .Q(\decoded_imm_uj[13] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _29710_ (.D(_03198_),
    .Q(\decoded_imm_uj[14] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29711_ (.D(_03199_),
    .Q(\decoded_imm_uj[15] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _29712_ (.D(_03200_),
    .Q(\decoded_imm_uj[16] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _29713_ (.D(_03201_),
    .Q(\decoded_imm_uj[17] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _29714_ (.D(_03202_),
    .Q(\decoded_imm_uj[18] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _29715_ (.D(_03203_),
    .Q(\decoded_imm_uj[19] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29716_ (.D(_03204_),
    .Q(\decoded_imm_uj[20] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29717_ (.D(_03205_),
    .Q(is_lb_lh_lw_lbu_lhu),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _29718_ (.D(_03206_),
    .Q(is_slli_srli_srai),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _29719_ (.D(_03207_),
    .Q(is_jalr_addi_slti_sltiu_xori_ori_andi),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _29720_ (.D(_03208_),
    .Q(is_sb_sh_sw),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29721_ (.D(_03209_),
    .Q(\cpuregs[13][0] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29722_ (.D(_03210_),
    .Q(\cpuregs[13][1] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29723_ (.D(_03211_),
    .Q(\cpuregs[13][2] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29724_ (.D(_03212_),
    .Q(\cpuregs[13][3] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29725_ (.D(_03213_),
    .Q(\cpuregs[13][4] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29726_ (.D(_03214_),
    .Q(\cpuregs[13][5] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29727_ (.D(_03215_),
    .Q(\cpuregs[13][6] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29728_ (.D(_03216_),
    .Q(\cpuregs[13][7] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29729_ (.D(_03217_),
    .Q(\cpuregs[13][8] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29730_ (.D(_03218_),
    .Q(\cpuregs[13][9] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29731_ (.D(_03219_),
    .Q(\cpuregs[13][10] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29732_ (.D(_03220_),
    .Q(\cpuregs[13][11] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29733_ (.D(_03221_),
    .Q(\cpuregs[13][12] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29734_ (.D(_03222_),
    .Q(\cpuregs[13][13] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29735_ (.D(_03223_),
    .Q(\cpuregs[13][14] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29736_ (.D(_03224_),
    .Q(\cpuregs[13][15] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29737_ (.D(_03225_),
    .Q(\cpuregs[13][16] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29738_ (.D(_03226_),
    .Q(\cpuregs[13][17] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29739_ (.D(_03227_),
    .Q(\cpuregs[13][18] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29740_ (.D(_03228_),
    .Q(\cpuregs[13][19] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29741_ (.D(_03229_),
    .Q(\cpuregs[13][20] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29742_ (.D(_03230_),
    .Q(\cpuregs[13][21] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29743_ (.D(_03231_),
    .Q(\cpuregs[13][22] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29744_ (.D(_03232_),
    .Q(\cpuregs[13][23] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29745_ (.D(_03233_),
    .Q(\cpuregs[13][24] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29746_ (.D(_03234_),
    .Q(\cpuregs[13][25] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29747_ (.D(_03235_),
    .Q(\cpuregs[13][26] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29748_ (.D(_03236_),
    .Q(\cpuregs[13][27] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29749_ (.D(_03237_),
    .Q(\cpuregs[13][28] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29750_ (.D(_03238_),
    .Q(\cpuregs[13][29] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29751_ (.D(_03239_),
    .Q(\cpuregs[13][30] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29752_ (.D(_03240_),
    .Q(\cpuregs[13][31] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29753_ (.D(_03241_),
    .Q(is_alu_reg_imm),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29754_ (.D(_03242_),
    .Q(is_alu_reg_reg),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _29755_ (.D(_03243_),
    .Q(net270),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _29756_ (.D(_03244_),
    .Q(net271),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _29757_ (.D(_03245_),
    .Q(net272),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _29758_ (.D(_03246_),
    .Q(net273),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _29759_ (.D(_03247_),
    .Q(\pcpi_mul.rs2[0] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29760_ (.D(_03248_),
    .Q(\pcpi_mul.rs2[1] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29761_ (.D(_03249_),
    .Q(\pcpi_mul.rs2[2] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _29762_ (.D(_03250_),
    .Q(\pcpi_mul.rs2[3] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29763_ (.D(_03251_),
    .Q(\pcpi_mul.rs2[4] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29764_ (.D(_03252_),
    .Q(\pcpi_mul.rs2[5] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _29765_ (.D(_03253_),
    .Q(\pcpi_mul.rs2[6] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29766_ (.D(_03254_),
    .Q(\pcpi_mul.rs2[7] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29767_ (.D(_03255_),
    .Q(\pcpi_mul.rs2[8] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _29768_ (.D(_03256_),
    .Q(\pcpi_mul.rs2[9] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29769_ (.D(_03257_),
    .Q(\pcpi_mul.rs2[10] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _29770_ (.D(_03258_),
    .Q(\pcpi_mul.rs2[11] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _29771_ (.D(_03259_),
    .Q(\pcpi_mul.rs2[12] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29772_ (.D(_03260_),
    .Q(\pcpi_mul.rs2[13] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29773_ (.D(_03261_),
    .Q(\pcpi_mul.rs2[14] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29774_ (.D(_03262_),
    .Q(\pcpi_mul.rs2[15] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _29775_ (.D(_03263_),
    .Q(\pcpi_mul.rs2[16] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _29776_ (.D(_03264_),
    .Q(\pcpi_mul.rs2[17] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _29777_ (.D(_03265_),
    .Q(\pcpi_mul.rs2[18] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _29778_ (.D(_03266_),
    .Q(\pcpi_mul.rs2[19] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _29779_ (.D(_03267_),
    .Q(\pcpi_mul.rs2[20] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _29780_ (.D(_03268_),
    .Q(\pcpi_mul.rs2[21] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _29781_ (.D(_03269_),
    .Q(\pcpi_mul.rs2[22] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _29782_ (.D(_03270_),
    .Q(\pcpi_mul.rs2[23] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _29783_ (.D(_03271_),
    .Q(\pcpi_mul.rs2[24] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _29784_ (.D(_03272_),
    .Q(\pcpi_mul.rs2[25] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _29785_ (.D(_03273_),
    .Q(\pcpi_mul.rs2[26] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _29786_ (.D(_03274_),
    .Q(\pcpi_mul.rs2[27] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _29787_ (.D(_03275_),
    .Q(\pcpi_mul.rs2[28] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _29788_ (.D(_03276_),
    .Q(\pcpi_mul.rs2[29] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29789_ (.D(_03277_),
    .Q(\pcpi_mul.rs2[30] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _29790_ (.D(_03278_),
    .Q(\pcpi_mul.rs2[31] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29791_ (.D(_03279_),
    .Q(\cpuregs[17][0] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29792_ (.D(_03280_),
    .Q(\cpuregs[17][1] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29793_ (.D(_03281_),
    .Q(\cpuregs[17][2] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29794_ (.D(_03282_),
    .Q(\cpuregs[17][3] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29795_ (.D(_03283_),
    .Q(\cpuregs[17][4] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29796_ (.D(_03284_),
    .Q(\cpuregs[17][5] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29797_ (.D(_03285_),
    .Q(\cpuregs[17][6] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29798_ (.D(_03286_),
    .Q(\cpuregs[17][7] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29799_ (.D(_03287_),
    .Q(\cpuregs[17][8] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29800_ (.D(_03288_),
    .Q(\cpuregs[17][9] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29801_ (.D(_03289_),
    .Q(\cpuregs[17][10] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29802_ (.D(_03290_),
    .Q(\cpuregs[17][11] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29803_ (.D(_03291_),
    .Q(\cpuregs[17][12] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29804_ (.D(_03292_),
    .Q(\cpuregs[17][13] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29805_ (.D(_03293_),
    .Q(\cpuregs[17][14] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29806_ (.D(_03294_),
    .Q(\cpuregs[17][15] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29807_ (.D(_03295_),
    .Q(\cpuregs[17][16] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29808_ (.D(_03296_),
    .Q(\cpuregs[17][17] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29809_ (.D(_03297_),
    .Q(\cpuregs[17][18] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29810_ (.D(_03298_),
    .Q(\cpuregs[17][19] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29811_ (.D(_03299_),
    .Q(\cpuregs[17][20] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29812_ (.D(_03300_),
    .Q(\cpuregs[17][21] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29813_ (.D(_03301_),
    .Q(\cpuregs[17][22] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29814_ (.D(_03302_),
    .Q(\cpuregs[17][23] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29815_ (.D(_03303_),
    .Q(\cpuregs[17][24] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29816_ (.D(_03304_),
    .Q(\cpuregs[17][25] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29817_ (.D(_03305_),
    .Q(\cpuregs[17][26] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29818_ (.D(_03306_),
    .Q(\cpuregs[17][27] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29819_ (.D(_03307_),
    .Q(\cpuregs[17][28] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29820_ (.D(_03308_),
    .Q(\cpuregs[17][29] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29821_ (.D(_03309_),
    .Q(\cpuregs[17][30] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29822_ (.D(_03310_),
    .Q(\cpuregs[17][31] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29823_ (.D(_03311_),
    .Q(\cpuregs[16][0] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29824_ (.D(_03312_),
    .Q(\cpuregs[16][1] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29825_ (.D(_03313_),
    .Q(\cpuregs[16][2] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29826_ (.D(_03314_),
    .Q(\cpuregs[16][3] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29827_ (.D(_03315_),
    .Q(\cpuregs[16][4] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29828_ (.D(_03316_),
    .Q(\cpuregs[16][5] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29829_ (.D(_03317_),
    .Q(\cpuregs[16][6] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29830_ (.D(_03318_),
    .Q(\cpuregs[16][7] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29831_ (.D(_03319_),
    .Q(\cpuregs[16][8] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29832_ (.D(_03320_),
    .Q(\cpuregs[16][9] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29833_ (.D(_03321_),
    .Q(\cpuregs[16][10] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29834_ (.D(_03322_),
    .Q(\cpuregs[16][11] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29835_ (.D(_03323_),
    .Q(\cpuregs[16][12] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29836_ (.D(_03324_),
    .Q(\cpuregs[16][13] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29837_ (.D(_03325_),
    .Q(\cpuregs[16][14] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29838_ (.D(_03326_),
    .Q(\cpuregs[16][15] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29839_ (.D(_03327_),
    .Q(\cpuregs[16][16] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29840_ (.D(_03328_),
    .Q(\cpuregs[16][17] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29841_ (.D(_03329_),
    .Q(\cpuregs[16][18] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29842_ (.D(_03330_),
    .Q(\cpuregs[16][19] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29843_ (.D(_03331_),
    .Q(\cpuregs[16][20] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29844_ (.D(_03332_),
    .Q(\cpuregs[16][21] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29845_ (.D(_03333_),
    .Q(\cpuregs[16][22] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29846_ (.D(_03334_),
    .Q(\cpuregs[16][23] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29847_ (.D(_03335_),
    .Q(\cpuregs[16][24] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29848_ (.D(_03336_),
    .Q(\cpuregs[16][25] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29849_ (.D(_03337_),
    .Q(\cpuregs[16][26] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29850_ (.D(_03338_),
    .Q(\cpuregs[16][27] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29851_ (.D(_03339_),
    .Q(\cpuregs[16][28] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29852_ (.D(_03340_),
    .Q(\cpuregs[16][29] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29853_ (.D(_03341_),
    .Q(\cpuregs[16][30] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29854_ (.D(_03342_),
    .Q(\cpuregs[16][31] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29855_ (.D(_03343_),
    .Q(\cpuregs[12][0] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29856_ (.D(_03344_),
    .Q(\cpuregs[12][1] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29857_ (.D(_03345_),
    .Q(\cpuregs[12][2] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29858_ (.D(_03346_),
    .Q(\cpuregs[12][3] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29859_ (.D(_03347_),
    .Q(\cpuregs[12][4] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29860_ (.D(_03348_),
    .Q(\cpuregs[12][5] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29861_ (.D(_03349_),
    .Q(\cpuregs[12][6] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29862_ (.D(_03350_),
    .Q(\cpuregs[12][7] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29863_ (.D(_03351_),
    .Q(\cpuregs[12][8] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29864_ (.D(_03352_),
    .Q(\cpuregs[12][9] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29865_ (.D(_03353_),
    .Q(\cpuregs[12][10] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29866_ (.D(_03354_),
    .Q(\cpuregs[12][11] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29867_ (.D(_03355_),
    .Q(\cpuregs[12][12] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29868_ (.D(_03356_),
    .Q(\cpuregs[12][13] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29869_ (.D(_03357_),
    .Q(\cpuregs[12][14] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29870_ (.D(_03358_),
    .Q(\cpuregs[12][15] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29871_ (.D(_03359_),
    .Q(\cpuregs[12][16] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29872_ (.D(_03360_),
    .Q(\cpuregs[12][17] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29873_ (.D(_03361_),
    .Q(\cpuregs[12][18] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29874_ (.D(_03362_),
    .Q(\cpuregs[12][19] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29875_ (.D(_03363_),
    .Q(\cpuregs[12][20] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29876_ (.D(_03364_),
    .Q(\cpuregs[12][21] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29877_ (.D(_03365_),
    .Q(\cpuregs[12][22] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29878_ (.D(_03366_),
    .Q(\cpuregs[12][23] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29879_ (.D(_03367_),
    .Q(\cpuregs[12][24] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29880_ (.D(_03368_),
    .Q(\cpuregs[12][25] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29881_ (.D(_03369_),
    .Q(\cpuregs[12][26] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29882_ (.D(_03370_),
    .Q(\cpuregs[12][27] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29883_ (.D(_03371_),
    .Q(\cpuregs[12][28] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29884_ (.D(_03372_),
    .Q(\cpuregs[12][29] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29885_ (.D(_03373_),
    .Q(\cpuregs[12][30] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29886_ (.D(_03374_),
    .Q(\cpuregs[12][31] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29887_ (.D(_03375_),
    .Q(\cpuregs[1][0] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29888_ (.D(_03376_),
    .Q(\cpuregs[1][1] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29889_ (.D(_03377_),
    .Q(\cpuregs[1][2] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29890_ (.D(_03378_),
    .Q(\cpuregs[1][3] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29891_ (.D(_03379_),
    .Q(\cpuregs[1][4] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29892_ (.D(_03380_),
    .Q(\cpuregs[1][5] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29893_ (.D(_03381_),
    .Q(\cpuregs[1][6] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29894_ (.D(_03382_),
    .Q(\cpuregs[1][7] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29895_ (.D(_03383_),
    .Q(\cpuregs[1][8] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29896_ (.D(_03384_),
    .Q(\cpuregs[1][9] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29897_ (.D(_03385_),
    .Q(\cpuregs[1][10] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29898_ (.D(_03386_),
    .Q(\cpuregs[1][11] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29899_ (.D(_03387_),
    .Q(\cpuregs[1][12] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29900_ (.D(_03388_),
    .Q(\cpuregs[1][13] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29901_ (.D(_03389_),
    .Q(\cpuregs[1][14] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29902_ (.D(_03390_),
    .Q(\cpuregs[1][15] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29903_ (.D(_03391_),
    .Q(\cpuregs[1][16] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29904_ (.D(_03392_),
    .Q(\cpuregs[1][17] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29905_ (.D(_03393_),
    .Q(\cpuregs[1][18] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29906_ (.D(_03394_),
    .Q(\cpuregs[1][19] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29907_ (.D(_03395_),
    .Q(\cpuregs[1][20] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29908_ (.D(_03396_),
    .Q(\cpuregs[1][21] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29909_ (.D(_03397_),
    .Q(\cpuregs[1][22] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29910_ (.D(_03398_),
    .Q(\cpuregs[1][23] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29911_ (.D(_03399_),
    .Q(\cpuregs[1][24] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29912_ (.D(_03400_),
    .Q(\cpuregs[1][25] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29913_ (.D(_03401_),
    .Q(\cpuregs[1][26] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29914_ (.D(_03402_),
    .Q(\cpuregs[1][27] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29915_ (.D(_03403_),
    .Q(\cpuregs[1][28] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29916_ (.D(_03404_),
    .Q(\cpuregs[1][29] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29917_ (.D(_03405_),
    .Q(\cpuregs[1][30] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29918_ (.D(_03406_),
    .Q(\cpuregs[1][31] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29919_ (.D(_03407_),
    .Q(\cpuregs[3][0] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29920_ (.D(_03408_),
    .Q(\cpuregs[3][1] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29921_ (.D(_03409_),
    .Q(\cpuregs[3][2] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29922_ (.D(_03410_),
    .Q(\cpuregs[3][3] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29923_ (.D(_03411_),
    .Q(\cpuregs[3][4] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29924_ (.D(_03412_),
    .Q(\cpuregs[3][5] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29925_ (.D(_03413_),
    .Q(\cpuregs[3][6] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29926_ (.D(_03414_),
    .Q(\cpuregs[3][7] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29927_ (.D(_03415_),
    .Q(\cpuregs[3][8] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29928_ (.D(_03416_),
    .Q(\cpuregs[3][9] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29929_ (.D(_03417_),
    .Q(\cpuregs[3][10] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29930_ (.D(_03418_),
    .Q(\cpuregs[3][11] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29931_ (.D(_03419_),
    .Q(\cpuregs[3][12] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29932_ (.D(_03420_),
    .Q(\cpuregs[3][13] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29933_ (.D(_03421_),
    .Q(\cpuregs[3][14] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29934_ (.D(_03422_),
    .Q(\cpuregs[3][15] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29935_ (.D(_03423_),
    .Q(\cpuregs[3][16] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29936_ (.D(_03424_),
    .Q(\cpuregs[3][17] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29937_ (.D(_03425_),
    .Q(\cpuregs[3][18] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29938_ (.D(_03426_),
    .Q(\cpuregs[3][19] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29939_ (.D(_03427_),
    .Q(\cpuregs[3][20] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29940_ (.D(_03428_),
    .Q(\cpuregs[3][21] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29941_ (.D(_03429_),
    .Q(\cpuregs[3][22] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29942_ (.D(_03430_),
    .Q(\cpuregs[3][23] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29943_ (.D(_03431_),
    .Q(\cpuregs[3][24] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29944_ (.D(_03432_),
    .Q(\cpuregs[3][25] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29945_ (.D(_03433_),
    .Q(\cpuregs[3][26] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29946_ (.D(_03434_),
    .Q(\cpuregs[3][27] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29947_ (.D(_03435_),
    .Q(\cpuregs[3][28] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29948_ (.D(_03436_),
    .Q(\cpuregs[3][29] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29949_ (.D(_03437_),
    .Q(\cpuregs[3][30] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29950_ (.D(_03438_),
    .Q(\cpuregs[3][31] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29951_ (.D(_03439_),
    .Q(\cpuregs[11][0] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29952_ (.D(_03440_),
    .Q(\cpuregs[11][1] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29953_ (.D(_03441_),
    .Q(\cpuregs[11][2] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29954_ (.D(_03442_),
    .Q(\cpuregs[11][3] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29955_ (.D(_03443_),
    .Q(\cpuregs[11][4] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29956_ (.D(_03444_),
    .Q(\cpuregs[11][5] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29957_ (.D(_03445_),
    .Q(\cpuregs[11][6] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29958_ (.D(_03446_),
    .Q(\cpuregs[11][7] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29959_ (.D(_03447_),
    .Q(\cpuregs[11][8] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29960_ (.D(_03448_),
    .Q(\cpuregs[11][9] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29961_ (.D(_03449_),
    .Q(\cpuregs[11][10] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29962_ (.D(_03450_),
    .Q(\cpuregs[11][11] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29963_ (.D(_03451_),
    .Q(\cpuregs[11][12] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29964_ (.D(_03452_),
    .Q(\cpuregs[11][13] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29965_ (.D(_03453_),
    .Q(\cpuregs[11][14] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29966_ (.D(_03454_),
    .Q(\cpuregs[11][15] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29967_ (.D(_03455_),
    .Q(\cpuregs[11][16] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29968_ (.D(_03456_),
    .Q(\cpuregs[11][17] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29969_ (.D(_03457_),
    .Q(\cpuregs[11][18] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29970_ (.D(_03458_),
    .Q(\cpuregs[11][19] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29971_ (.D(_03459_),
    .Q(\cpuregs[11][20] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29972_ (.D(_03460_),
    .Q(\cpuregs[11][21] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29973_ (.D(_03461_),
    .Q(\cpuregs[11][22] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29974_ (.D(_03462_),
    .Q(\cpuregs[11][23] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29975_ (.D(_03463_),
    .Q(\cpuregs[11][24] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29976_ (.D(_03464_),
    .Q(\cpuregs[11][25] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29977_ (.D(_03465_),
    .Q(\cpuregs[11][26] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29978_ (.D(_03466_),
    .Q(\cpuregs[11][27] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29979_ (.D(_03467_),
    .Q(\cpuregs[11][28] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29980_ (.D(_03468_),
    .Q(\cpuregs[11][29] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29981_ (.D(_03469_),
    .Q(\cpuregs[11][30] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29982_ (.D(_03470_),
    .Q(\cpuregs[11][31] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29983_ (.D(_03471_),
    .Q(\cpuregs[15][0] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29984_ (.D(_03472_),
    .Q(\cpuregs[15][1] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29985_ (.D(_03473_),
    .Q(\cpuregs[15][2] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29986_ (.D(_03474_),
    .Q(\cpuregs[15][3] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29987_ (.D(_03475_),
    .Q(\cpuregs[15][4] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29988_ (.D(_03476_),
    .Q(\cpuregs[15][5] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29989_ (.D(_03477_),
    .Q(\cpuregs[15][6] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29990_ (.D(_03478_),
    .Q(\cpuregs[15][7] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29991_ (.D(_03479_),
    .Q(\cpuregs[15][8] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29992_ (.D(_03480_),
    .Q(\cpuregs[15][9] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29993_ (.D(_03481_),
    .Q(\cpuregs[15][10] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29994_ (.D(_03482_),
    .Q(\cpuregs[15][11] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29995_ (.D(_03483_),
    .Q(\cpuregs[15][12] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29996_ (.D(_03484_),
    .Q(\cpuregs[15][13] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29997_ (.D(_03485_),
    .Q(\cpuregs[15][14] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29998_ (.D(_03486_),
    .Q(\cpuregs[15][15] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _29999_ (.D(_03487_),
    .Q(\cpuregs[15][16] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30000_ (.D(_03488_),
    .Q(\cpuregs[15][17] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30001_ (.D(_03489_),
    .Q(\cpuregs[15][18] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30002_ (.D(_03490_),
    .Q(\cpuregs[15][19] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30003_ (.D(_03491_),
    .Q(\cpuregs[15][20] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30004_ (.D(_03492_),
    .Q(\cpuregs[15][21] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30005_ (.D(_03493_),
    .Q(\cpuregs[15][22] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30006_ (.D(_03494_),
    .Q(\cpuregs[15][23] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30007_ (.D(_03495_),
    .Q(\cpuregs[15][24] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30008_ (.D(_03496_),
    .Q(\cpuregs[15][25] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30009_ (.D(_03497_),
    .Q(\cpuregs[15][26] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30010_ (.D(_03498_),
    .Q(\cpuregs[15][27] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30011_ (.D(_03499_),
    .Q(\cpuregs[15][28] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30012_ (.D(_03500_),
    .Q(\cpuregs[15][29] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30013_ (.D(_03501_),
    .Q(\cpuregs[15][30] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30014_ (.D(_03502_),
    .Q(\cpuregs[15][31] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30015_ (.D(_03503_),
    .Q(\latched_rd[4] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30016_ (.D(_03504_),
    .Q(\cpuregs[7][0] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30017_ (.D(_03505_),
    .Q(\cpuregs[7][1] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30018_ (.D(_03506_),
    .Q(\cpuregs[7][2] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30019_ (.D(_03507_),
    .Q(\cpuregs[7][3] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30020_ (.D(_03508_),
    .Q(\cpuregs[7][4] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30021_ (.D(_03509_),
    .Q(\cpuregs[7][5] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30022_ (.D(_03510_),
    .Q(\cpuregs[7][6] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30023_ (.D(_03511_),
    .Q(\cpuregs[7][7] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30024_ (.D(_03512_),
    .Q(\cpuregs[7][8] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30025_ (.D(_03513_),
    .Q(\cpuregs[7][9] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30026_ (.D(_03514_),
    .Q(\cpuregs[7][10] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30027_ (.D(_03515_),
    .Q(\cpuregs[7][11] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30028_ (.D(_03516_),
    .Q(\cpuregs[7][12] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30029_ (.D(_03517_),
    .Q(\cpuregs[7][13] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30030_ (.D(_03518_),
    .Q(\cpuregs[7][14] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30031_ (.D(_03519_),
    .Q(\cpuregs[7][15] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30032_ (.D(_03520_),
    .Q(\cpuregs[7][16] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30033_ (.D(_03521_),
    .Q(\cpuregs[7][17] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30034_ (.D(_03522_),
    .Q(\cpuregs[7][18] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30035_ (.D(_03523_),
    .Q(\cpuregs[7][19] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30036_ (.D(_03524_),
    .Q(\cpuregs[7][20] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30037_ (.D(_03525_),
    .Q(\cpuregs[7][21] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30038_ (.D(_03526_),
    .Q(\cpuregs[7][22] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30039_ (.D(_03527_),
    .Q(\cpuregs[7][23] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30040_ (.D(_03528_),
    .Q(\cpuregs[7][24] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30041_ (.D(_03529_),
    .Q(\cpuregs[7][25] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30042_ (.D(_03530_),
    .Q(\cpuregs[7][26] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30043_ (.D(_03531_),
    .Q(\cpuregs[7][27] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30044_ (.D(_03532_),
    .Q(\cpuregs[7][28] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30045_ (.D(_03533_),
    .Q(\cpuregs[7][29] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30046_ (.D(_03534_),
    .Q(\cpuregs[7][30] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30047_ (.D(_03535_),
    .Q(\cpuregs[7][31] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _30048_ (.D(_03536_),
    .Q(net238),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _30049_ (.D(_03537_),
    .Q(net249),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _30050_ (.D(_03538_),
    .Q(net260),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _30051_ (.D(_03539_),
    .Q(net263),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _30052_ (.D(_03540_),
    .Q(net264),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _30053_ (.D(_03541_),
    .Q(net265),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _30054_ (.D(_03542_),
    .Q(net266),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _30055_ (.D(_03543_),
    .Q(net267),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _30056_ (.D(_03544_),
    .Q(net268),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _30057_ (.D(_03545_),
    .Q(net269),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _30058_ (.D(_03546_),
    .Q(net239),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _30059_ (.D(_03547_),
    .Q(net240),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _30060_ (.D(_03548_),
    .Q(net241),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _30061_ (.D(_03549_),
    .Q(net242),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _30062_ (.D(_03550_),
    .Q(net243),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _30063_ (.D(_03551_),
    .Q(net244),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _30064_ (.D(_03552_),
    .Q(net245),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _30065_ (.D(_03553_),
    .Q(net246),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _30066_ (.D(_03554_),
    .Q(net247),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _30067_ (.D(_03555_),
    .Q(net248),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _30068_ (.D(_03556_),
    .Q(net250),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _30069_ (.D(_03557_),
    .Q(net251),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _30070_ (.D(_03558_),
    .Q(net252),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _30071_ (.D(_03559_),
    .Q(net253),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _30072_ (.D(_03560_),
    .Q(net254),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _30073_ (.D(_03561_),
    .Q(net255),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _30074_ (.D(_03562_),
    .Q(net256),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _30075_ (.D(_03563_),
    .Q(net257),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _30076_ (.D(_03564_),
    .Q(net258),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _30077_ (.D(_03565_),
    .Q(net259),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _30078_ (.D(_03566_),
    .Q(net261),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _30079_ (.D(_03567_),
    .Q(net262),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30080_ (.D(_03568_),
    .Q(\cpuregs[19][0] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30081_ (.D(_03569_),
    .Q(\cpuregs[19][1] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30082_ (.D(_03570_),
    .Q(\cpuregs[19][2] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30083_ (.D(_03571_),
    .Q(\cpuregs[19][3] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30084_ (.D(_03572_),
    .Q(\cpuregs[19][4] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30085_ (.D(_03573_),
    .Q(\cpuregs[19][5] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30086_ (.D(_03574_),
    .Q(\cpuregs[19][6] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30087_ (.D(_03575_),
    .Q(\cpuregs[19][7] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30088_ (.D(_03576_),
    .Q(\cpuregs[19][8] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30089_ (.D(_03577_),
    .Q(\cpuregs[19][9] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30090_ (.D(_03578_),
    .Q(\cpuregs[19][10] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30091_ (.D(_03579_),
    .Q(\cpuregs[19][11] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30092_ (.D(_03580_),
    .Q(\cpuregs[19][12] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30093_ (.D(_03581_),
    .Q(\cpuregs[19][13] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30094_ (.D(_03582_),
    .Q(\cpuregs[19][14] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30095_ (.D(_03583_),
    .Q(\cpuregs[19][15] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30096_ (.D(_03584_),
    .Q(\cpuregs[19][16] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30097_ (.D(_03585_),
    .Q(\cpuregs[19][17] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30098_ (.D(_03586_),
    .Q(\cpuregs[19][18] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30099_ (.D(_03587_),
    .Q(\cpuregs[19][19] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30100_ (.D(_03588_),
    .Q(\cpuregs[19][20] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30101_ (.D(_03589_),
    .Q(\cpuregs[19][21] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30102_ (.D(_03590_),
    .Q(\cpuregs[19][22] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30103_ (.D(_03591_),
    .Q(\cpuregs[19][23] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30104_ (.D(_03592_),
    .Q(\cpuregs[19][24] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30105_ (.D(_03593_),
    .Q(\cpuregs[19][25] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30106_ (.D(_03594_),
    .Q(\cpuregs[19][26] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30107_ (.D(_03595_),
    .Q(\cpuregs[19][27] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30108_ (.D(_03596_),
    .Q(\cpuregs[19][28] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30109_ (.D(_03597_),
    .Q(\cpuregs[19][29] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30110_ (.D(_03598_),
    .Q(\cpuregs[19][30] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30111_ (.D(_03599_),
    .Q(\cpuregs[19][31] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30112_ (.D(_03600_),
    .Q(\cpuregs[4][0] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30113_ (.D(_03601_),
    .Q(\cpuregs[4][1] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30114_ (.D(_03602_),
    .Q(\cpuregs[4][2] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30115_ (.D(_03603_),
    .Q(\cpuregs[4][3] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30116_ (.D(_03604_),
    .Q(\cpuregs[4][4] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30117_ (.D(_03605_),
    .Q(\cpuregs[4][5] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30118_ (.D(_03606_),
    .Q(\cpuregs[4][6] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30119_ (.D(_03607_),
    .Q(\cpuregs[4][7] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30120_ (.D(_03608_),
    .Q(\cpuregs[4][8] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30121_ (.D(_03609_),
    .Q(\cpuregs[4][9] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30122_ (.D(_03610_),
    .Q(\cpuregs[4][10] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30123_ (.D(_03611_),
    .Q(\cpuregs[4][11] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30124_ (.D(_03612_),
    .Q(\cpuregs[4][12] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30125_ (.D(_03613_),
    .Q(\cpuregs[4][13] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30126_ (.D(_03614_),
    .Q(\cpuregs[4][14] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30127_ (.D(_03615_),
    .Q(\cpuregs[4][15] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30128_ (.D(_03616_),
    .Q(\cpuregs[4][16] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30129_ (.D(_03617_),
    .Q(\cpuregs[4][17] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30130_ (.D(_03618_),
    .Q(\cpuregs[4][18] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30131_ (.D(_03619_),
    .Q(\cpuregs[4][19] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30132_ (.D(_03620_),
    .Q(\cpuregs[4][20] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30133_ (.D(_03621_),
    .Q(\cpuregs[4][21] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30134_ (.D(_03622_),
    .Q(\cpuregs[4][22] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30135_ (.D(_03623_),
    .Q(\cpuregs[4][23] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30136_ (.D(_03624_),
    .Q(\cpuregs[4][24] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30137_ (.D(_03625_),
    .Q(\cpuregs[4][25] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30138_ (.D(_03626_),
    .Q(\cpuregs[4][26] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30139_ (.D(_03627_),
    .Q(\cpuregs[4][27] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30140_ (.D(_03628_),
    .Q(\cpuregs[4][28] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30141_ (.D(_03629_),
    .Q(\cpuregs[4][29] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30142_ (.D(_03630_),
    .Q(\cpuregs[4][30] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30143_ (.D(_03631_),
    .Q(\cpuregs[4][31] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _30144_ (.D(_03632_),
    .Q(net200),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _30145_ (.D(_03633_),
    .Q(net211),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _30146_ (.D(_03634_),
    .Q(net222),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _30147_ (.D(_03635_),
    .Q(net225),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _30148_ (.D(_03636_),
    .Q(net226),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _30149_ (.D(_03637_),
    .Q(net227),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _30150_ (.D(_03638_),
    .Q(net228),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _30151_ (.D(_03639_),
    .Q(net229),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _30152_ (.D(_03640_),
    .Q(net368),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _30153_ (.D(_03641_),
    .Q(net369),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _30154_ (.D(_03642_),
    .Q(net339),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _30155_ (.D(_03643_),
    .Q(net340),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _30156_ (.D(_03644_),
    .Q(net341),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _30157_ (.D(_03645_),
    .Q(net342),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _30158_ (.D(_03646_),
    .Q(net343),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _30159_ (.D(_03647_),
    .Q(net344),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _30160_ (.D(_03648_),
    .Q(net345),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _30161_ (.D(_03649_),
    .Q(net346),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _30162_ (.D(_03650_),
    .Q(net347),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _30163_ (.D(_03651_),
    .Q(net348),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _30164_ (.D(_03652_),
    .Q(net350),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _30165_ (.D(_03653_),
    .Q(net351),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _30166_ (.D(_03654_),
    .Q(net352),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _30167_ (.D(_03655_),
    .Q(net353),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _30168_ (.D(_03656_),
    .Q(net354),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _30169_ (.D(_03657_),
    .Q(net355),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _30170_ (.D(_03658_),
    .Q(net356),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _30171_ (.D(_03659_),
    .Q(net357),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _30172_ (.D(_03660_),
    .Q(net358),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _30173_ (.D(_03661_),
    .Q(net359),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _30174_ (.D(_03662_),
    .Q(net361),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _30175_ (.D(_03663_),
    .Q(net362),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30176_ (.D(_03664_),
    .Q(\cpuregs[9][0] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30177_ (.D(_03665_),
    .Q(\cpuregs[9][1] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30178_ (.D(_03666_),
    .Q(\cpuregs[9][2] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30179_ (.D(_03667_),
    .Q(\cpuregs[9][3] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30180_ (.D(_03668_),
    .Q(\cpuregs[9][4] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30181_ (.D(_03669_),
    .Q(\cpuregs[9][5] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30182_ (.D(_03670_),
    .Q(\cpuregs[9][6] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30183_ (.D(_03671_),
    .Q(\cpuregs[9][7] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30184_ (.D(_03672_),
    .Q(\cpuregs[9][8] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30185_ (.D(_03673_),
    .Q(\cpuregs[9][9] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30186_ (.D(_03674_),
    .Q(\cpuregs[9][10] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30187_ (.D(_03675_),
    .Q(\cpuregs[9][11] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30188_ (.D(_03676_),
    .Q(\cpuregs[9][12] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30189_ (.D(_03677_),
    .Q(\cpuregs[9][13] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30190_ (.D(_03678_),
    .Q(\cpuregs[9][14] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30191_ (.D(_03679_),
    .Q(\cpuregs[9][15] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30192_ (.D(_03680_),
    .Q(\cpuregs[9][16] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30193_ (.D(_03681_),
    .Q(\cpuregs[9][17] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30194_ (.D(_03682_),
    .Q(\cpuregs[9][18] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30195_ (.D(_03683_),
    .Q(\cpuregs[9][19] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30196_ (.D(_03684_),
    .Q(\cpuregs[9][20] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30197_ (.D(_03685_),
    .Q(\cpuregs[9][21] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30198_ (.D(_03686_),
    .Q(\cpuregs[9][22] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30199_ (.D(_03687_),
    .Q(\cpuregs[9][23] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30200_ (.D(_03688_),
    .Q(\cpuregs[9][24] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30201_ (.D(_03689_),
    .Q(\cpuregs[9][25] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30202_ (.D(_03690_),
    .Q(\cpuregs[9][26] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30203_ (.D(_03691_),
    .Q(\cpuregs[9][27] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30204_ (.D(_03692_),
    .Q(\cpuregs[9][28] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30205_ (.D(_03693_),
    .Q(\cpuregs[9][29] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30206_ (.D(_03694_),
    .Q(\cpuregs[9][30] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30207_ (.D(_03695_),
    .Q(\cpuregs[9][31] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30208_ (.D(_03696_),
    .Q(\cpuregs[6][0] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30209_ (.D(_03697_),
    .Q(\cpuregs[6][1] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30210_ (.D(_03698_),
    .Q(\cpuregs[6][2] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30211_ (.D(_03699_),
    .Q(\cpuregs[6][3] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30212_ (.D(_03700_),
    .Q(\cpuregs[6][4] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30213_ (.D(_03701_),
    .Q(\cpuregs[6][5] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30214_ (.D(_03702_),
    .Q(\cpuregs[6][6] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30215_ (.D(_03703_),
    .Q(\cpuregs[6][7] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30216_ (.D(_03704_),
    .Q(\cpuregs[6][8] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30217_ (.D(_03705_),
    .Q(\cpuregs[6][9] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30218_ (.D(_03706_),
    .Q(\cpuregs[6][10] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30219_ (.D(_03707_),
    .Q(\cpuregs[6][11] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30220_ (.D(_03708_),
    .Q(\cpuregs[6][12] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30221_ (.D(_03709_),
    .Q(\cpuregs[6][13] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30222_ (.D(_03710_),
    .Q(\cpuregs[6][14] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30223_ (.D(_03711_),
    .Q(\cpuregs[6][15] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30224_ (.D(_03712_),
    .Q(\cpuregs[6][16] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30225_ (.D(_03713_),
    .Q(\cpuregs[6][17] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30226_ (.D(_03714_),
    .Q(\cpuregs[6][18] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30227_ (.D(_03715_),
    .Q(\cpuregs[6][19] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30228_ (.D(_03716_),
    .Q(\cpuregs[6][20] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30229_ (.D(_03717_),
    .Q(\cpuregs[6][21] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30230_ (.D(_03718_),
    .Q(\cpuregs[6][22] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30231_ (.D(_03719_),
    .Q(\cpuregs[6][23] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30232_ (.D(_03720_),
    .Q(\cpuregs[6][24] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30233_ (.D(_03721_),
    .Q(\cpuregs[6][25] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30234_ (.D(_03722_),
    .Q(\cpuregs[6][26] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30235_ (.D(_03723_),
    .Q(\cpuregs[6][27] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30236_ (.D(_03724_),
    .Q(\cpuregs[6][28] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30237_ (.D(_03725_),
    .Q(\cpuregs[6][29] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30238_ (.D(_03726_),
    .Q(\cpuregs[6][30] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30239_ (.D(_03727_),
    .Q(\cpuregs[6][31] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30240_ (.D(_03728_),
    .Q(\pcpi_mul.active[0] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _30241_ (.D(_03729_),
    .Q(\pcpi_mul.active[1] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _30242_ (.D(_03730_),
    .Q(net408),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30243_ (.D(_03731_),
    .Q(\count_cycle[0] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30244_ (.D(_03732_),
    .Q(\count_cycle[1] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30245_ (.D(_03733_),
    .Q(\count_cycle[2] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30246_ (.D(_03734_),
    .Q(\count_cycle[3] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30247_ (.D(_03735_),
    .Q(\count_cycle[4] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30248_ (.D(_03736_),
    .Q(\count_cycle[5] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30249_ (.D(_03737_),
    .Q(\count_cycle[6] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30250_ (.D(_03738_),
    .Q(\count_cycle[7] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30251_ (.D(_03739_),
    .Q(\count_cycle[8] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30252_ (.D(_03740_),
    .Q(\count_cycle[9] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30253_ (.D(_03741_),
    .Q(\count_cycle[10] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30254_ (.D(_03742_),
    .Q(\count_cycle[11] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30255_ (.D(_03743_),
    .Q(\count_cycle[12] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30256_ (.D(_03744_),
    .Q(\count_cycle[13] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30257_ (.D(_03745_),
    .Q(\count_cycle[14] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30258_ (.D(_03746_),
    .Q(\count_cycle[15] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30259_ (.D(_03747_),
    .Q(\count_cycle[16] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30260_ (.D(_03748_),
    .Q(\count_cycle[17] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30261_ (.D(_03749_),
    .Q(\count_cycle[18] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30262_ (.D(_03750_),
    .Q(\count_cycle[19] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30263_ (.D(_03751_),
    .Q(\count_cycle[20] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30264_ (.D(_03752_),
    .Q(\count_cycle[21] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30265_ (.D(_03753_),
    .Q(\count_cycle[22] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30266_ (.D(_03754_),
    .Q(\count_cycle[23] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30267_ (.D(_03755_),
    .Q(\count_cycle[24] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30268_ (.D(_03756_),
    .Q(\count_cycle[25] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30269_ (.D(_03757_),
    .Q(\count_cycle[26] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30270_ (.D(_03758_),
    .Q(\count_cycle[27] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30271_ (.D(_03759_),
    .Q(\count_cycle[28] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30272_ (.D(_03760_),
    .Q(\count_cycle[29] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30273_ (.D(_03761_),
    .Q(\count_cycle[30] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30274_ (.D(_03762_),
    .Q(\count_cycle[31] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30275_ (.D(_03763_),
    .Q(\count_cycle[32] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30276_ (.D(_03764_),
    .Q(\count_cycle[33] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30277_ (.D(_03765_),
    .Q(\count_cycle[34] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30278_ (.D(_03766_),
    .Q(\count_cycle[35] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30279_ (.D(_03767_),
    .Q(\count_cycle[36] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30280_ (.D(_03768_),
    .Q(\count_cycle[37] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30281_ (.D(_03769_),
    .Q(\count_cycle[38] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30282_ (.D(_03770_),
    .Q(\count_cycle[39] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30283_ (.D(_03771_),
    .Q(\count_cycle[40] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30284_ (.D(_03772_),
    .Q(\count_cycle[41] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30285_ (.D(_03773_),
    .Q(\count_cycle[42] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30286_ (.D(_03774_),
    .Q(\count_cycle[43] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30287_ (.D(_03775_),
    .Q(\count_cycle[44] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30288_ (.D(_03776_),
    .Q(\count_cycle[45] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30289_ (.D(_03777_),
    .Q(\count_cycle[46] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30290_ (.D(_03778_),
    .Q(\count_cycle[47] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30291_ (.D(_03779_),
    .Q(\count_cycle[48] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30292_ (.D(_03780_),
    .Q(\count_cycle[49] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30293_ (.D(_03781_),
    .Q(\count_cycle[50] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30294_ (.D(_03782_),
    .Q(\count_cycle[51] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30295_ (.D(_03783_),
    .Q(\count_cycle[52] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30296_ (.D(_03784_),
    .Q(\count_cycle[53] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30297_ (.D(_03785_),
    .Q(\count_cycle[54] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30298_ (.D(_03786_),
    .Q(\count_cycle[55] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30299_ (.D(_03787_),
    .Q(\count_cycle[56] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30300_ (.D(_03788_),
    .Q(\count_cycle[57] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30301_ (.D(_03789_),
    .Q(\count_cycle[58] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30302_ (.D(_03790_),
    .Q(\count_cycle[59] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30303_ (.D(_03791_),
    .Q(\count_cycle[60] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30304_ (.D(_03792_),
    .Q(\count_cycle[61] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30305_ (.D(_03793_),
    .Q(\count_cycle[62] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30306_ (.D(_03794_),
    .Q(\count_cycle[63] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30307_ (.D(_03795_),
    .Q(\timer[0] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30308_ (.D(_03796_),
    .Q(\timer[1] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30309_ (.D(_03797_),
    .Q(\timer[2] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30310_ (.D(_03798_),
    .Q(\timer[3] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30311_ (.D(_03799_),
    .Q(\timer[4] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30312_ (.D(_03800_),
    .Q(\timer[5] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30313_ (.D(_03801_),
    .Q(\timer[6] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30314_ (.D(_03802_),
    .Q(\timer[7] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30315_ (.D(_03803_),
    .Q(\timer[8] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30316_ (.D(_03804_),
    .Q(\timer[9] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30317_ (.D(_03805_),
    .Q(\timer[10] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30318_ (.D(_03806_),
    .Q(\timer[11] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30319_ (.D(_03807_),
    .Q(\timer[12] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30320_ (.D(_03808_),
    .Q(\timer[13] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30321_ (.D(_03809_),
    .Q(\timer[14] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30322_ (.D(_03810_),
    .Q(\timer[15] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30323_ (.D(_03811_),
    .Q(\timer[16] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _30324_ (.D(_03812_),
    .Q(\timer[17] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30325_ (.D(_03813_),
    .Q(\timer[18] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30326_ (.D(_03814_),
    .Q(\timer[19] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30327_ (.D(_03815_),
    .Q(\timer[20] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30328_ (.D(_03816_),
    .Q(\timer[21] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30329_ (.D(_03817_),
    .Q(\timer[22] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30330_ (.D(_03818_),
    .Q(\timer[23] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30331_ (.D(_03819_),
    .Q(\timer[24] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _30332_ (.D(_03820_),
    .Q(\timer[25] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30333_ (.D(_03821_),
    .Q(\timer[26] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30334_ (.D(_03822_),
    .Q(\timer[27] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30335_ (.D(_03823_),
    .Q(\timer[28] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30336_ (.D(_03824_),
    .Q(\timer[29] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30337_ (.D(_03825_),
    .Q(\timer[30] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _30338_ (.D(_03826_),
    .Q(\timer[31] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30339_ (.D(_03827_),
    .Q(pcpi_timeout),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30340_ (.D(_03828_),
    .Q(decoder_pseudo_trigger),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30341_ (.D(_03829_),
    .Q(is_compare),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30342_ (.D(_03830_),
    .Q(do_waitirq),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _30343_ (.D(_03831_),
    .Q(net237),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _30344_ (.D(_03832_),
    .Q(net370),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _30345_ (.D(_03833_),
    .Q(net102),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _30346_ (.D(_03834_),
    .Q(net113),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _30347_ (.D(_03835_),
    .Q(net124),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _30348_ (.D(_03836_),
    .Q(net127),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _30349_ (.D(_03837_),
    .Q(net128),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _30350_ (.D(_03838_),
    .Q(net129),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _30351_ (.D(_03839_),
    .Q(net130),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _30352_ (.D(_03840_),
    .Q(net131),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _30353_ (.D(_03841_),
    .Q(net132),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _30354_ (.D(_03842_),
    .Q(net133),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _30355_ (.D(_03843_),
    .Q(net103),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _30356_ (.D(_03844_),
    .Q(net104),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _30357_ (.D(_03845_),
    .Q(net105),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _30358_ (.D(_03846_),
    .Q(net106),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _30359_ (.D(_03847_),
    .Q(net107),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _30360_ (.D(_03848_),
    .Q(net108),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _30361_ (.D(_03849_),
    .Q(net109),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _30362_ (.D(_03850_),
    .Q(net110),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30363_ (.D(_03851_),
    .Q(net111),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _30364_ (.D(_03852_),
    .Q(net112),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _30365_ (.D(_03853_),
    .Q(net114),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _30366_ (.D(_03854_),
    .Q(net115),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _30367_ (.D(_03855_),
    .Q(net116),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _30368_ (.D(_03856_),
    .Q(net117),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _30369_ (.D(_03857_),
    .Q(net118),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _30370_ (.D(_03858_),
    .Q(net119),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _30371_ (.D(_03859_),
    .Q(net120),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _30372_ (.D(_03860_),
    .Q(net121),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _30373_ (.D(_03861_),
    .Q(net122),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _30374_ (.D(_03862_),
    .Q(net123),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _30375_ (.D(_03863_),
    .Q(net125),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _30376_ (.D(_03864_),
    .Q(net126),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30377_ (.D(_03865_),
    .Q(\count_instr[0] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30378_ (.D(_03866_),
    .Q(\count_instr[1] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30379_ (.D(_03867_),
    .Q(\count_instr[2] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30380_ (.D(_03868_),
    .Q(\count_instr[3] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30381_ (.D(_03869_),
    .Q(\count_instr[4] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30382_ (.D(_03870_),
    .Q(\count_instr[5] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30383_ (.D(_03871_),
    .Q(\count_instr[6] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30384_ (.D(_03872_),
    .Q(\count_instr[7] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30385_ (.D(_03873_),
    .Q(\count_instr[8] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30386_ (.D(_03874_),
    .Q(\count_instr[9] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30387_ (.D(_03875_),
    .Q(\count_instr[10] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30388_ (.D(_03876_),
    .Q(\count_instr[11] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30389_ (.D(_03877_),
    .Q(\count_instr[12] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30390_ (.D(_03878_),
    .Q(\count_instr[13] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30391_ (.D(_03879_),
    .Q(\count_instr[14] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30392_ (.D(_03880_),
    .Q(\count_instr[15] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30393_ (.D(_03881_),
    .Q(\count_instr[16] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30394_ (.D(_03882_),
    .Q(\count_instr[17] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30395_ (.D(_03883_),
    .Q(\count_instr[18] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30396_ (.D(_03884_),
    .Q(\count_instr[19] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30397_ (.D(_03885_),
    .Q(\count_instr[20] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30398_ (.D(_03886_),
    .Q(\count_instr[21] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30399_ (.D(_03887_),
    .Q(\count_instr[22] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30400_ (.D(_03888_),
    .Q(\count_instr[23] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30401_ (.D(_03889_),
    .Q(\count_instr[24] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30402_ (.D(_03890_),
    .Q(\count_instr[25] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30403_ (.D(_03891_),
    .Q(\count_instr[26] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30404_ (.D(_03892_),
    .Q(\count_instr[27] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30405_ (.D(_03893_),
    .Q(\count_instr[28] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30406_ (.D(_03894_),
    .Q(\count_instr[29] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30407_ (.D(_03895_),
    .Q(\count_instr[30] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30408_ (.D(_03896_),
    .Q(\count_instr[31] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30409_ (.D(_03897_),
    .Q(\count_instr[32] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30410_ (.D(_03898_),
    .Q(\count_instr[33] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30411_ (.D(_03899_),
    .Q(\count_instr[34] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30412_ (.D(_03900_),
    .Q(\count_instr[35] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30413_ (.D(_03901_),
    .Q(\count_instr[36] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30414_ (.D(_03902_),
    .Q(\count_instr[37] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30415_ (.D(_03903_),
    .Q(\count_instr[38] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30416_ (.D(_03904_),
    .Q(\count_instr[39] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30417_ (.D(_03905_),
    .Q(\count_instr[40] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30418_ (.D(_03906_),
    .Q(\count_instr[41] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30419_ (.D(_03907_),
    .Q(\count_instr[42] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30420_ (.D(_03908_),
    .Q(\count_instr[43] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30421_ (.D(_03909_),
    .Q(\count_instr[44] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30422_ (.D(_03910_),
    .Q(\count_instr[45] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30423_ (.D(_03911_),
    .Q(\count_instr[46] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30424_ (.D(_03912_),
    .Q(\count_instr[47] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30425_ (.D(_03913_),
    .Q(\count_instr[48] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30426_ (.D(_03914_),
    .Q(\count_instr[49] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30427_ (.D(_03915_),
    .Q(\count_instr[50] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30428_ (.D(_03916_),
    .Q(\count_instr[51] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30429_ (.D(_03917_),
    .Q(\count_instr[52] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30430_ (.D(_03918_),
    .Q(\count_instr[53] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30431_ (.D(_03919_),
    .Q(\count_instr[54] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30432_ (.D(_03920_),
    .Q(\count_instr[55] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30433_ (.D(_03921_),
    .Q(\count_instr[56] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30434_ (.D(_03922_),
    .Q(\count_instr[57] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30435_ (.D(_03923_),
    .Q(\count_instr[58] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30436_ (.D(_03924_),
    .Q(\count_instr[59] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30437_ (.D(_03925_),
    .Q(\count_instr[60] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30438_ (.D(_03926_),
    .Q(\count_instr[61] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30439_ (.D(_03927_),
    .Q(\count_instr[62] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30440_ (.D(_03928_),
    .Q(\count_instr[63] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _30441_ (.D(_03929_),
    .Q(\reg_pc[1] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _30442_ (.D(_03930_),
    .Q(\reg_pc[2] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30443_ (.D(_03931_),
    .Q(\reg_pc[3] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30444_ (.D(_03932_),
    .Q(\reg_pc[4] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30445_ (.D(_03933_),
    .Q(\reg_pc[5] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30446_ (.D(_03934_),
    .Q(\reg_pc[6] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _30447_ (.D(_03935_),
    .Q(\reg_pc[7] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30448_ (.D(_03936_),
    .Q(\reg_pc[8] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _30449_ (.D(_03937_),
    .Q(\reg_pc[9] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30450_ (.D(_03938_),
    .Q(\reg_pc[10] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30451_ (.D(_03939_),
    .Q(\reg_pc[11] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30452_ (.D(_03940_),
    .Q(\reg_pc[12] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30453_ (.D(_03941_),
    .Q(\reg_pc[13] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30454_ (.D(_03942_),
    .Q(\reg_pc[14] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30455_ (.D(_03943_),
    .Q(\reg_pc[15] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30456_ (.D(_03944_),
    .Q(\reg_pc[16] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _30457_ (.D(_03945_),
    .Q(\reg_pc[17] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30458_ (.D(_03946_),
    .Q(\reg_pc[18] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30459_ (.D(_03947_),
    .Q(\reg_pc[19] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _30460_ (.D(_03948_),
    .Q(\reg_pc[20] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30461_ (.D(_03949_),
    .Q(\reg_pc[21] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30462_ (.D(_03950_),
    .Q(\reg_pc[22] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30463_ (.D(_03951_),
    .Q(\reg_pc[23] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30464_ (.D(_03952_),
    .Q(\reg_pc[24] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30465_ (.D(_03953_),
    .Q(\reg_pc[25] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30466_ (.D(_03954_),
    .Q(\reg_pc[26] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30467_ (.D(_03955_),
    .Q(\reg_pc[27] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30468_ (.D(_03956_),
    .Q(\reg_pc[28] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30469_ (.D(_03957_),
    .Q(\reg_pc[29] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30470_ (.D(_03958_),
    .Q(\reg_pc[30] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30471_ (.D(_03959_),
    .Q(\reg_pc[31] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30472_ (.D(_03960_),
    .Q(\reg_next_pc[1] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _30473_ (.D(_03961_),
    .Q(\reg_next_pc[2] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30474_ (.D(_03962_),
    .Q(\reg_next_pc[3] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30475_ (.D(_03963_),
    .Q(\reg_next_pc[4] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30476_ (.D(_03964_),
    .Q(\reg_next_pc[5] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30477_ (.D(_03965_),
    .Q(\reg_next_pc[6] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30478_ (.D(_03966_),
    .Q(\reg_next_pc[7] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30479_ (.D(_03967_),
    .Q(\reg_next_pc[8] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30480_ (.D(_03968_),
    .Q(\reg_next_pc[9] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30481_ (.D(_03969_),
    .Q(\reg_next_pc[10] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30482_ (.D(_03970_),
    .Q(\reg_next_pc[11] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30483_ (.D(_03971_),
    .Q(\reg_next_pc[12] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30484_ (.D(_03972_),
    .Q(\reg_next_pc[13] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30485_ (.D(_03973_),
    .Q(\reg_next_pc[14] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30486_ (.D(_03974_),
    .Q(\reg_next_pc[15] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30487_ (.D(_03975_),
    .Q(\reg_next_pc[16] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30488_ (.D(_03976_),
    .Q(\reg_next_pc[17] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30489_ (.D(_03977_),
    .Q(\reg_next_pc[18] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30490_ (.D(_03978_),
    .Q(\reg_next_pc[19] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30491_ (.D(_03979_),
    .Q(\reg_next_pc[20] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30492_ (.D(_03980_),
    .Q(\reg_next_pc[21] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30493_ (.D(_03981_),
    .Q(\reg_next_pc[22] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30494_ (.D(_03982_),
    .Q(\reg_next_pc[23] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30495_ (.D(_03983_),
    .Q(\reg_next_pc[24] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30496_ (.D(_03984_),
    .Q(\reg_next_pc[25] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30497_ (.D(_03985_),
    .Q(\reg_next_pc[26] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30498_ (.D(_03986_),
    .Q(\reg_next_pc[27] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30499_ (.D(_03987_),
    .Q(\reg_next_pc[28] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30500_ (.D(_03988_),
    .Q(\reg_next_pc[29] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30501_ (.D(_03989_),
    .Q(\reg_next_pc[30] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30502_ (.D(_03990_),
    .Q(\reg_next_pc[31] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30503_ (.D(_03991_),
    .Q(mem_do_rdata),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30504_ (.D(_03992_),
    .Q(mem_do_wdata),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30505_ (.D(_03993_),
    .Q(\pcpi_timeout_counter[0] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30506_ (.D(_03994_),
    .Q(\pcpi_timeout_counter[1] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30507_ (.D(_03995_),
    .Q(\pcpi_timeout_counter[2] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30508_ (.D(_03996_),
    .Q(\pcpi_timeout_counter[3] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30509_ (.D(_03997_),
    .Q(instr_beq),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30510_ (.D(_03998_),
    .Q(instr_bne),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30511_ (.D(_03999_),
    .Q(instr_blt),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30512_ (.D(_04000_),
    .Q(instr_bge),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30513_ (.D(_04001_),
    .Q(instr_bltu),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30514_ (.D(_04002_),
    .Q(instr_bgeu),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30515_ (.D(_04003_),
    .Q(instr_addi),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30516_ (.D(_04004_),
    .Q(instr_slti),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30517_ (.D(_04005_),
    .Q(instr_sltiu),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30518_ (.D(_04006_),
    .Q(instr_xori),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _30519_ (.D(_04007_),
    .Q(instr_ori),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _30520_ (.D(_04008_),
    .Q(instr_andi),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30521_ (.D(_04009_),
    .Q(instr_add),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _30522_ (.D(_04010_),
    .Q(instr_sub),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30523_ (.D(_04011_),
    .Q(instr_sll),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30524_ (.D(_04012_),
    .Q(instr_slt),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30525_ (.D(_04013_),
    .Q(instr_sltu),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30526_ (.D(_04014_),
    .Q(instr_xor),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30527_ (.D(_04015_),
    .Q(instr_srl),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _30528_ (.D(_04016_),
    .Q(instr_sra),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _30529_ (.D(_04017_),
    .Q(instr_or),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _30530_ (.D(_04018_),
    .Q(instr_and),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30531_ (.D(_04019_),
    .Q(\decoded_rs1[0] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30532_ (.D(_04020_),
    .Q(\decoded_rs1[1] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30533_ (.D(_04021_),
    .Q(\decoded_rs1[2] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30534_ (.D(_04022_),
    .Q(\decoded_rs1[3] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30535_ (.D(_04023_),
    .Q(is_beq_bne_blt_bge_bltu_bgeu),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30536_ (.D(_04024_),
    .Q(net166),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30537_ (.D(_04025_),
    .Q(\irq_mask[0] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30538_ (.D(_04026_),
    .Q(\irq_mask[1] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30539_ (.D(_04027_),
    .Q(\irq_mask[2] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30540_ (.D(_04028_),
    .Q(\irq_mask[3] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30541_ (.D(_04029_),
    .Q(\irq_mask[4] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30542_ (.D(_04030_),
    .Q(\irq_mask[5] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30543_ (.D(_04031_),
    .Q(\irq_mask[6] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30544_ (.D(_04032_),
    .Q(\irq_mask[7] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30545_ (.D(_04033_),
    .Q(\irq_mask[8] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30546_ (.D(_04034_),
    .Q(\irq_mask[9] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30547_ (.D(_04035_),
    .Q(\irq_mask[10] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30548_ (.D(_04036_),
    .Q(\irq_mask[11] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30549_ (.D(_04037_),
    .Q(\irq_mask[12] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30550_ (.D(_04038_),
    .Q(\irq_mask[13] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30551_ (.D(_04039_),
    .Q(\irq_mask[14] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30552_ (.D(_04040_),
    .Q(\irq_mask[15] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30553_ (.D(_04041_),
    .Q(\irq_mask[16] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30554_ (.D(_04042_),
    .Q(\irq_mask[17] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30555_ (.D(_04043_),
    .Q(\irq_mask[18] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30556_ (.D(_04044_),
    .Q(\irq_mask[19] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30557_ (.D(_04045_),
    .Q(\irq_mask[20] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30558_ (.D(_04046_),
    .Q(\irq_mask[21] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30559_ (.D(_04047_),
    .Q(\irq_mask[22] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30560_ (.D(_04048_),
    .Q(\irq_mask[23] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30561_ (.D(_04049_),
    .Q(\irq_mask[24] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30562_ (.D(_04050_),
    .Q(\irq_mask[25] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30563_ (.D(_04051_),
    .Q(\irq_mask[26] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30564_ (.D(_04052_),
    .Q(\irq_mask[27] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30565_ (.D(_04053_),
    .Q(\irq_mask[28] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30566_ (.D(_04054_),
    .Q(\irq_mask[29] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30567_ (.D(_04055_),
    .Q(\irq_mask[30] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30568_ (.D(_04056_),
    .Q(\irq_mask[31] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30569_ (.D(_04057_),
    .Q(mem_do_prefetch),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30570_ (.D(_04058_),
    .Q(mem_do_rinst),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30571_ (.D(_04059_),
    .Q(\irq_state[0] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _30572_ (.D(_04060_),
    .Q(\irq_state[1] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _30573_ (.D(_04061_),
    .Q(latched_store),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _30574_ (.D(_04062_),
    .Q(latched_stalu),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _30575_ (.D(_04063_),
    .Q(\pcpi_mul.rs2[32] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30576_ (.D(_04064_),
    .Q(\pcpi_mul.rs1[32] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30577_ (.D(_04065_),
    .Q(irq_delay),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30578_ (.D(_04066_),
    .Q(\decoded_rs1[4] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30579_ (.D(_04067_),
    .Q(\mem_state[0] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30580_ (.D(_04068_),
    .Q(\mem_state[1] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30581_ (.D(_04069_),
    .Q(latched_branch),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _30582_ (.D(_04070_),
    .Q(latched_is_lh),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _30583_ (.D(_04071_),
    .Q(latched_is_lb),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30584_ (.D(_04072_),
    .Q(irq_active),
    .CLK(clk));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__decap_3 PHY_204 ();
 sky130_fd_sc_hd__decap_3 PHY_205 ();
 sky130_fd_sc_hd__decap_3 PHY_206 ();
 sky130_fd_sc_hd__decap_3 PHY_207 ();
 sky130_fd_sc_hd__decap_3 PHY_208 ();
 sky130_fd_sc_hd__decap_3 PHY_209 ();
 sky130_fd_sc_hd__decap_3 PHY_210 ();
 sky130_fd_sc_hd__decap_3 PHY_211 ();
 sky130_fd_sc_hd__decap_3 PHY_212 ();
 sky130_fd_sc_hd__decap_3 PHY_213 ();
 sky130_fd_sc_hd__decap_3 PHY_214 ();
 sky130_fd_sc_hd__decap_3 PHY_215 ();
 sky130_fd_sc_hd__decap_3 PHY_216 ();
 sky130_fd_sc_hd__decap_3 PHY_217 ();
 sky130_fd_sc_hd__decap_3 PHY_218 ();
 sky130_fd_sc_hd__decap_3 PHY_219 ();
 sky130_fd_sc_hd__decap_3 PHY_220 ();
 sky130_fd_sc_hd__decap_3 PHY_221 ();
 sky130_fd_sc_hd__decap_3 PHY_222 ();
 sky130_fd_sc_hd__decap_3 PHY_223 ();
 sky130_fd_sc_hd__decap_3 PHY_224 ();
 sky130_fd_sc_hd__decap_3 PHY_225 ();
 sky130_fd_sc_hd__decap_3 PHY_226 ();
 sky130_fd_sc_hd__decap_3 PHY_227 ();
 sky130_fd_sc_hd__decap_3 PHY_228 ();
 sky130_fd_sc_hd__decap_3 PHY_229 ();
 sky130_fd_sc_hd__decap_3 PHY_230 ();
 sky130_fd_sc_hd__decap_3 PHY_231 ();
 sky130_fd_sc_hd__decap_3 PHY_232 ();
 sky130_fd_sc_hd__decap_3 PHY_233 ();
 sky130_fd_sc_hd__decap_3 PHY_234 ();
 sky130_fd_sc_hd__decap_3 PHY_235 ();
 sky130_fd_sc_hd__decap_3 PHY_236 ();
 sky130_fd_sc_hd__decap_3 PHY_237 ();
 sky130_fd_sc_hd__decap_3 PHY_238 ();
 sky130_fd_sc_hd__decap_3 PHY_239 ();
 sky130_fd_sc_hd__decap_3 PHY_240 ();
 sky130_fd_sc_hd__decap_3 PHY_241 ();
 sky130_fd_sc_hd__decap_3 PHY_242 ();
 sky130_fd_sc_hd__decap_3 PHY_243 ();
 sky130_fd_sc_hd__decap_3 PHY_244 ();
 sky130_fd_sc_hd__decap_3 PHY_245 ();
 sky130_fd_sc_hd__decap_3 PHY_246 ();
 sky130_fd_sc_hd__decap_3 PHY_247 ();
 sky130_fd_sc_hd__decap_3 PHY_248 ();
 sky130_fd_sc_hd__decap_3 PHY_249 ();
 sky130_fd_sc_hd__decap_3 PHY_250 ();
 sky130_fd_sc_hd__decap_3 PHY_251 ();
 sky130_fd_sc_hd__decap_3 PHY_252 ();
 sky130_fd_sc_hd__decap_3 PHY_253 ();
 sky130_fd_sc_hd__decap_3 PHY_254 ();
 sky130_fd_sc_hd__decap_3 PHY_255 ();
 sky130_fd_sc_hd__decap_3 PHY_256 ();
 sky130_fd_sc_hd__decap_3 PHY_257 ();
 sky130_fd_sc_hd__decap_3 PHY_258 ();
 sky130_fd_sc_hd__decap_3 PHY_259 ();
 sky130_fd_sc_hd__decap_3 PHY_260 ();
 sky130_fd_sc_hd__decap_3 PHY_261 ();
 sky130_fd_sc_hd__decap_3 PHY_262 ();
 sky130_fd_sc_hd__decap_3 PHY_263 ();
 sky130_fd_sc_hd__decap_3 PHY_264 ();
 sky130_fd_sc_hd__decap_3 PHY_265 ();
 sky130_fd_sc_hd__decap_3 PHY_266 ();
 sky130_fd_sc_hd__decap_3 PHY_267 ();
 sky130_fd_sc_hd__decap_3 PHY_268 ();
 sky130_fd_sc_hd__decap_3 PHY_269 ();
 sky130_fd_sc_hd__decap_3 PHY_270 ();
 sky130_fd_sc_hd__decap_3 PHY_271 ();
 sky130_fd_sc_hd__decap_3 PHY_272 ();
 sky130_fd_sc_hd__decap_3 PHY_273 ();
 sky130_fd_sc_hd__decap_3 PHY_274 ();
 sky130_fd_sc_hd__decap_3 PHY_275 ();
 sky130_fd_sc_hd__decap_3 PHY_276 ();
 sky130_fd_sc_hd__decap_3 PHY_277 ();
 sky130_fd_sc_hd__decap_3 PHY_278 ();
 sky130_fd_sc_hd__decap_3 PHY_279 ();
 sky130_fd_sc_hd__decap_3 PHY_280 ();
 sky130_fd_sc_hd__decap_3 PHY_281 ();
 sky130_fd_sc_hd__decap_3 PHY_282 ();
 sky130_fd_sc_hd__decap_3 PHY_283 ();
 sky130_fd_sc_hd__decap_3 PHY_284 ();
 sky130_fd_sc_hd__decap_3 PHY_285 ();
 sky130_fd_sc_hd__decap_3 PHY_286 ();
 sky130_fd_sc_hd__decap_3 PHY_287 ();
 sky130_fd_sc_hd__decap_3 PHY_288 ();
 sky130_fd_sc_hd__decap_3 PHY_289 ();
 sky130_fd_sc_hd__decap_3 PHY_290 ();
 sky130_fd_sc_hd__decap_3 PHY_291 ();
 sky130_fd_sc_hd__decap_3 PHY_292 ();
 sky130_fd_sc_hd__decap_3 PHY_293 ();
 sky130_fd_sc_hd__decap_3 PHY_294 ();
 sky130_fd_sc_hd__decap_3 PHY_295 ();
 sky130_fd_sc_hd__decap_3 PHY_296 ();
 sky130_fd_sc_hd__decap_3 PHY_297 ();
 sky130_fd_sc_hd__decap_3 PHY_298 ();
 sky130_fd_sc_hd__decap_3 PHY_299 ();
 sky130_fd_sc_hd__decap_3 PHY_300 ();
 sky130_fd_sc_hd__decap_3 PHY_301 ();
 sky130_fd_sc_hd__decap_3 PHY_302 ();
 sky130_fd_sc_hd__decap_3 PHY_303 ();
 sky130_fd_sc_hd__decap_3 PHY_304 ();
 sky130_fd_sc_hd__decap_3 PHY_305 ();
 sky130_fd_sc_hd__decap_3 PHY_306 ();
 sky130_fd_sc_hd__decap_3 PHY_307 ();
 sky130_fd_sc_hd__decap_3 PHY_308 ();
 sky130_fd_sc_hd__decap_3 PHY_309 ();
 sky130_fd_sc_hd__decap_3 PHY_310 ();
 sky130_fd_sc_hd__decap_3 PHY_311 ();
 sky130_fd_sc_hd__decap_3 PHY_312 ();
 sky130_fd_sc_hd__decap_3 PHY_313 ();
 sky130_fd_sc_hd__decap_3 PHY_314 ();
 sky130_fd_sc_hd__decap_3 PHY_315 ();
 sky130_fd_sc_hd__decap_3 PHY_316 ();
 sky130_fd_sc_hd__decap_3 PHY_317 ();
 sky130_fd_sc_hd__decap_3 PHY_318 ();
 sky130_fd_sc_hd__decap_3 PHY_319 ();
 sky130_fd_sc_hd__decap_3 PHY_320 ();
 sky130_fd_sc_hd__decap_3 PHY_321 ();
 sky130_fd_sc_hd__decap_3 PHY_322 ();
 sky130_fd_sc_hd__decap_3 PHY_323 ();
 sky130_fd_sc_hd__decap_3 PHY_324 ();
 sky130_fd_sc_hd__decap_3 PHY_325 ();
 sky130_fd_sc_hd__decap_3 PHY_326 ();
 sky130_fd_sc_hd__decap_3 PHY_327 ();
 sky130_fd_sc_hd__decap_3 PHY_328 ();
 sky130_fd_sc_hd__decap_3 PHY_329 ();
 sky130_fd_sc_hd__decap_3 PHY_330 ();
 sky130_fd_sc_hd__decap_3 PHY_331 ();
 sky130_fd_sc_hd__decap_3 PHY_332 ();
 sky130_fd_sc_hd__decap_3 PHY_333 ();
 sky130_fd_sc_hd__decap_3 PHY_334 ();
 sky130_fd_sc_hd__decap_3 PHY_335 ();
 sky130_fd_sc_hd__decap_3 PHY_336 ();
 sky130_fd_sc_hd__decap_3 PHY_337 ();
 sky130_fd_sc_hd__decap_3 PHY_338 ();
 sky130_fd_sc_hd__decap_3 PHY_339 ();
 sky130_fd_sc_hd__decap_3 PHY_340 ();
 sky130_fd_sc_hd__decap_3 PHY_341 ();
 sky130_fd_sc_hd__decap_3 PHY_342 ();
 sky130_fd_sc_hd__decap_3 PHY_343 ();
 sky130_fd_sc_hd__decap_3 PHY_344 ();
 sky130_fd_sc_hd__decap_3 PHY_345 ();
 sky130_fd_sc_hd__decap_3 PHY_346 ();
 sky130_fd_sc_hd__decap_3 PHY_347 ();
 sky130_fd_sc_hd__decap_3 PHY_348 ();
 sky130_fd_sc_hd__decap_3 PHY_349 ();
 sky130_fd_sc_hd__decap_3 PHY_350 ();
 sky130_fd_sc_hd__decap_3 PHY_351 ();
 sky130_fd_sc_hd__decap_3 PHY_352 ();
 sky130_fd_sc_hd__decap_3 PHY_353 ();
 sky130_fd_sc_hd__decap_3 PHY_354 ();
 sky130_fd_sc_hd__decap_3 PHY_355 ();
 sky130_fd_sc_hd__decap_3 PHY_356 ();
 sky130_fd_sc_hd__decap_3 PHY_357 ();
 sky130_fd_sc_hd__decap_3 PHY_358 ();
 sky130_fd_sc_hd__decap_3 PHY_359 ();
 sky130_fd_sc_hd__decap_3 PHY_360 ();
 sky130_fd_sc_hd__decap_3 PHY_361 ();
 sky130_fd_sc_hd__decap_3 PHY_362 ();
 sky130_fd_sc_hd__decap_3 PHY_363 ();
 sky130_fd_sc_hd__decap_3 PHY_364 ();
 sky130_fd_sc_hd__decap_3 PHY_365 ();
 sky130_fd_sc_hd__decap_3 PHY_366 ();
 sky130_fd_sc_hd__decap_3 PHY_367 ();
 sky130_fd_sc_hd__decap_3 PHY_368 ();
 sky130_fd_sc_hd__decap_3 PHY_369 ();
 sky130_fd_sc_hd__decap_3 PHY_370 ();
 sky130_fd_sc_hd__decap_3 PHY_371 ();
 sky130_fd_sc_hd__decap_3 PHY_372 ();
 sky130_fd_sc_hd__decap_3 PHY_373 ();
 sky130_fd_sc_hd__decap_3 PHY_374 ();
 sky130_fd_sc_hd__decap_3 PHY_375 ();
 sky130_fd_sc_hd__decap_3 PHY_376 ();
 sky130_fd_sc_hd__decap_3 PHY_377 ();
 sky130_fd_sc_hd__decap_3 PHY_378 ();
 sky130_fd_sc_hd__decap_3 PHY_379 ();
 sky130_fd_sc_hd__decap_3 PHY_380 ();
 sky130_fd_sc_hd__decap_3 PHY_381 ();
 sky130_fd_sc_hd__decap_3 PHY_382 ();
 sky130_fd_sc_hd__decap_3 PHY_383 ();
 sky130_fd_sc_hd__decap_3 PHY_384 ();
 sky130_fd_sc_hd__decap_3 PHY_385 ();
 sky130_fd_sc_hd__decap_3 PHY_386 ();
 sky130_fd_sc_hd__decap_3 PHY_387 ();
 sky130_fd_sc_hd__decap_3 PHY_388 ();
 sky130_fd_sc_hd__decap_3 PHY_389 ();
 sky130_fd_sc_hd__decap_3 PHY_390 ();
 sky130_fd_sc_hd__decap_3 PHY_391 ();
 sky130_fd_sc_hd__decap_3 PHY_392 ();
 sky130_fd_sc_hd__decap_3 PHY_393 ();
 sky130_fd_sc_hd__decap_3 PHY_394 ();
 sky130_fd_sc_hd__decap_3 PHY_395 ();
 sky130_fd_sc_hd__decap_3 PHY_396 ();
 sky130_fd_sc_hd__decap_3 PHY_397 ();
 sky130_fd_sc_hd__decap_3 PHY_398 ();
 sky130_fd_sc_hd__decap_3 PHY_399 ();
 sky130_fd_sc_hd__decap_3 PHY_400 ();
 sky130_fd_sc_hd__decap_3 PHY_401 ();
 sky130_fd_sc_hd__decap_3 PHY_402 ();
 sky130_fd_sc_hd__decap_3 PHY_403 ();
 sky130_fd_sc_hd__decap_3 PHY_404 ();
 sky130_fd_sc_hd__decap_3 PHY_405 ();
 sky130_fd_sc_hd__decap_3 PHY_406 ();
 sky130_fd_sc_hd__decap_3 PHY_407 ();
 sky130_fd_sc_hd__decap_3 PHY_408 ();
 sky130_fd_sc_hd__decap_3 PHY_409 ();
 sky130_fd_sc_hd__decap_3 PHY_410 ();
 sky130_fd_sc_hd__decap_3 PHY_411 ();
 sky130_fd_sc_hd__decap_3 PHY_412 ();
 sky130_fd_sc_hd__decap_3 PHY_413 ();
 sky130_fd_sc_hd__decap_3 PHY_414 ();
 sky130_fd_sc_hd__decap_3 PHY_415 ();
 sky130_fd_sc_hd__decap_3 PHY_416 ();
 sky130_fd_sc_hd__decap_3 PHY_417 ();
 sky130_fd_sc_hd__decap_3 PHY_418 ();
 sky130_fd_sc_hd__decap_3 PHY_419 ();
 sky130_fd_sc_hd__decap_3 PHY_420 ();
 sky130_fd_sc_hd__decap_3 PHY_421 ();
 sky130_fd_sc_hd__decap_3 PHY_422 ();
 sky130_fd_sc_hd__decap_3 PHY_423 ();
 sky130_fd_sc_hd__decap_3 PHY_424 ();
 sky130_fd_sc_hd__decap_3 PHY_425 ();
 sky130_fd_sc_hd__decap_3 PHY_426 ();
 sky130_fd_sc_hd__decap_3 PHY_427 ();
 sky130_fd_sc_hd__decap_3 PHY_428 ();
 sky130_fd_sc_hd__decap_3 PHY_429 ();
 sky130_fd_sc_hd__decap_3 PHY_430 ();
 sky130_fd_sc_hd__decap_3 PHY_431 ();
 sky130_fd_sc_hd__decap_3 PHY_432 ();
 sky130_fd_sc_hd__decap_3 PHY_433 ();
 sky130_fd_sc_hd__decap_3 PHY_434 ();
 sky130_fd_sc_hd__decap_3 PHY_435 ();
 sky130_fd_sc_hd__decap_3 PHY_436 ();
 sky130_fd_sc_hd__decap_3 PHY_437 ();
 sky130_fd_sc_hd__decap_3 PHY_438 ();
 sky130_fd_sc_hd__decap_3 PHY_439 ();
 sky130_fd_sc_hd__decap_3 PHY_440 ();
 sky130_fd_sc_hd__decap_3 PHY_441 ();
 sky130_fd_sc_hd__decap_3 PHY_442 ();
 sky130_fd_sc_hd__decap_3 PHY_443 ();
 sky130_fd_sc_hd__decap_3 PHY_444 ();
 sky130_fd_sc_hd__decap_3 PHY_445 ();
 sky130_fd_sc_hd__decap_3 PHY_446 ();
 sky130_fd_sc_hd__decap_3 PHY_447 ();
 sky130_fd_sc_hd__decap_3 PHY_448 ();
 sky130_fd_sc_hd__decap_3 PHY_449 ();
 sky130_fd_sc_hd__decap_3 PHY_450 ();
 sky130_fd_sc_hd__decap_3 PHY_451 ();
 sky130_fd_sc_hd__decap_3 PHY_452 ();
 sky130_fd_sc_hd__decap_3 PHY_453 ();
 sky130_fd_sc_hd__decap_3 PHY_454 ();
 sky130_fd_sc_hd__decap_3 PHY_455 ();
 sky130_fd_sc_hd__decap_3 PHY_456 ();
 sky130_fd_sc_hd__decap_3 PHY_457 ();
 sky130_fd_sc_hd__decap_3 PHY_458 ();
 sky130_fd_sc_hd__decap_3 PHY_459 ();
 sky130_fd_sc_hd__decap_3 PHY_460 ();
 sky130_fd_sc_hd__decap_3 PHY_461 ();
 sky130_fd_sc_hd__decap_3 PHY_462 ();
 sky130_fd_sc_hd__decap_3 PHY_463 ();
 sky130_fd_sc_hd__decap_3 PHY_464 ();
 sky130_fd_sc_hd__decap_3 PHY_465 ();
 sky130_fd_sc_hd__decap_3 PHY_466 ();
 sky130_fd_sc_hd__decap_3 PHY_467 ();
 sky130_fd_sc_hd__decap_3 PHY_468 ();
 sky130_fd_sc_hd__decap_3 PHY_469 ();
 sky130_fd_sc_hd__decap_3 PHY_470 ();
 sky130_fd_sc_hd__decap_3 PHY_471 ();
 sky130_fd_sc_hd__decap_3 PHY_472 ();
 sky130_fd_sc_hd__decap_3 PHY_473 ();
 sky130_fd_sc_hd__decap_3 PHY_474 ();
 sky130_fd_sc_hd__decap_3 PHY_475 ();
 sky130_fd_sc_hd__decap_3 PHY_476 ();
 sky130_fd_sc_hd__decap_3 PHY_477 ();
 sky130_fd_sc_hd__decap_3 PHY_478 ();
 sky130_fd_sc_hd__decap_3 PHY_479 ();
 sky130_fd_sc_hd__decap_3 PHY_480 ();
 sky130_fd_sc_hd__decap_3 PHY_481 ();
 sky130_fd_sc_hd__decap_3 PHY_482 ();
 sky130_fd_sc_hd__decap_3 PHY_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6581 ();
 sky130_fd_sc_hd__buf_6 input1 (.A(irq[0]),
    .X(net1));
 sky130_fd_sc_hd__buf_8 input2 (.A(irq[10]),
    .X(net2));
 sky130_fd_sc_hd__buf_4 input3 (.A(irq[11]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_4 input4 (.A(irq[12]),
    .X(net4));
 sky130_fd_sc_hd__buf_6 input5 (.A(irq[13]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_4 input6 (.A(irq[14]),
    .X(net6));
 sky130_fd_sc_hd__buf_8 input7 (.A(irq[15]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_4 input8 (.A(irq[16]),
    .X(net8));
 sky130_fd_sc_hd__buf_4 input9 (.A(irq[17]),
    .X(net9));
 sky130_fd_sc_hd__buf_1 input10 (.A(irq[18]),
    .X(net10));
 sky130_fd_sc_hd__buf_1 input11 (.A(irq[19]),
    .X(net11));
 sky130_fd_sc_hd__buf_4 input12 (.A(irq[1]),
    .X(net12));
 sky130_fd_sc_hd__buf_1 input13 (.A(irq[20]),
    .X(net13));
 sky130_fd_sc_hd__buf_8 input14 (.A(irq[21]),
    .X(net14));
 sky130_fd_sc_hd__buf_1 input15 (.A(irq[22]),
    .X(net15));
 sky130_fd_sc_hd__buf_2 input16 (.A(irq[23]),
    .X(net16));
 sky130_fd_sc_hd__buf_4 input17 (.A(irq[24]),
    .X(net17));
 sky130_fd_sc_hd__buf_4 input18 (.A(irq[25]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_4 input19 (.A(irq[26]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_2 input20 (.A(irq[27]),
    .X(net20));
 sky130_fd_sc_hd__buf_1 input21 (.A(irq[28]),
    .X(net21));
 sky130_fd_sc_hd__buf_4 input22 (.A(irq[29]),
    .X(net22));
 sky130_fd_sc_hd__buf_6 input23 (.A(irq[2]),
    .X(net23));
 sky130_fd_sc_hd__buf_4 input24 (.A(irq[30]),
    .X(net24));
 sky130_fd_sc_hd__buf_6 input25 (.A(irq[31]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_4 input26 (.A(irq[3]),
    .X(net26));
 sky130_fd_sc_hd__buf_6 input27 (.A(irq[4]),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_4 input28 (.A(irq[5]),
    .X(net28));
 sky130_fd_sc_hd__buf_6 input29 (.A(irq[6]),
    .X(net29));
 sky130_fd_sc_hd__buf_8 input30 (.A(irq[7]),
    .X(net30));
 sky130_fd_sc_hd__buf_2 input31 (.A(irq[8]),
    .X(net31));
 sky130_fd_sc_hd__buf_6 input32 (.A(irq[9]),
    .X(net32));
 sky130_fd_sc_hd__buf_6 input33 (.A(mem_rdata[0]),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_4 input34 (.A(mem_rdata[10]),
    .X(net34));
 sky130_fd_sc_hd__buf_6 input35 (.A(mem_rdata[11]),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_8 input36 (.A(mem_rdata[12]),
    .X(net36));
 sky130_fd_sc_hd__buf_4 input37 (.A(mem_rdata[13]),
    .X(net37));
 sky130_fd_sc_hd__buf_6 input38 (.A(mem_rdata[14]),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_8 input39 (.A(mem_rdata[15]),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_4 input40 (.A(mem_rdata[16]),
    .X(net40));
 sky130_fd_sc_hd__buf_6 input41 (.A(mem_rdata[17]),
    .X(net41));
 sky130_fd_sc_hd__buf_6 input42 (.A(mem_rdata[18]),
    .X(net42));
 sky130_fd_sc_hd__buf_6 input43 (.A(mem_rdata[19]),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_8 input44 (.A(mem_rdata[1]),
    .X(net44));
 sky130_fd_sc_hd__buf_1 input45 (.A(mem_rdata[20]),
    .X(net45));
 sky130_fd_sc_hd__buf_4 input46 (.A(mem_rdata[21]),
    .X(net46));
 sky130_fd_sc_hd__buf_4 input47 (.A(mem_rdata[22]),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_4 input48 (.A(mem_rdata[23]),
    .X(net48));
 sky130_fd_sc_hd__buf_4 input49 (.A(mem_rdata[24]),
    .X(net49));
 sky130_fd_sc_hd__buf_6 input50 (.A(mem_rdata[25]),
    .X(net50));
 sky130_fd_sc_hd__buf_4 input51 (.A(mem_rdata[26]),
    .X(net51));
 sky130_fd_sc_hd__buf_6 input52 (.A(mem_rdata[27]),
    .X(net52));
 sky130_fd_sc_hd__buf_4 input53 (.A(mem_rdata[28]),
    .X(net53));
 sky130_fd_sc_hd__buf_6 input54 (.A(mem_rdata[29]),
    .X(net54));
 sky130_fd_sc_hd__buf_6 input55 (.A(mem_rdata[2]),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_8 input56 (.A(mem_rdata[30]),
    .X(net56));
 sky130_fd_sc_hd__buf_6 input57 (.A(mem_rdata[31]),
    .X(net57));
 sky130_fd_sc_hd__buf_6 input58 (.A(mem_rdata[3]),
    .X(net58));
 sky130_fd_sc_hd__buf_6 input59 (.A(mem_rdata[4]),
    .X(net59));
 sky130_fd_sc_hd__buf_6 input60 (.A(mem_rdata[5]),
    .X(net60));
 sky130_fd_sc_hd__buf_6 input61 (.A(mem_rdata[6]),
    .X(net61));
 sky130_fd_sc_hd__buf_4 input62 (.A(mem_rdata[7]),
    .X(net62));
 sky130_fd_sc_hd__buf_6 input63 (.A(mem_rdata[8]),
    .X(net63));
 sky130_fd_sc_hd__clkbuf_4 input64 (.A(mem_rdata[9]),
    .X(net64));
 sky130_fd_sc_hd__buf_8 input65 (.A(mem_ready),
    .X(net65));
 sky130_fd_sc_hd__buf_1 input66 (.A(pcpi_rd[0]),
    .X(net66));
 sky130_fd_sc_hd__buf_1 input67 (.A(pcpi_rd[10]),
    .X(net67));
 sky130_fd_sc_hd__buf_1 input68 (.A(pcpi_rd[11]),
    .X(net68));
 sky130_fd_sc_hd__buf_1 input69 (.A(pcpi_rd[12]),
    .X(net69));
 sky130_fd_sc_hd__buf_1 input70 (.A(pcpi_rd[13]),
    .X(net70));
 sky130_fd_sc_hd__buf_1 input71 (.A(pcpi_rd[14]),
    .X(net71));
 sky130_fd_sc_hd__buf_1 input72 (.A(pcpi_rd[15]),
    .X(net72));
 sky130_fd_sc_hd__buf_1 input73 (.A(pcpi_rd[16]),
    .X(net73));
 sky130_fd_sc_hd__buf_1 input74 (.A(pcpi_rd[17]),
    .X(net74));
 sky130_fd_sc_hd__buf_1 input75 (.A(pcpi_rd[18]),
    .X(net75));
 sky130_fd_sc_hd__buf_1 input76 (.A(pcpi_rd[19]),
    .X(net76));
 sky130_fd_sc_hd__buf_1 input77 (.A(pcpi_rd[1]),
    .X(net77));
 sky130_fd_sc_hd__buf_1 input78 (.A(pcpi_rd[20]),
    .X(net78));
 sky130_fd_sc_hd__buf_1 input79 (.A(pcpi_rd[21]),
    .X(net79));
 sky130_fd_sc_hd__buf_1 input80 (.A(pcpi_rd[22]),
    .X(net80));
 sky130_fd_sc_hd__buf_1 input81 (.A(pcpi_rd[23]),
    .X(net81));
 sky130_fd_sc_hd__buf_1 input82 (.A(pcpi_rd[24]),
    .X(net82));
 sky130_fd_sc_hd__buf_1 input83 (.A(pcpi_rd[25]),
    .X(net83));
 sky130_fd_sc_hd__buf_1 input84 (.A(pcpi_rd[26]),
    .X(net84));
 sky130_fd_sc_hd__buf_1 input85 (.A(pcpi_rd[27]),
    .X(net85));
 sky130_fd_sc_hd__buf_1 input86 (.A(pcpi_rd[28]),
    .X(net86));
 sky130_fd_sc_hd__buf_1 input87 (.A(pcpi_rd[29]),
    .X(net87));
 sky130_fd_sc_hd__buf_1 input88 (.A(pcpi_rd[2]),
    .X(net88));
 sky130_fd_sc_hd__buf_1 input89 (.A(pcpi_rd[30]),
    .X(net89));
 sky130_fd_sc_hd__buf_1 input90 (.A(pcpi_rd[31]),
    .X(net90));
 sky130_fd_sc_hd__buf_1 input91 (.A(pcpi_rd[3]),
    .X(net91));
 sky130_fd_sc_hd__buf_1 input92 (.A(pcpi_rd[4]),
    .X(net92));
 sky130_fd_sc_hd__buf_1 input93 (.A(pcpi_rd[5]),
    .X(net93));
 sky130_fd_sc_hd__buf_1 input94 (.A(pcpi_rd[6]),
    .X(net94));
 sky130_fd_sc_hd__buf_1 input95 (.A(pcpi_rd[7]),
    .X(net95));
 sky130_fd_sc_hd__buf_1 input96 (.A(pcpi_rd[8]),
    .X(net96));
 sky130_fd_sc_hd__buf_1 input97 (.A(pcpi_rd[9]),
    .X(net97));
 sky130_fd_sc_hd__buf_1 input98 (.A(pcpi_ready),
    .X(net98));
 sky130_fd_sc_hd__buf_1 input99 (.A(pcpi_wait),
    .X(net99));
 sky130_fd_sc_hd__buf_1 input100 (.A(pcpi_wr),
    .X(net100));
 sky130_fd_sc_hd__buf_4 input101 (.A(resetn),
    .X(net101));
 sky130_fd_sc_hd__clkbuf_2 output102 (.A(net102),
    .X(eoi[0]));
 sky130_fd_sc_hd__clkbuf_2 output103 (.A(net103),
    .X(eoi[10]));
 sky130_fd_sc_hd__clkbuf_2 output104 (.A(net104),
    .X(eoi[11]));
 sky130_fd_sc_hd__clkbuf_2 output105 (.A(net105),
    .X(eoi[12]));
 sky130_fd_sc_hd__clkbuf_2 output106 (.A(net106),
    .X(eoi[13]));
 sky130_fd_sc_hd__clkbuf_2 output107 (.A(net107),
    .X(eoi[14]));
 sky130_fd_sc_hd__clkbuf_2 output108 (.A(net108),
    .X(eoi[15]));
 sky130_fd_sc_hd__clkbuf_2 output109 (.A(net109),
    .X(eoi[16]));
 sky130_fd_sc_hd__clkbuf_2 output110 (.A(net110),
    .X(eoi[17]));
 sky130_fd_sc_hd__clkbuf_2 output111 (.A(net111),
    .X(eoi[18]));
 sky130_fd_sc_hd__clkbuf_2 output112 (.A(net112),
    .X(eoi[19]));
 sky130_fd_sc_hd__clkbuf_2 output113 (.A(net113),
    .X(eoi[1]));
 sky130_fd_sc_hd__clkbuf_2 output114 (.A(net114),
    .X(eoi[20]));
 sky130_fd_sc_hd__clkbuf_2 output115 (.A(net115),
    .X(eoi[21]));
 sky130_fd_sc_hd__clkbuf_2 output116 (.A(net116),
    .X(eoi[22]));
 sky130_fd_sc_hd__clkbuf_2 output117 (.A(net117),
    .X(eoi[23]));
 sky130_fd_sc_hd__clkbuf_2 output118 (.A(net118),
    .X(eoi[24]));
 sky130_fd_sc_hd__clkbuf_2 output119 (.A(net119),
    .X(eoi[25]));
 sky130_fd_sc_hd__clkbuf_2 output120 (.A(net120),
    .X(eoi[26]));
 sky130_fd_sc_hd__clkbuf_2 output121 (.A(net121),
    .X(eoi[27]));
 sky130_fd_sc_hd__clkbuf_2 output122 (.A(net122),
    .X(eoi[28]));
 sky130_fd_sc_hd__clkbuf_2 output123 (.A(net123),
    .X(eoi[29]));
 sky130_fd_sc_hd__clkbuf_2 output124 (.A(net124),
    .X(eoi[2]));
 sky130_fd_sc_hd__clkbuf_2 output125 (.A(net125),
    .X(eoi[30]));
 sky130_fd_sc_hd__clkbuf_2 output126 (.A(net126),
    .X(eoi[31]));
 sky130_fd_sc_hd__clkbuf_2 output127 (.A(net127),
    .X(eoi[3]));
 sky130_fd_sc_hd__clkbuf_2 output128 (.A(net128),
    .X(eoi[4]));
 sky130_fd_sc_hd__clkbuf_2 output129 (.A(net129),
    .X(eoi[5]));
 sky130_fd_sc_hd__clkbuf_2 output130 (.A(net130),
    .X(eoi[6]));
 sky130_fd_sc_hd__clkbuf_2 output131 (.A(net131),
    .X(eoi[7]));
 sky130_fd_sc_hd__clkbuf_2 output132 (.A(net132),
    .X(eoi[8]));
 sky130_fd_sc_hd__clkbuf_2 output133 (.A(net133),
    .X(eoi[9]));
 sky130_fd_sc_hd__clkbuf_2 output134 (.A(net134),
    .X(mem_addr[0]));
 sky130_fd_sc_hd__clkbuf_2 output135 (.A(net135),
    .X(mem_addr[10]));
 sky130_fd_sc_hd__clkbuf_2 output136 (.A(net136),
    .X(mem_addr[11]));
 sky130_fd_sc_hd__clkbuf_2 output137 (.A(net137),
    .X(mem_addr[12]));
 sky130_fd_sc_hd__clkbuf_2 output138 (.A(net138),
    .X(mem_addr[13]));
 sky130_fd_sc_hd__clkbuf_2 output139 (.A(net139),
    .X(mem_addr[14]));
 sky130_fd_sc_hd__clkbuf_2 output140 (.A(net140),
    .X(mem_addr[15]));
 sky130_fd_sc_hd__clkbuf_2 output141 (.A(net141),
    .X(mem_addr[16]));
 sky130_fd_sc_hd__clkbuf_2 output142 (.A(net142),
    .X(mem_addr[17]));
 sky130_fd_sc_hd__clkbuf_2 output143 (.A(net143),
    .X(mem_addr[18]));
 sky130_fd_sc_hd__clkbuf_2 output144 (.A(net144),
    .X(mem_addr[19]));
 sky130_fd_sc_hd__clkbuf_2 output145 (.A(net145),
    .X(mem_addr[1]));
 sky130_fd_sc_hd__clkbuf_2 output146 (.A(net146),
    .X(mem_addr[20]));
 sky130_fd_sc_hd__clkbuf_2 output147 (.A(net147),
    .X(mem_addr[21]));
 sky130_fd_sc_hd__clkbuf_2 output148 (.A(net148),
    .X(mem_addr[22]));
 sky130_fd_sc_hd__clkbuf_2 output149 (.A(net149),
    .X(mem_addr[23]));
 sky130_fd_sc_hd__clkbuf_2 output150 (.A(net150),
    .X(mem_addr[24]));
 sky130_fd_sc_hd__clkbuf_2 output151 (.A(net151),
    .X(mem_addr[25]));
 sky130_fd_sc_hd__clkbuf_2 output152 (.A(net152),
    .X(mem_addr[26]));
 sky130_fd_sc_hd__clkbuf_2 output153 (.A(net153),
    .X(mem_addr[27]));
 sky130_fd_sc_hd__clkbuf_2 output154 (.A(net154),
    .X(mem_addr[28]));
 sky130_fd_sc_hd__clkbuf_2 output155 (.A(net155),
    .X(mem_addr[29]));
 sky130_fd_sc_hd__clkbuf_2 output156 (.A(net156),
    .X(mem_addr[2]));
 sky130_fd_sc_hd__clkbuf_2 output157 (.A(net157),
    .X(mem_addr[30]));
 sky130_fd_sc_hd__clkbuf_2 output158 (.A(net158),
    .X(mem_addr[31]));
 sky130_fd_sc_hd__clkbuf_2 output159 (.A(net159),
    .X(mem_addr[3]));
 sky130_fd_sc_hd__clkbuf_2 output160 (.A(net160),
    .X(mem_addr[4]));
 sky130_fd_sc_hd__clkbuf_2 output161 (.A(net161),
    .X(mem_addr[5]));
 sky130_fd_sc_hd__clkbuf_2 output162 (.A(net162),
    .X(mem_addr[6]));
 sky130_fd_sc_hd__clkbuf_2 output163 (.A(net163),
    .X(mem_addr[7]));
 sky130_fd_sc_hd__clkbuf_2 output164 (.A(net164),
    .X(mem_addr[8]));
 sky130_fd_sc_hd__clkbuf_2 output165 (.A(net165),
    .X(mem_addr[9]));
 sky130_fd_sc_hd__clkbuf_2 output166 (.A(net166),
    .X(mem_instr));
 sky130_fd_sc_hd__clkbuf_2 output167 (.A(net167),
    .X(mem_la_addr[0]));
 sky130_fd_sc_hd__clkbuf_2 output168 (.A(net168),
    .X(mem_la_addr[10]));
 sky130_fd_sc_hd__clkbuf_2 output169 (.A(net169),
    .X(mem_la_addr[11]));
 sky130_fd_sc_hd__clkbuf_2 output170 (.A(net170),
    .X(mem_la_addr[12]));
 sky130_fd_sc_hd__clkbuf_2 output171 (.A(net171),
    .X(mem_la_addr[13]));
 sky130_fd_sc_hd__clkbuf_2 output172 (.A(net172),
    .X(mem_la_addr[14]));
 sky130_fd_sc_hd__clkbuf_2 output173 (.A(net173),
    .X(mem_la_addr[15]));
 sky130_fd_sc_hd__clkbuf_2 output174 (.A(net174),
    .X(mem_la_addr[16]));
 sky130_fd_sc_hd__clkbuf_2 output175 (.A(net175),
    .X(mem_la_addr[17]));
 sky130_fd_sc_hd__clkbuf_2 output176 (.A(net176),
    .X(mem_la_addr[18]));
 sky130_fd_sc_hd__clkbuf_2 output177 (.A(net177),
    .X(mem_la_addr[19]));
 sky130_fd_sc_hd__clkbuf_2 output178 (.A(net178),
    .X(mem_la_addr[1]));
 sky130_fd_sc_hd__clkbuf_2 output179 (.A(net179),
    .X(mem_la_addr[20]));
 sky130_fd_sc_hd__clkbuf_2 output180 (.A(net180),
    .X(mem_la_addr[21]));
 sky130_fd_sc_hd__clkbuf_2 output181 (.A(net181),
    .X(mem_la_addr[22]));
 sky130_fd_sc_hd__clkbuf_2 output182 (.A(net182),
    .X(mem_la_addr[23]));
 sky130_fd_sc_hd__clkbuf_2 output183 (.A(net183),
    .X(mem_la_addr[24]));
 sky130_fd_sc_hd__clkbuf_2 output184 (.A(net184),
    .X(mem_la_addr[25]));
 sky130_fd_sc_hd__clkbuf_2 output185 (.A(net185),
    .X(mem_la_addr[26]));
 sky130_fd_sc_hd__clkbuf_2 output186 (.A(net186),
    .X(mem_la_addr[27]));
 sky130_fd_sc_hd__clkbuf_2 output187 (.A(net187),
    .X(mem_la_addr[28]));
 sky130_fd_sc_hd__clkbuf_2 output188 (.A(net188),
    .X(mem_la_addr[29]));
 sky130_fd_sc_hd__clkbuf_2 output189 (.A(net189),
    .X(mem_la_addr[2]));
 sky130_fd_sc_hd__clkbuf_2 output190 (.A(net190),
    .X(mem_la_addr[30]));
 sky130_fd_sc_hd__clkbuf_2 output191 (.A(net191),
    .X(mem_la_addr[31]));
 sky130_fd_sc_hd__clkbuf_2 output192 (.A(net192),
    .X(mem_la_addr[3]));
 sky130_fd_sc_hd__clkbuf_2 output193 (.A(net193),
    .X(mem_la_addr[4]));
 sky130_fd_sc_hd__clkbuf_2 output194 (.A(net194),
    .X(mem_la_addr[5]));
 sky130_fd_sc_hd__clkbuf_2 output195 (.A(net195),
    .X(mem_la_addr[6]));
 sky130_fd_sc_hd__clkbuf_2 output196 (.A(net196),
    .X(mem_la_addr[7]));
 sky130_fd_sc_hd__clkbuf_2 output197 (.A(net197),
    .X(mem_la_addr[8]));
 sky130_fd_sc_hd__clkbuf_2 output198 (.A(net198),
    .X(mem_la_addr[9]));
 sky130_fd_sc_hd__clkbuf_2 output199 (.A(net199),
    .X(mem_la_read));
 sky130_fd_sc_hd__clkbuf_2 output200 (.A(net200),
    .X(mem_la_wdata[0]));
 sky130_fd_sc_hd__clkbuf_2 output201 (.A(net201),
    .X(mem_la_wdata[10]));
 sky130_fd_sc_hd__clkbuf_2 output202 (.A(net202),
    .X(mem_la_wdata[11]));
 sky130_fd_sc_hd__clkbuf_2 output203 (.A(net203),
    .X(mem_la_wdata[12]));
 sky130_fd_sc_hd__clkbuf_2 output204 (.A(net204),
    .X(mem_la_wdata[13]));
 sky130_fd_sc_hd__clkbuf_2 output205 (.A(net205),
    .X(mem_la_wdata[14]));
 sky130_fd_sc_hd__clkbuf_2 output206 (.A(net206),
    .X(mem_la_wdata[15]));
 sky130_fd_sc_hd__clkbuf_2 output207 (.A(net207),
    .X(mem_la_wdata[16]));
 sky130_fd_sc_hd__clkbuf_2 output208 (.A(net208),
    .X(mem_la_wdata[17]));
 sky130_fd_sc_hd__clkbuf_2 output209 (.A(net209),
    .X(mem_la_wdata[18]));
 sky130_fd_sc_hd__clkbuf_2 output210 (.A(net210),
    .X(mem_la_wdata[19]));
 sky130_fd_sc_hd__clkbuf_2 output211 (.A(net211),
    .X(mem_la_wdata[1]));
 sky130_fd_sc_hd__clkbuf_2 output212 (.A(net212),
    .X(mem_la_wdata[20]));
 sky130_fd_sc_hd__clkbuf_2 output213 (.A(net213),
    .X(mem_la_wdata[21]));
 sky130_fd_sc_hd__clkbuf_2 output214 (.A(net214),
    .X(mem_la_wdata[22]));
 sky130_fd_sc_hd__clkbuf_2 output215 (.A(net215),
    .X(mem_la_wdata[23]));
 sky130_fd_sc_hd__clkbuf_2 output216 (.A(net216),
    .X(mem_la_wdata[24]));
 sky130_fd_sc_hd__clkbuf_2 output217 (.A(net217),
    .X(mem_la_wdata[25]));
 sky130_fd_sc_hd__clkbuf_2 output218 (.A(net218),
    .X(mem_la_wdata[26]));
 sky130_fd_sc_hd__clkbuf_2 output219 (.A(net219),
    .X(mem_la_wdata[27]));
 sky130_fd_sc_hd__clkbuf_2 output220 (.A(net220),
    .X(mem_la_wdata[28]));
 sky130_fd_sc_hd__clkbuf_2 output221 (.A(net221),
    .X(mem_la_wdata[29]));
 sky130_fd_sc_hd__clkbuf_2 output222 (.A(net222),
    .X(mem_la_wdata[2]));
 sky130_fd_sc_hd__clkbuf_2 output223 (.A(net223),
    .X(mem_la_wdata[30]));
 sky130_fd_sc_hd__clkbuf_2 output224 (.A(net224),
    .X(mem_la_wdata[31]));
 sky130_fd_sc_hd__clkbuf_2 output225 (.A(net225),
    .X(mem_la_wdata[3]));
 sky130_fd_sc_hd__clkbuf_2 output226 (.A(net226),
    .X(mem_la_wdata[4]));
 sky130_fd_sc_hd__clkbuf_2 output227 (.A(net227),
    .X(mem_la_wdata[5]));
 sky130_fd_sc_hd__clkbuf_2 output228 (.A(net228),
    .X(mem_la_wdata[6]));
 sky130_fd_sc_hd__clkbuf_2 output229 (.A(net229),
    .X(mem_la_wdata[7]));
 sky130_fd_sc_hd__clkbuf_2 output230 (.A(net230),
    .X(mem_la_wdata[8]));
 sky130_fd_sc_hd__clkbuf_2 output231 (.A(net231),
    .X(mem_la_wdata[9]));
 sky130_fd_sc_hd__clkbuf_2 output232 (.A(net232),
    .X(mem_la_write));
 sky130_fd_sc_hd__clkbuf_2 output233 (.A(net233),
    .X(mem_la_wstrb[0]));
 sky130_fd_sc_hd__clkbuf_2 output234 (.A(net234),
    .X(mem_la_wstrb[1]));
 sky130_fd_sc_hd__clkbuf_2 output235 (.A(net235),
    .X(mem_la_wstrb[2]));
 sky130_fd_sc_hd__clkbuf_2 output236 (.A(net236),
    .X(mem_la_wstrb[3]));
 sky130_fd_sc_hd__clkbuf_2 output237 (.A(net237),
    .X(mem_valid));
 sky130_fd_sc_hd__clkbuf_2 output238 (.A(net238),
    .X(mem_wdata[0]));
 sky130_fd_sc_hd__clkbuf_2 output239 (.A(net239),
    .X(mem_wdata[10]));
 sky130_fd_sc_hd__clkbuf_2 output240 (.A(net240),
    .X(mem_wdata[11]));
 sky130_fd_sc_hd__clkbuf_2 output241 (.A(net241),
    .X(mem_wdata[12]));
 sky130_fd_sc_hd__clkbuf_2 output242 (.A(net242),
    .X(mem_wdata[13]));
 sky130_fd_sc_hd__clkbuf_2 output243 (.A(net243),
    .X(mem_wdata[14]));
 sky130_fd_sc_hd__clkbuf_2 output244 (.A(net244),
    .X(mem_wdata[15]));
 sky130_fd_sc_hd__clkbuf_2 output245 (.A(net245),
    .X(mem_wdata[16]));
 sky130_fd_sc_hd__clkbuf_2 output246 (.A(net246),
    .X(mem_wdata[17]));
 sky130_fd_sc_hd__clkbuf_2 output247 (.A(net247),
    .X(mem_wdata[18]));
 sky130_fd_sc_hd__clkbuf_2 output248 (.A(net248),
    .X(mem_wdata[19]));
 sky130_fd_sc_hd__clkbuf_2 output249 (.A(net249),
    .X(mem_wdata[1]));
 sky130_fd_sc_hd__clkbuf_2 output250 (.A(net250),
    .X(mem_wdata[20]));
 sky130_fd_sc_hd__clkbuf_2 output251 (.A(net251),
    .X(mem_wdata[21]));
 sky130_fd_sc_hd__clkbuf_2 output252 (.A(net252),
    .X(mem_wdata[22]));
 sky130_fd_sc_hd__clkbuf_2 output253 (.A(net253),
    .X(mem_wdata[23]));
 sky130_fd_sc_hd__clkbuf_2 output254 (.A(net254),
    .X(mem_wdata[24]));
 sky130_fd_sc_hd__clkbuf_2 output255 (.A(net255),
    .X(mem_wdata[25]));
 sky130_fd_sc_hd__clkbuf_2 output256 (.A(net256),
    .X(mem_wdata[26]));
 sky130_fd_sc_hd__clkbuf_2 output257 (.A(net257),
    .X(mem_wdata[27]));
 sky130_fd_sc_hd__clkbuf_2 output258 (.A(net258),
    .X(mem_wdata[28]));
 sky130_fd_sc_hd__clkbuf_2 output259 (.A(net259),
    .X(mem_wdata[29]));
 sky130_fd_sc_hd__clkbuf_2 output260 (.A(net260),
    .X(mem_wdata[2]));
 sky130_fd_sc_hd__clkbuf_2 output261 (.A(net261),
    .X(mem_wdata[30]));
 sky130_fd_sc_hd__clkbuf_2 output262 (.A(net262),
    .X(mem_wdata[31]));
 sky130_fd_sc_hd__clkbuf_2 output263 (.A(net263),
    .X(mem_wdata[3]));
 sky130_fd_sc_hd__clkbuf_2 output264 (.A(net264),
    .X(mem_wdata[4]));
 sky130_fd_sc_hd__clkbuf_2 output265 (.A(net265),
    .X(mem_wdata[5]));
 sky130_fd_sc_hd__clkbuf_2 output266 (.A(net266),
    .X(mem_wdata[6]));
 sky130_fd_sc_hd__clkbuf_2 output267 (.A(net267),
    .X(mem_wdata[7]));
 sky130_fd_sc_hd__clkbuf_2 output268 (.A(net268),
    .X(mem_wdata[8]));
 sky130_fd_sc_hd__clkbuf_2 output269 (.A(net269),
    .X(mem_wdata[9]));
 sky130_fd_sc_hd__clkbuf_2 output270 (.A(net270),
    .X(mem_wstrb[0]));
 sky130_fd_sc_hd__clkbuf_2 output271 (.A(net271),
    .X(mem_wstrb[1]));
 sky130_fd_sc_hd__clkbuf_2 output272 (.A(net272),
    .X(mem_wstrb[2]));
 sky130_fd_sc_hd__clkbuf_2 output273 (.A(net273),
    .X(mem_wstrb[3]));
 sky130_fd_sc_hd__clkbuf_2 output274 (.A(net274),
    .X(pcpi_insn[0]));
 sky130_fd_sc_hd__clkbuf_2 output275 (.A(net275),
    .X(pcpi_insn[10]));
 sky130_fd_sc_hd__clkbuf_2 output276 (.A(net276),
    .X(pcpi_insn[11]));
 sky130_fd_sc_hd__clkbuf_2 output277 (.A(net277),
    .X(pcpi_insn[12]));
 sky130_fd_sc_hd__clkbuf_2 output278 (.A(net278),
    .X(pcpi_insn[13]));
 sky130_fd_sc_hd__clkbuf_2 output279 (.A(net279),
    .X(pcpi_insn[14]));
 sky130_fd_sc_hd__clkbuf_2 output280 (.A(net280),
    .X(pcpi_insn[15]));
 sky130_fd_sc_hd__clkbuf_2 output281 (.A(net281),
    .X(pcpi_insn[16]));
 sky130_fd_sc_hd__clkbuf_2 output282 (.A(net282),
    .X(pcpi_insn[17]));
 sky130_fd_sc_hd__clkbuf_2 output283 (.A(net283),
    .X(pcpi_insn[18]));
 sky130_fd_sc_hd__clkbuf_2 output284 (.A(net284),
    .X(pcpi_insn[19]));
 sky130_fd_sc_hd__clkbuf_2 output285 (.A(net285),
    .X(pcpi_insn[1]));
 sky130_fd_sc_hd__clkbuf_2 output286 (.A(net286),
    .X(pcpi_insn[20]));
 sky130_fd_sc_hd__clkbuf_2 output287 (.A(net287),
    .X(pcpi_insn[21]));
 sky130_fd_sc_hd__clkbuf_2 output288 (.A(net288),
    .X(pcpi_insn[22]));
 sky130_fd_sc_hd__clkbuf_2 output289 (.A(net289),
    .X(pcpi_insn[23]));
 sky130_fd_sc_hd__clkbuf_2 output290 (.A(net290),
    .X(pcpi_insn[24]));
 sky130_fd_sc_hd__clkbuf_2 output291 (.A(net291),
    .X(pcpi_insn[25]));
 sky130_fd_sc_hd__clkbuf_2 output292 (.A(net292),
    .X(pcpi_insn[26]));
 sky130_fd_sc_hd__clkbuf_2 output293 (.A(net293),
    .X(pcpi_insn[27]));
 sky130_fd_sc_hd__clkbuf_2 output294 (.A(net294),
    .X(pcpi_insn[28]));
 sky130_fd_sc_hd__clkbuf_2 output295 (.A(net295),
    .X(pcpi_insn[29]));
 sky130_fd_sc_hd__clkbuf_2 output296 (.A(net296),
    .X(pcpi_insn[2]));
 sky130_fd_sc_hd__clkbuf_2 output297 (.A(net297),
    .X(pcpi_insn[30]));
 sky130_fd_sc_hd__clkbuf_2 output298 (.A(net298),
    .X(pcpi_insn[31]));
 sky130_fd_sc_hd__clkbuf_2 output299 (.A(net299),
    .X(pcpi_insn[3]));
 sky130_fd_sc_hd__clkbuf_2 output300 (.A(net300),
    .X(pcpi_insn[4]));
 sky130_fd_sc_hd__clkbuf_2 output301 (.A(net301),
    .X(pcpi_insn[5]));
 sky130_fd_sc_hd__clkbuf_2 output302 (.A(net302),
    .X(pcpi_insn[6]));
 sky130_fd_sc_hd__clkbuf_2 output303 (.A(net303),
    .X(pcpi_insn[7]));
 sky130_fd_sc_hd__clkbuf_2 output304 (.A(net304),
    .X(pcpi_insn[8]));
 sky130_fd_sc_hd__clkbuf_2 output305 (.A(net305),
    .X(pcpi_insn[9]));
 sky130_fd_sc_hd__clkbuf_2 output306 (.A(net306),
    .X(pcpi_rs1[0]));
 sky130_fd_sc_hd__clkbuf_2 output307 (.A(net307),
    .X(pcpi_rs1[10]));
 sky130_fd_sc_hd__clkbuf_2 output308 (.A(net308),
    .X(pcpi_rs1[11]));
 sky130_fd_sc_hd__clkbuf_2 output309 (.A(net309),
    .X(pcpi_rs1[12]));
 sky130_fd_sc_hd__clkbuf_2 output310 (.A(net310),
    .X(pcpi_rs1[13]));
 sky130_fd_sc_hd__clkbuf_2 output311 (.A(net311),
    .X(pcpi_rs1[14]));
 sky130_fd_sc_hd__clkbuf_2 output312 (.A(net312),
    .X(pcpi_rs1[15]));
 sky130_fd_sc_hd__clkbuf_2 output313 (.A(net313),
    .X(pcpi_rs1[16]));
 sky130_fd_sc_hd__clkbuf_2 output314 (.A(net314),
    .X(pcpi_rs1[17]));
 sky130_fd_sc_hd__clkbuf_2 output315 (.A(net315),
    .X(pcpi_rs1[18]));
 sky130_fd_sc_hd__clkbuf_2 output316 (.A(net316),
    .X(pcpi_rs1[19]));
 sky130_fd_sc_hd__clkbuf_2 output317 (.A(net317),
    .X(pcpi_rs1[1]));
 sky130_fd_sc_hd__clkbuf_2 output318 (.A(net318),
    .X(pcpi_rs1[20]));
 sky130_fd_sc_hd__clkbuf_2 output319 (.A(net319),
    .X(pcpi_rs1[21]));
 sky130_fd_sc_hd__clkbuf_2 output320 (.A(net320),
    .X(pcpi_rs1[22]));
 sky130_fd_sc_hd__clkbuf_2 output321 (.A(net321),
    .X(pcpi_rs1[23]));
 sky130_fd_sc_hd__clkbuf_2 output322 (.A(net322),
    .X(pcpi_rs1[24]));
 sky130_fd_sc_hd__clkbuf_2 output323 (.A(net323),
    .X(pcpi_rs1[25]));
 sky130_fd_sc_hd__clkbuf_2 output324 (.A(net324),
    .X(pcpi_rs1[26]));
 sky130_fd_sc_hd__clkbuf_2 output325 (.A(net325),
    .X(pcpi_rs1[27]));
 sky130_fd_sc_hd__clkbuf_2 output326 (.A(net326),
    .X(pcpi_rs1[28]));
 sky130_fd_sc_hd__clkbuf_2 output327 (.A(net327),
    .X(pcpi_rs1[29]));
 sky130_fd_sc_hd__clkbuf_2 output328 (.A(net328),
    .X(pcpi_rs1[2]));
 sky130_fd_sc_hd__clkbuf_2 output329 (.A(net329),
    .X(pcpi_rs1[30]));
 sky130_fd_sc_hd__clkbuf_2 output330 (.A(net330),
    .X(pcpi_rs1[31]));
 sky130_fd_sc_hd__clkbuf_2 output331 (.A(net331),
    .X(pcpi_rs1[3]));
 sky130_fd_sc_hd__clkbuf_2 output332 (.A(net332),
    .X(pcpi_rs1[4]));
 sky130_fd_sc_hd__clkbuf_2 output333 (.A(net333),
    .X(pcpi_rs1[5]));
 sky130_fd_sc_hd__clkbuf_2 output334 (.A(net334),
    .X(pcpi_rs1[6]));
 sky130_fd_sc_hd__clkbuf_2 output335 (.A(net335),
    .X(pcpi_rs1[7]));
 sky130_fd_sc_hd__clkbuf_2 output336 (.A(net336),
    .X(pcpi_rs1[8]));
 sky130_fd_sc_hd__clkbuf_2 output337 (.A(net337),
    .X(pcpi_rs1[9]));
 sky130_fd_sc_hd__clkbuf_2 output338 (.A(net338),
    .X(pcpi_rs2[0]));
 sky130_fd_sc_hd__clkbuf_2 output339 (.A(net339),
    .X(pcpi_rs2[10]));
 sky130_fd_sc_hd__clkbuf_2 output340 (.A(net340),
    .X(pcpi_rs2[11]));
 sky130_fd_sc_hd__clkbuf_2 output341 (.A(net341),
    .X(pcpi_rs2[12]));
 sky130_fd_sc_hd__clkbuf_2 output342 (.A(net342),
    .X(pcpi_rs2[13]));
 sky130_fd_sc_hd__clkbuf_2 output343 (.A(net343),
    .X(pcpi_rs2[14]));
 sky130_fd_sc_hd__clkbuf_2 output344 (.A(net344),
    .X(pcpi_rs2[15]));
 sky130_fd_sc_hd__clkbuf_2 output345 (.A(net345),
    .X(pcpi_rs2[16]));
 sky130_fd_sc_hd__clkbuf_2 output346 (.A(net346),
    .X(pcpi_rs2[17]));
 sky130_fd_sc_hd__clkbuf_2 output347 (.A(net347),
    .X(pcpi_rs2[18]));
 sky130_fd_sc_hd__clkbuf_2 output348 (.A(net348),
    .X(pcpi_rs2[19]));
 sky130_fd_sc_hd__clkbuf_2 output349 (.A(net349),
    .X(pcpi_rs2[1]));
 sky130_fd_sc_hd__clkbuf_2 output350 (.A(net350),
    .X(pcpi_rs2[20]));
 sky130_fd_sc_hd__clkbuf_2 output351 (.A(net351),
    .X(pcpi_rs2[21]));
 sky130_fd_sc_hd__clkbuf_2 output352 (.A(net352),
    .X(pcpi_rs2[22]));
 sky130_fd_sc_hd__clkbuf_2 output353 (.A(net353),
    .X(pcpi_rs2[23]));
 sky130_fd_sc_hd__clkbuf_2 output354 (.A(net354),
    .X(pcpi_rs2[24]));
 sky130_fd_sc_hd__clkbuf_2 output355 (.A(net355),
    .X(pcpi_rs2[25]));
 sky130_fd_sc_hd__clkbuf_2 output356 (.A(net356),
    .X(pcpi_rs2[26]));
 sky130_fd_sc_hd__clkbuf_2 output357 (.A(net357),
    .X(pcpi_rs2[27]));
 sky130_fd_sc_hd__clkbuf_2 output358 (.A(net358),
    .X(pcpi_rs2[28]));
 sky130_fd_sc_hd__clkbuf_2 output359 (.A(net359),
    .X(pcpi_rs2[29]));
 sky130_fd_sc_hd__clkbuf_2 output360 (.A(net360),
    .X(pcpi_rs2[2]));
 sky130_fd_sc_hd__clkbuf_2 output361 (.A(net361),
    .X(pcpi_rs2[30]));
 sky130_fd_sc_hd__clkbuf_2 output362 (.A(net362),
    .X(pcpi_rs2[31]));
 sky130_fd_sc_hd__clkbuf_2 output363 (.A(net363),
    .X(pcpi_rs2[3]));
 sky130_fd_sc_hd__clkbuf_2 output364 (.A(net364),
    .X(pcpi_rs2[4]));
 sky130_fd_sc_hd__clkbuf_2 output365 (.A(net365),
    .X(pcpi_rs2[5]));
 sky130_fd_sc_hd__clkbuf_2 output366 (.A(net366),
    .X(pcpi_rs2[6]));
 sky130_fd_sc_hd__clkbuf_2 output367 (.A(net367),
    .X(pcpi_rs2[7]));
 sky130_fd_sc_hd__clkbuf_2 output368 (.A(net368),
    .X(pcpi_rs2[8]));
 sky130_fd_sc_hd__clkbuf_2 output369 (.A(net369),
    .X(pcpi_rs2[9]));
 sky130_fd_sc_hd__clkbuf_2 output370 (.A(net370),
    .X(pcpi_valid));
 sky130_fd_sc_hd__clkbuf_2 output371 (.A(net371),
    .X(trace_data[0]));
 sky130_fd_sc_hd__clkbuf_2 output372 (.A(net372),
    .X(trace_data[10]));
 sky130_fd_sc_hd__clkbuf_2 output373 (.A(net373),
    .X(trace_data[11]));
 sky130_fd_sc_hd__clkbuf_2 output374 (.A(net374),
    .X(trace_data[12]));
 sky130_fd_sc_hd__clkbuf_2 output375 (.A(net375),
    .X(trace_data[13]));
 sky130_fd_sc_hd__clkbuf_2 output376 (.A(net376),
    .X(trace_data[14]));
 sky130_fd_sc_hd__clkbuf_2 output377 (.A(net377),
    .X(trace_data[15]));
 sky130_fd_sc_hd__clkbuf_2 output378 (.A(net378),
    .X(trace_data[16]));
 sky130_fd_sc_hd__clkbuf_2 output379 (.A(net379),
    .X(trace_data[17]));
 sky130_fd_sc_hd__clkbuf_2 output380 (.A(net380),
    .X(trace_data[18]));
 sky130_fd_sc_hd__clkbuf_2 output381 (.A(net381),
    .X(trace_data[19]));
 sky130_fd_sc_hd__clkbuf_2 output382 (.A(net382),
    .X(trace_data[1]));
 sky130_fd_sc_hd__clkbuf_2 output383 (.A(net383),
    .X(trace_data[20]));
 sky130_fd_sc_hd__clkbuf_2 output384 (.A(net384),
    .X(trace_data[21]));
 sky130_fd_sc_hd__clkbuf_2 output385 (.A(net385),
    .X(trace_data[22]));
 sky130_fd_sc_hd__clkbuf_2 output386 (.A(net386),
    .X(trace_data[23]));
 sky130_fd_sc_hd__clkbuf_2 output387 (.A(net387),
    .X(trace_data[24]));
 sky130_fd_sc_hd__clkbuf_2 output388 (.A(net388),
    .X(trace_data[25]));
 sky130_fd_sc_hd__clkbuf_2 output389 (.A(net389),
    .X(trace_data[26]));
 sky130_fd_sc_hd__clkbuf_2 output390 (.A(net390),
    .X(trace_data[27]));
 sky130_fd_sc_hd__clkbuf_2 output391 (.A(net391),
    .X(trace_data[28]));
 sky130_fd_sc_hd__clkbuf_2 output392 (.A(net392),
    .X(trace_data[29]));
 sky130_fd_sc_hd__clkbuf_2 output393 (.A(net393),
    .X(trace_data[2]));
 sky130_fd_sc_hd__clkbuf_2 output394 (.A(net394),
    .X(trace_data[30]));
 sky130_fd_sc_hd__clkbuf_2 output395 (.A(net395),
    .X(trace_data[31]));
 sky130_fd_sc_hd__clkbuf_2 output396 (.A(net396),
    .X(trace_data[32]));
 sky130_fd_sc_hd__clkbuf_2 output397 (.A(net397),
    .X(trace_data[33]));
 sky130_fd_sc_hd__clkbuf_2 output398 (.A(net398),
    .X(trace_data[34]));
 sky130_fd_sc_hd__clkbuf_2 output399 (.A(net399),
    .X(trace_data[35]));
 sky130_fd_sc_hd__clkbuf_2 output400 (.A(net400),
    .X(trace_data[3]));
 sky130_fd_sc_hd__clkbuf_2 output401 (.A(net401),
    .X(trace_data[4]));
 sky130_fd_sc_hd__clkbuf_2 output402 (.A(net402),
    .X(trace_data[5]));
 sky130_fd_sc_hd__clkbuf_2 output403 (.A(net403),
    .X(trace_data[6]));
 sky130_fd_sc_hd__clkbuf_2 output404 (.A(net404),
    .X(trace_data[7]));
 sky130_fd_sc_hd__clkbuf_2 output405 (.A(net405),
    .X(trace_data[8]));
 sky130_fd_sc_hd__clkbuf_2 output406 (.A(net406),
    .X(trace_data[9]));
 sky130_fd_sc_hd__clkbuf_2 output407 (.A(net407),
    .X(trace_valid));
 sky130_fd_sc_hd__clkbuf_2 output408 (.A(net408),
    .X(trap));
 sky130_fd_sc_hd__buf_6 repeater409 (.A(_01208_),
    .X(net409));
 sky130_fd_sc_hd__buf_8 repeater410 (.A(_00308_),
    .X(net410));
 sky130_fd_sc_hd__buf_6 repeater411 (.A(_00308_),
    .X(net411));
 sky130_fd_sc_hd__buf_12 repeater412 (.A(_14285_),
    .X(net412));
 sky130_fd_sc_hd__buf_6 repeater413 (.A(_11844_),
    .X(net413));
 sky130_fd_sc_hd__clkbuf_16 repeater414 (.A(_02069_),
    .X(net414));
 sky130_fd_sc_hd__buf_8 repeater415 (.A(mem_xfer),
    .X(net415));
 sky130_fd_sc_hd__buf_8 repeater416 (.A(net419),
    .X(net416));
 sky130_fd_sc_hd__buf_8 repeater417 (.A(net418),
    .X(net417));
 sky130_fd_sc_hd__buf_6 repeater418 (.A(net419),
    .X(net418));
 sky130_fd_sc_hd__buf_8 repeater419 (.A(_00301_),
    .X(net419));
 sky130_fd_sc_hd__buf_8 repeater420 (.A(net421),
    .X(net420));
 sky130_fd_sc_hd__buf_6 repeater421 (.A(_01683_),
    .X(net421));
 sky130_fd_sc_hd__buf_8 repeater422 (.A(_01683_),
    .X(net422));
 sky130_fd_sc_hd__buf_8 repeater423 (.A(net424),
    .X(net423));
 sky130_fd_sc_hd__buf_8 repeater424 (.A(_00297_),
    .X(net424));
 sky130_fd_sc_hd__buf_8 repeater425 (.A(_00292_),
    .X(net425));
 sky130_fd_sc_hd__buf_8 repeater426 (.A(_01714_),
    .X(net426));
 sky130_fd_sc_hd__buf_12 repeater427 (.A(net428),
    .X(net427));
 sky130_fd_sc_hd__buf_12 repeater428 (.A(_00368_),
    .X(net428));
 sky130_fd_sc_hd__buf_6 repeater429 (.A(net430),
    .X(net429));
 sky130_fd_sc_hd__buf_4 repeater430 (.A(_01717_),
    .X(net430));
 sky130_fd_sc_hd__buf_12 repeater431 (.A(_00309_),
    .X(net431));
 sky130_fd_sc_hd__buf_12 repeater432 (.A(net435),
    .X(net432));
 sky130_fd_sc_hd__clkbuf_8 repeater433 (.A(net435),
    .X(net433));
 sky130_fd_sc_hd__buf_12 repeater434 (.A(net436),
    .X(net434));
 sky130_fd_sc_hd__buf_8 repeater435 (.A(net436),
    .X(net435));
 sky130_fd_sc_hd__buf_12 repeater436 (.A(net437),
    .X(net436));
 sky130_fd_sc_hd__buf_12 repeater437 (.A(net438),
    .X(net437));
 sky130_fd_sc_hd__buf_12 repeater438 (.A(net439),
    .X(net438));
 sky130_fd_sc_hd__buf_8 repeater439 (.A(net442),
    .X(net439));
 sky130_fd_sc_hd__buf_12 repeater440 (.A(net441),
    .X(net440));
 sky130_fd_sc_hd__clkbuf_8 repeater441 (.A(net443),
    .X(net441));
 sky130_fd_sc_hd__buf_12 repeater442 (.A(net443),
    .X(net442));
 sky130_fd_sc_hd__buf_12 repeater443 (.A(_00357_),
    .X(net443));
 sky130_fd_sc_hd__buf_12 repeater444 (.A(net446),
    .X(net444));
 sky130_fd_sc_hd__buf_8 repeater445 (.A(net446),
    .X(net445));
 sky130_fd_sc_hd__buf_12 repeater446 (.A(net447),
    .X(net446));
 sky130_fd_sc_hd__buf_12 repeater447 (.A(net448),
    .X(net447));
 sky130_fd_sc_hd__buf_12 repeater448 (.A(net450),
    .X(net448));
 sky130_fd_sc_hd__buf_12 repeater449 (.A(_00358_),
    .X(net449));
 sky130_fd_sc_hd__buf_12 repeater450 (.A(_00358_),
    .X(net450));
 sky130_fd_sc_hd__buf_12 repeater451 (.A(_00360_),
    .X(net451));
 sky130_fd_sc_hd__buf_8 repeater452 (.A(_00360_),
    .X(net452));
 sky130_fd_sc_hd__buf_12 repeater453 (.A(net454),
    .X(net453));
 sky130_fd_sc_hd__buf_12 repeater454 (.A(_00362_),
    .X(net454));
 sky130_fd_sc_hd__buf_8 repeater455 (.A(_01816_),
    .X(net455));
 sky130_fd_sc_hd__buf_8 repeater456 (.A(_01304_),
    .X(net456));
 sky130_fd_sc_hd__buf_4 repeater457 (.A(_01304_),
    .X(net457));
 sky130_fd_sc_hd__clkbuf_16 repeater458 (.A(net226),
    .X(net458));
 sky130_fd_sc_hd__clkbuf_16 repeater459 (.A(net225),
    .X(net459));
 sky130_fd_sc_hd__clkbuf_16 repeater460 (.A(net222),
    .X(net460));
 sky130_fd_sc_hd__clkbuf_16 repeater461 (.A(net211),
    .X(net461));
 sky130_fd_sc_hd__clkbuf_16 repeater462 (.A(net200),
    .X(net462));
 sky130_fd_sc_hd__clkbuf_16 repeater463 (.A(\cpu_state[3] ),
    .X(net463));
 sky130_fd_sc_hd__buf_8 repeater464 (.A(net45),
    .X(net464));
 sky130_fd_sc_hd__buf_8 repeater465 (.A(net21),
    .X(net465));
 sky130_fd_sc_hd__buf_8 repeater466 (.A(net20),
    .X(net466));
 sky130_fd_sc_hd__buf_8 repeater467 (.A(net13),
    .X(net467));
endmodule
